* Substrate SPICE library
* This is a generated file. Be careful when editing manually: this file may be overwritten.


.SUBCKT sky130_fd_sc_hs__nand2_4 A B VGND VNB VPB VPWR Y

  X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X1 Y A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X2 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X3 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X4 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X5 a_27_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X6 Y A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X7 VPWR B Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X8 Y B VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X9 a_27_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X11 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740


.ENDS sky130_fd_sc_hs__nand2_4

.SUBCKT sky130_fd_sc_hs__nand2_4_wrapper A B VGND VNB VPB VPWR Y

  X0 A B VGND VNB VPB VPWR Y sky130_fd_sc_hs__nand2_4

.ENDS sky130_fd_sc_hs__nand2_4_wrapper

.SUBCKT sky130_fd_sc_hs__nand2_8 A B VGND VNB VPB VPWR Y

  X0 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X1 Y A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X2 Y B VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X3 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X4 Y A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X5 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X6 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X7 a_27_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X9 Y A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X10 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X11 a_27_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X12 VPWR B Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X13 VPWR B Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X14 a_27_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X15 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X16 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X17 VGND B a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X18 a_27_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X19 Y B VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X20 a_27_74# A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X21 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X22 Y A a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X23 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120


.ENDS sky130_fd_sc_hs__nand2_8

.SUBCKT sky130_fd_sc_hs__nand2_8_wrapper A B VGND VNB VPB VPWR Y

  X0 A B VGND VNB VPB VPWR Y sky130_fd_sc_hs__nand2_8

.ENDS sky130_fd_sc_hs__nand2_8_wrapper

.SUBCKT mos_w5000_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=5.000


.ENDS mos_w5000_l150_m1_nf1_id1

.SUBCKT mos_w3230_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=3.230


.ENDS mos_w3230_l150_m1_nf1_id1

.SUBCKT mos_w800_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.800


.ENDS mos_w800_l150_m1_nf1_id1

.SUBCKT mos_w500_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.500


.ENDS mos_w500_l150_m1_nf1_id1

.SUBCKT precharge vdd bl br en_b

  Xbl_pull_up bl en_b vdd vdd mos_w800_l150_m1_nf1_id1
  Xbr_pull_up br en_b vdd vdd mos_w800_l150_m1_nf1_id1
  Xequalizer bl en_b br vdd mos_w500_l150_m1_nf1_id1

.ENDS precharge

.SUBCKT sky130_fd_sc_hs__and2_4 A B VGND VNB VPB VPWR X

  X0 VPWR a_83_269# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X1 VPWR B a_83_269# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.840

  X2 VPWR a_83_269# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X3 a_504_119# B VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X4 a_83_269# A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.840

  X5 VGND B a_504_119# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X6 VGND a_83_269# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X7 a_83_269# B VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.840

  X8 X a_83_269# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X9 VGND a_83_269# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X10 X a_83_269# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X11 X a_83_269# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X12 a_504_119# A a_83_269# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X13 a_83_269# A a_504_119# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X14 VPWR A a_83_269# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.840

  X15 X a_83_269# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740


.ENDS sky130_fd_sc_hs__and2_4

.SUBCKT sky130_fd_sc_hs__and2_4_wrapper A B VGND VNB VPB VPWR X

  X0 A B VGND VNB VPB VPWR X sky130_fd_sc_hs__and2_4

.ENDS sky130_fd_sc_hs__and2_4_wrapper

.SUBCKT mos_w2000_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=2.000


.ENDS mos_w2000_l150_m1_nf1_id0

.SUBCKT mos_w2500_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=2.500


.ENDS mos_w2500_l150_m1_nf1_id1

.SUBCKT nand2 vdd vss a b y

  Xn1 x a vss vss mos_w2000_l150_m1_nf1_id0
  Xn2 y b x vss mos_w2000_l150_m1_nf1_id0
  Xp1 y a vdd vdd mos_w2500_l150_m1_nf1_id1
  Xp2 y b vdd vdd mos_w2500_l150_m1_nf1_id1

.ENDS nand2

.SUBCKT folded_inv_1 vdd vss a y

  XMP0 y a vdd vdd mos_w5000_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w2000_l150_m1_nf1_id0
  XMP1 y a vdd vdd mos_w5000_l150_m1_nf1_id1
  XMN1 y a vss vss mos_w2000_l150_m1_nf1_id0

.ENDS folded_inv_1

.SUBCKT and2 vdd a b y yb vss

  X0 vdd vss a b yb nand2
  X0_1 vdd vss yb y folded_inv_1

.ENDS and2

.SUBCKT sky130_fd_sc_hs__dfrbp_2 CLK D RESET_B VGND VNB VPB VPWR Q Q_N

  X0 a_1800_291# a_1586_149# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.420

  X1 VGND CLK a_728_331# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X2 Q a_2363_352# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X3 VPWR CLK a_728_331# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X4 a_1499_149# a_728_331# a_1586_149# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.420

  X5 a_536_81# a_331_392# a_614_81# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.420

  X6 a_156_74# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.420

  X7 a_298_294# a_818_418# a_614_81# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.420

  X8 a_70_74# a_728_331# a_298_294# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.420

  X9 a_331_392# a_728_331# a_1586_149# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X10 a_70_74# D a_156_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.420

  X11 a_818_418# a_728_331# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X12 a_818_418# a_728_331# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X13 a_1586_149# a_818_418# a_1755_389# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.420

  X14 Q_N a_1586_149# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X15 a_298_294# a_818_418# a_70_74# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.420

  X16 VGND RESET_B a_536_81# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.420

  X17 a_1755_389# a_1800_291# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.420

  X18 a_1586_149# a_818_418# a_331_392# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X19 Q a_2363_352# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X20 VGND a_1586_149# Q_N VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X21 VGND a_1586_149# a_2363_352# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X22 VPWR a_298_294# a_331_392# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X23 a_298_294# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.420

  X24 a_1499_149# a_1800_291# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.420

  X25 VPWR a_331_392# a_683_485# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.420

  X26 VPWR D a_70_74# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.420

  X27 VPWR RESET_B a_1800_291# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.420

  X28 a_1974_74# a_1586_149# a_1800_291# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.420

  X29 a_70_74# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.420

  X30 Q_N a_1586_149# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X31 VPWR a_1586_149# a_2363_352# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X32 VGND a_2363_352# Q VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X33 VPWR a_1586_149# Q_N VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X34 VGND RESET_B a_1974_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.420

  X35 a_683_485# a_728_331# a_298_294# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.420

  X36 VGND a_298_294# a_331_392# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X37 VPWR a_2363_352# Q VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120


.ENDS sky130_fd_sc_hs__dfrbp_2

.SUBCKT sky130_fd_sc_hs__dfrbp_2_wrapper CLK D RESET_B VGND VNB VPB VPWR Q Q_N

  X0 CLK D RESET_B VGND VNB VPB VPWR Q Q_N sky130_fd_sc_hs__dfrbp_2

.ENDS sky130_fd_sc_hs__dfrbp_2_wrapper

.SUBCKT sramgen_svt_inv_2 A VGND VNB VPB VPWR Y

  X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X2 VGND A Y VNB sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.740

  X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.740


.ENDS sramgen_svt_inv_2

.SUBCKT sramgen_svt_inv_2_wrapper A VGND VNB VPB VPWR Y

  X0 A VGND VNB VPB VPWR Y sramgen_svt_inv_2

.ENDS sramgen_svt_inv_2_wrapper

.SUBCKT sramgen_svt_inv_4 A VGND VNB VPB VPWR Y

  X0 VGND A Y VNB sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.740

  X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.740

  X4 Y A VGND VNB sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.740

  X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.740


.ENDS sramgen_svt_inv_4

.SUBCKT sramgen_svt_inv_4_wrapper A VGND VNB VPB VPWR Y

  X0 A VGND VNB VPB VPWR Y sramgen_svt_inv_4

.ENDS sramgen_svt_inv_4_wrapper

.SUBCKT svt_inv_chain_22 din dout vdd vss

  Xinv0 din vss vss vdd vdd x[0] sramgen_svt_inv_2_wrapper
  Xinv1 x[0] vss vss vdd vdd x[1] sramgen_svt_inv_2_wrapper
  Xinv2 x[1] vss vss vdd vdd x[2] sramgen_svt_inv_2_wrapper
  Xinv3 x[2] vss vss vdd vdd x[3] sramgen_svt_inv_2_wrapper
  Xinv4 x[3] vss vss vdd vdd x[4] sramgen_svt_inv_2_wrapper
  Xinv5 x[4] vss vss vdd vdd x[5] sramgen_svt_inv_2_wrapper
  Xinv6 x[5] vss vss vdd vdd x[6] sramgen_svt_inv_2_wrapper
  Xinv7 x[6] vss vss vdd vdd x[7] sramgen_svt_inv_2_wrapper
  Xinv8 x[7] vss vss vdd vdd x[8] sramgen_svt_inv_2_wrapper
  Xinv9 x[8] vss vss vdd vdd x[9] sramgen_svt_inv_2_wrapper
  Xinv10 x[9] vss vss vdd vdd x[10] sramgen_svt_inv_2_wrapper
  Xinv11 x[10] vss vss vdd vdd x[11] sramgen_svt_inv_2_wrapper
  Xinv12 x[11] vss vss vdd vdd x[12] sramgen_svt_inv_2_wrapper
  Xinv13 x[12] vss vss vdd vdd x[13] sramgen_svt_inv_2_wrapper
  Xinv14 x[13] vss vss vdd vdd x[14] sramgen_svt_inv_2_wrapper
  Xinv15 x[14] vss vss vdd vdd x[15] sramgen_svt_inv_2_wrapper
  Xinv16 x[15] vss vss vdd vdd x[16] sramgen_svt_inv_2_wrapper
  Xinv17 x[16] vss vss vdd vdd x[17] sramgen_svt_inv_2_wrapper
  Xinv18 x[17] vss vss vdd vdd x[18] sramgen_svt_inv_2_wrapper
  Xinv19 x[18] vss vss vdd vdd x[19] sramgen_svt_inv_2_wrapper
  Xinv20 x[19] vss vss vdd vdd x[20] sramgen_svt_inv_2_wrapper
  Xinv21 x[20] vss vss vdd vdd dout sramgen_svt_inv_4_wrapper

.ENDS svt_inv_chain_22

.SUBCKT mos_w700_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=0.700


.ENDS mos_w700_l150_m1_nf1_id1

.SUBCKT mos_w700_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.700


.ENDS mos_w700_l150_m1_nf1_id0

.SUBCKT multi_finger_inv_4 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP8 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP9 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP10 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP11 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP12 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP13 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP14 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP15 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP16 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP17 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP18 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP19 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP20 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP21 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP22 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP23 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP24 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP25 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP26 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP27 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP28 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP29 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP30 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP31 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP32 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP33 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP34 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP35 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP36 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP37 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP38 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP39 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP40 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP41 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP42 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP43 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP44 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP45 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP46 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP47 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP48 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP49 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP50 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP51 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP52 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP53 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP54 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN3 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN4 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN5 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN6 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN7 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN8 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN9 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN10 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN11 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN12 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN13 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN14 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN15 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN16 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN17 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN18 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN19 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN20 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN21 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_4

.SUBCKT multi_finger_inv_13 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP8 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP9 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP10 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP11 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP12 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP13 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP14 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP15 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP16 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP17 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP18 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP19 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP20 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP21 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP22 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP23 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP24 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP25 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP26 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP27 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP28 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP29 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP30 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP31 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP32 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP33 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP34 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP35 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP36 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP37 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP38 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP39 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP40 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP41 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP42 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP43 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP44 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP45 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP46 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP47 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP48 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP49 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP50 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP51 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN3 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN4 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN5 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN6 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN7 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN8 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN9 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN10 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN11 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN12 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN13 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN14 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN15 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN16 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN17 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN18 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN19 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN20 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_13

.SUBCKT mos_w1000_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000


.ENDS mos_w1000_l150_m1_nf1_id1

.SUBCKT mos_w600_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.600


.ENDS mos_w600_l150_m1_nf1_id0

.SUBCKT folded_inv_6 vdd vss a y

  XMP0 y a vdd vdd mos_w1000_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w600_l150_m1_nf1_id0
  XMP1 y a vdd vdd mos_w1000_l150_m1_nf1_id1
  XMN1 y a vss vss mos_w600_l150_m1_nf1_id0

.ENDS folded_inv_6

.SUBCKT mos_w1000_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=1.000


.ENDS mos_w1000_l150_m1_nf1_id0

.SUBCKT diff_latch vdd vss din1 din2 dout1 dout2

  Xinbuf_1 vdd vss din1 rst folded_inv_6
  Xinbuf_2 vdd vss din2 set folded_inv_6
  Xoutbuf_1 vdd vss q dout2 folded_inv_6
  Xoutbuf_2 vdd vss qb dout1 folded_inv_6
  Xinvq_1 vdd vss q qb folded_inv_6
  Xinvq_2 vdd vss qb q folded_inv_6
  XMN10 q rst vss vss mos_w1000_l150_m1_nf1_id0
  XMN11 q rst vss vss mos_w1000_l150_m1_nf1_id0
  XMN20 qb set vss vss mos_w1000_l150_m1_nf1_id0
  XMN21 qb set vss vss mos_w1000_l150_m1_nf1_id0

.ENDS diff_latch

.SUBCKT sky130_fd_sc_hs__inv_2 A VGND VNB VPB VPWR Y

  X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X2 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X3 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740


.ENDS sky130_fd_sc_hs__inv_2

.SUBCKT decoder_stage vdd vss y[0] y[1] y[2] y[3] y[4] y[5] y[6] y[7] y[8] y[9] y[10] y[11] y_b[0] y_b[1] y_b[2] y_b[3] y_b[4] y_b[5] y_b[6] y_b[7] y_b[8] y_b[9] y_b[10] y_b[11] wl_en in[0] in[1] in[2] in[3] in[4] in[5] in[6] in[7] in[8] in[9] in[10] in[11]

  Xgate_0_0_0 vdd wl_en in[0] y[0] y_b[0] vss and2
  Xgate_0_1_0 vdd wl_en in[1] y[1] y_b[1] vss and2
  Xgate_0_2_0 vdd wl_en in[2] y[2] y_b[2] vss and2
  Xgate_0_3_0 vdd wl_en in[3] y[3] y_b[3] vss and2
  Xgate_0_4_0 vdd wl_en in[4] y[4] y_b[4] vss and2
  Xgate_0_5_0 vdd wl_en in[5] y[5] y_b[5] vss and2
  Xgate_0_6_0 vdd wl_en in[6] y[6] y_b[6] vss and2
  Xgate_0_7_0 vdd wl_en in[7] y[7] y_b[7] vss and2
  Xgate_0_8_0 vdd wl_en in[8] y[8] y_b[8] vss and2
  Xgate_0_9_0 vdd wl_en in[9] y[9] y_b[9] vss and2
  Xgate_0_10_0 vdd wl_en in[10] y[10] y_b[10] vss and2
  Xgate_0_11_0 vdd wl_en in[11] y[11] y_b[11] vss and2

.ENDS decoder_stage

.SUBCKT mos_w3000_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=3.000


.ENDS mos_w3000_l150_m1_nf1_id0

.SUBCKT nand3 vdd vss a b c y

  Xn1 x1 a vss vss mos_w3000_l150_m1_nf1_id0
  Xn2 x2 b x1 vss mos_w3000_l150_m1_nf1_id0
  Xn3 y c x2 vss mos_w3000_l150_m1_nf1_id0
  Xp1 y a vdd vdd mos_w2500_l150_m1_nf1_id1
  Xp2 y b vdd vdd mos_w2500_l150_m1_nf1_id1
  Xp3 y c vdd vdd mos_w2500_l150_m1_nf1_id1

.ENDS nand3

.SUBCKT mos_w3800_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=3.800


.ENDS mos_w3800_l150_m1_nf1_id1

.SUBCKT mos_w1530_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=1.530


.ENDS mos_w1530_l150_m1_nf1_id0

.SUBCKT folded_inv_4 vdd vss a y

  XMP0 y a vdd vdd mos_w3800_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w1530_l150_m1_nf1_id0
  XMP1 y a vdd vdd mos_w3800_l150_m1_nf1_id1
  XMN1 y a vss vss mos_w1530_l150_m1_nf1_id0

.ENDS folded_inv_4

.SUBCKT decoder_stage_8 vdd vss y[0] y[1] y[2] y[3] y[4] y[5] y[6] y[7] y_b[0] y_b[1] y_b[2] y_b[3] y_b[4] y_b[5] y_b[6] y_b[7] predecode_0_0 predecode_0_1 predecode_1_0 predecode_1_1 predecode_2_0 predecode_2_1

  Xgate_0_0_0 vdd vss predecode_0_0 predecode_1_0 predecode_2_0 y_b[0] nand3
  Xgate_0_1_0 vdd vss predecode_0_1 predecode_1_0 predecode_2_0 y_b[1] nand3
  Xgate_0_2_0 vdd vss predecode_0_0 predecode_1_1 predecode_2_0 y_b[2] nand3
  Xgate_0_3_0 vdd vss predecode_0_1 predecode_1_1 predecode_2_0 y_b[3] nand3
  Xgate_0_4_0 vdd vss predecode_0_0 predecode_1_0 predecode_2_1 y_b[4] nand3
  Xgate_0_5_0 vdd vss predecode_0_1 predecode_1_0 predecode_2_1 y_b[5] nand3
  Xgate_0_6_0 vdd vss predecode_0_0 predecode_1_1 predecode_2_1 y_b[6] nand3
  Xgate_0_7_0 vdd vss predecode_0_1 predecode_1_1 predecode_2_1 y_b[7] nand3
  Xgate_1_0_0 vdd vss y_b[0] y[0] folded_inv_4
  Xgate_1_1_0 vdd vss y_b[1] y[1] folded_inv_4
  Xgate_1_2_0 vdd vss y_b[2] y[2] folded_inv_4
  Xgate_1_3_0 vdd vss y_b[3] y[3] folded_inv_4
  Xgate_1_4_0 vdd vss y_b[4] y[4] folded_inv_4
  Xgate_1_5_0 vdd vss y_b[5] y[5] folded_inv_4
  Xgate_1_6_0 vdd vss y_b[6] y[6] folded_inv_4
  Xgate_1_7_0 vdd vss y_b[7] y[7] folded_inv_4

.ENDS decoder_stage_8

.SUBCKT decoder_2 vdd vss y[0] y[1] y[2] y[3] y[4] y[5] y[6] y[7] y_b[0] y_b[1] y_b[2] y_b[3] y_b[4] y_b[5] y_b[6] y_b[7] predecode_0_0 predecode_0_1 predecode_1_0 predecode_1_1 predecode_2_0 predecode_2_1

  X0 vdd vss y[0] y[1] y[2] y[3] y[4] y[5] y[6] y[7] y_b[0] y_b[1] y_b[2] y_b[3] y_b[4] y_b[5] y_b[6] y_b[7] predecode_0_0 predecode_0_1 predecode_1_0 predecode_1_1 predecode_2_0 predecode_2_1 decoder_stage_8

.ENDS decoder_2

.SUBCKT mos_w2650_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=2.650


.ENDS mos_w2650_l150_m1_nf1_id1

.SUBCKT mos_w1050_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=1.050


.ENDS mos_w1050_l150_m1_nf1_id0

.SUBCKT folded_inv_5 vdd vss a y

  XMP0 y a vdd vdd mos_w2650_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w1050_l150_m1_nf1_id0
  XMP1 y a vdd vdd mos_w2650_l150_m1_nf1_id1
  XMN1 y a vss vss mos_w1050_l150_m1_nf1_id0

.ENDS folded_inv_5

.SUBCKT and2_1 vdd a b y yb vss

  X0 vdd vss a b yb nand2
  X0_1 vdd vss yb y folded_inv_5

.ENDS and2_1

.SUBCKT multi_finger_inv_14 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP8 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP9 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP10 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP11 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP12 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP13 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP14 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP15 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP16 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN3 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN4 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN5 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN6 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_14

.SUBCKT multi_finger_inv_15 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP8 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP9 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP10 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP11 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP12 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP13 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP14 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP15 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP16 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP17 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP18 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP19 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP20 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP21 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP22 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP23 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP24 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP25 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP26 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP27 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP28 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP29 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP30 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP31 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP32 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP33 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP34 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP35 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP36 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN3 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN4 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN5 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN6 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN7 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN8 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN9 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN10 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN11 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN12 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN13 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN14 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_15

.SUBCKT multi_finger_inv_16 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP8 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP9 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP10 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP11 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP12 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP13 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP14 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP15 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP16 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP17 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP18 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP19 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP20 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP21 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP22 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP23 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP24 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP25 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP26 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP27 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP28 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP29 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP30 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP31 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP32 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP33 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP34 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP35 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP36 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP37 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP38 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP39 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP40 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP41 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP42 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP43 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP44 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP45 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP46 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP47 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP48 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP49 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP50 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP51 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP52 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP53 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP54 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP55 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP56 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP57 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP58 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP59 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP60 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP61 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP62 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP63 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP64 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP65 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP66 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP67 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP68 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP69 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP70 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP71 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP72 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP73 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP74 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP75 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP76 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP77 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP78 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP79 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP80 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP81 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN3 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN4 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN5 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN6 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN7 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN8 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN9 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN10 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN11 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN12 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN13 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN14 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN15 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN16 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN17 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN18 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN19 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN20 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN21 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN22 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN23 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN24 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN25 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN26 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN27 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN28 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN29 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN30 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN31 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN32 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_16

.SUBCKT multi_finger_inv_17 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP8 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP9 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP10 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP11 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP12 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP13 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP14 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP15 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP16 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP17 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP18 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP19 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP20 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP21 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP22 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP23 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP24 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP25 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP26 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP27 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP28 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP29 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP30 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP31 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP32 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP33 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP34 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP35 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP36 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP37 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP38 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP39 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP40 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP41 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP42 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP43 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP44 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP45 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP46 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP47 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP48 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP49 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP50 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP51 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP52 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP53 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP54 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP55 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP56 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP57 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP58 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP59 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP60 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP61 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP62 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP63 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP64 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP65 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP66 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP67 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP68 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP69 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP70 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP71 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP72 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP73 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP74 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP75 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP76 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP77 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP78 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP79 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP80 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP81 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP82 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP83 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP84 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP85 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP86 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP87 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP88 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP89 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP90 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP91 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP92 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP93 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP94 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP95 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP96 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP97 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP98 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP99 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP100 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP101 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP102 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP103 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP104 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP105 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP106 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP107 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP108 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP109 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP110 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP111 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP112 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP113 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP114 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP115 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP116 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP117 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP118 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP119 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP120 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP121 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP122 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP123 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP124 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP125 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP126 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP127 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP128 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP129 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP130 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP131 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP132 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP133 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP134 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP135 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP136 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP137 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP138 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP139 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP140 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP141 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP142 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP143 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP144 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP145 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP146 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP147 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP148 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP149 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP150 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP151 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP152 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP153 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP154 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP155 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP156 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP157 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP158 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP159 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP160 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP161 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP162 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP163 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP164 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP165 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP166 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP167 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP168 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP169 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP170 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP171 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP172 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP173 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP174 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP175 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP176 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP177 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP178 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP179 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN3 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN4 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN5 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN6 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN7 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN8 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN9 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN10 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN11 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN12 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN13 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN14 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN15 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN16 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN17 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN18 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN19 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN20 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN21 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN22 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN23 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN24 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN25 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN26 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN27 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN28 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN29 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN30 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN31 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN32 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN33 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN34 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN35 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN36 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN37 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN38 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN39 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN40 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN41 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN42 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN43 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN44 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN45 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN46 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN47 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN48 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN49 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN50 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN51 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN52 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN53 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN54 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN55 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN56 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN57 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN58 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN59 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN60 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN61 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN62 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN63 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN64 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN65 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN66 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN67 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN68 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN69 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN70 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN71 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_17

.SUBCKT decoder_stage_5 vdd vss y[0] y[1] y[2] y[3] y[4] y[5] y[6] y[7] y[8] y[9] y[10] y[11] y[12] y[13] y[14] y[15] y[16] y[17] y[18] y[19] y[20] y[21] y[22] y[23] y[24] y[25] y[26] y[27] y[28] y[29] y[30] y[31] y[32] y[33] y[34] y[35] y[36] y[37] y[38] y[39] y[40] y[41] y[42] y[43] y[44] y[45] y[46] y[47] y[48] y[49] y[50] y[51] y[52] y[53] y[54] y[55] y[56] y[57] y[58] y[59] y[60] y[61] y[62] y[63] y_b[0] y_b[1] y_b[2] y_b[3] y_b[4] y_b[5] y_b[6] y_b[7] y_b[8] y_b[9] y_b[10] y_b[11] y_b[12] y_b[13] y_b[14] y_b[15] y_b[16] y_b[17] y_b[18] y_b[19] y_b[20] y_b[21] y_b[22] y_b[23] y_b[24] y_b[25] y_b[26] y_b[27] y_b[28] y_b[29] y_b[30] y_b[31] y_b[32] y_b[33] y_b[34] y_b[35] y_b[36] y_b[37] y_b[38] y_b[39] y_b[40] y_b[41] y_b[42] y_b[43] y_b[44] y_b[45] y_b[46] y_b[47] y_b[48] y_b[49] y_b[50] y_b[51] y_b[52] y_b[53] y_b[54] y_b[55] y_b[56] y_b[57] y_b[58] y_b[59] y_b[60] y_b[61] y_b[62] y_b[63] predecode_0_0 predecode_0_1 predecode_0_2 predecode_0_3 predecode_0_4 predecode_0_5 predecode_0_6 predecode_0_7 predecode_1_0 predecode_1_1 predecode_1_2 predecode_1_3 predecode_1_4 predecode_1_5 predecode_1_6 predecode_1_7

  Xgate_0_0_0 vdd predecode_0_0 predecode_1_0 x_0[0] y_b_noconn_0_0_0 vss and2_1
  Xgate_0_1_0 vdd predecode_0_1 predecode_1_0 x_0[1] y_b_noconn_0_1_0 vss and2_1
  Xgate_0_2_0 vdd predecode_0_2 predecode_1_0 x_0[2] y_b_noconn_0_2_0 vss and2_1
  Xgate_0_3_0 vdd predecode_0_3 predecode_1_0 x_0[3] y_b_noconn_0_3_0 vss and2_1
  Xgate_0_4_0 vdd predecode_0_4 predecode_1_0 x_0[4] y_b_noconn_0_4_0 vss and2_1
  Xgate_0_5_0 vdd predecode_0_5 predecode_1_0 x_0[5] y_b_noconn_0_5_0 vss and2_1
  Xgate_0_6_0 vdd predecode_0_6 predecode_1_0 x_0[6] y_b_noconn_0_6_0 vss and2_1
  Xgate_0_7_0 vdd predecode_0_7 predecode_1_0 x_0[7] y_b_noconn_0_7_0 vss and2_1
  Xgate_0_8_0 vdd predecode_0_0 predecode_1_1 x_0[8] y_b_noconn_0_8_0 vss and2_1
  Xgate_0_9_0 vdd predecode_0_1 predecode_1_1 x_0[9] y_b_noconn_0_9_0 vss and2_1
  Xgate_0_10_0 vdd predecode_0_2 predecode_1_1 x_0[10] y_b_noconn_0_10_0 vss and2_1
  Xgate_0_11_0 vdd predecode_0_3 predecode_1_1 x_0[11] y_b_noconn_0_11_0 vss and2_1
  Xgate_0_12_0 vdd predecode_0_4 predecode_1_1 x_0[12] y_b_noconn_0_12_0 vss and2_1
  Xgate_0_13_0 vdd predecode_0_5 predecode_1_1 x_0[13] y_b_noconn_0_13_0 vss and2_1
  Xgate_0_14_0 vdd predecode_0_6 predecode_1_1 x_0[14] y_b_noconn_0_14_0 vss and2_1
  Xgate_0_15_0 vdd predecode_0_7 predecode_1_1 x_0[15] y_b_noconn_0_15_0 vss and2_1
  Xgate_0_16_0 vdd predecode_0_0 predecode_1_2 x_0[16] y_b_noconn_0_16_0 vss and2_1
  Xgate_0_17_0 vdd predecode_0_1 predecode_1_2 x_0[17] y_b_noconn_0_17_0 vss and2_1
  Xgate_0_18_0 vdd predecode_0_2 predecode_1_2 x_0[18] y_b_noconn_0_18_0 vss and2_1
  Xgate_0_19_0 vdd predecode_0_3 predecode_1_2 x_0[19] y_b_noconn_0_19_0 vss and2_1
  Xgate_0_20_0 vdd predecode_0_4 predecode_1_2 x_0[20] y_b_noconn_0_20_0 vss and2_1
  Xgate_0_21_0 vdd predecode_0_5 predecode_1_2 x_0[21] y_b_noconn_0_21_0 vss and2_1
  Xgate_0_22_0 vdd predecode_0_6 predecode_1_2 x_0[22] y_b_noconn_0_22_0 vss and2_1
  Xgate_0_23_0 vdd predecode_0_7 predecode_1_2 x_0[23] y_b_noconn_0_23_0 vss and2_1
  Xgate_0_24_0 vdd predecode_0_0 predecode_1_3 x_0[24] y_b_noconn_0_24_0 vss and2_1
  Xgate_0_25_0 vdd predecode_0_1 predecode_1_3 x_0[25] y_b_noconn_0_25_0 vss and2_1
  Xgate_0_26_0 vdd predecode_0_2 predecode_1_3 x_0[26] y_b_noconn_0_26_0 vss and2_1
  Xgate_0_27_0 vdd predecode_0_3 predecode_1_3 x_0[27] y_b_noconn_0_27_0 vss and2_1
  Xgate_0_28_0 vdd predecode_0_4 predecode_1_3 x_0[28] y_b_noconn_0_28_0 vss and2_1
  Xgate_0_29_0 vdd predecode_0_5 predecode_1_3 x_0[29] y_b_noconn_0_29_0 vss and2_1
  Xgate_0_30_0 vdd predecode_0_6 predecode_1_3 x_0[30] y_b_noconn_0_30_0 vss and2_1
  Xgate_0_31_0 vdd predecode_0_7 predecode_1_3 x_0[31] y_b_noconn_0_31_0 vss and2_1
  Xgate_0_32_0 vdd predecode_0_0 predecode_1_4 x_0[32] y_b_noconn_0_32_0 vss and2_1
  Xgate_0_33_0 vdd predecode_0_1 predecode_1_4 x_0[33] y_b_noconn_0_33_0 vss and2_1
  Xgate_0_34_0 vdd predecode_0_2 predecode_1_4 x_0[34] y_b_noconn_0_34_0 vss and2_1
  Xgate_0_35_0 vdd predecode_0_3 predecode_1_4 x_0[35] y_b_noconn_0_35_0 vss and2_1
  Xgate_0_36_0 vdd predecode_0_4 predecode_1_4 x_0[36] y_b_noconn_0_36_0 vss and2_1
  Xgate_0_37_0 vdd predecode_0_5 predecode_1_4 x_0[37] y_b_noconn_0_37_0 vss and2_1
  Xgate_0_38_0 vdd predecode_0_6 predecode_1_4 x_0[38] y_b_noconn_0_38_0 vss and2_1
  Xgate_0_39_0 vdd predecode_0_7 predecode_1_4 x_0[39] y_b_noconn_0_39_0 vss and2_1
  Xgate_0_40_0 vdd predecode_0_0 predecode_1_5 x_0[40] y_b_noconn_0_40_0 vss and2_1
  Xgate_0_41_0 vdd predecode_0_1 predecode_1_5 x_0[41] y_b_noconn_0_41_0 vss and2_1
  Xgate_0_42_0 vdd predecode_0_2 predecode_1_5 x_0[42] y_b_noconn_0_42_0 vss and2_1
  Xgate_0_43_0 vdd predecode_0_3 predecode_1_5 x_0[43] y_b_noconn_0_43_0 vss and2_1
  Xgate_0_44_0 vdd predecode_0_4 predecode_1_5 x_0[44] y_b_noconn_0_44_0 vss and2_1
  Xgate_0_45_0 vdd predecode_0_5 predecode_1_5 x_0[45] y_b_noconn_0_45_0 vss and2_1
  Xgate_0_46_0 vdd predecode_0_6 predecode_1_5 x_0[46] y_b_noconn_0_46_0 vss and2_1
  Xgate_0_47_0 vdd predecode_0_7 predecode_1_5 x_0[47] y_b_noconn_0_47_0 vss and2_1
  Xgate_0_48_0 vdd predecode_0_0 predecode_1_6 x_0[48] y_b_noconn_0_48_0 vss and2_1
  Xgate_0_49_0 vdd predecode_0_1 predecode_1_6 x_0[49] y_b_noconn_0_49_0 vss and2_1
  Xgate_0_50_0 vdd predecode_0_2 predecode_1_6 x_0[50] y_b_noconn_0_50_0 vss and2_1
  Xgate_0_51_0 vdd predecode_0_3 predecode_1_6 x_0[51] y_b_noconn_0_51_0 vss and2_1
  Xgate_0_52_0 vdd predecode_0_4 predecode_1_6 x_0[52] y_b_noconn_0_52_0 vss and2_1
  Xgate_0_53_0 vdd predecode_0_5 predecode_1_6 x_0[53] y_b_noconn_0_53_0 vss and2_1
  Xgate_0_54_0 vdd predecode_0_6 predecode_1_6 x_0[54] y_b_noconn_0_54_0 vss and2_1
  Xgate_0_55_0 vdd predecode_0_7 predecode_1_6 x_0[55] y_b_noconn_0_55_0 vss and2_1
  Xgate_0_56_0 vdd predecode_0_0 predecode_1_7 x_0[56] y_b_noconn_0_56_0 vss and2_1
  Xgate_0_57_0 vdd predecode_0_1 predecode_1_7 x_0[57] y_b_noconn_0_57_0 vss and2_1
  Xgate_0_58_0 vdd predecode_0_2 predecode_1_7 x_0[58] y_b_noconn_0_58_0 vss and2_1
  Xgate_0_59_0 vdd predecode_0_3 predecode_1_7 x_0[59] y_b_noconn_0_59_0 vss and2_1
  Xgate_0_60_0 vdd predecode_0_4 predecode_1_7 x_0[60] y_b_noconn_0_60_0 vss and2_1
  Xgate_0_61_0 vdd predecode_0_5 predecode_1_7 x_0[61] y_b_noconn_0_61_0 vss and2_1
  Xgate_0_62_0 vdd predecode_0_6 predecode_1_7 x_0[62] y_b_noconn_0_62_0 vss and2_1
  Xgate_0_63_0 vdd predecode_0_7 predecode_1_7 x_0[63] y_b_noconn_0_63_0 vss and2_1
  Xgate_1_0_0 vdd vss x_0[0] x_1[0] multi_finger_inv_14
  Xgate_1_1_0 vdd vss x_0[1] x_1[1] multi_finger_inv_14
  Xgate_1_2_0 vdd vss x_0[2] x_1[2] multi_finger_inv_14
  Xgate_1_3_0 vdd vss x_0[3] x_1[3] multi_finger_inv_14
  Xgate_1_4_0 vdd vss x_0[4] x_1[4] multi_finger_inv_14
  Xgate_1_5_0 vdd vss x_0[5] x_1[5] multi_finger_inv_14
  Xgate_1_6_0 vdd vss x_0[6] x_1[6] multi_finger_inv_14
  Xgate_1_7_0 vdd vss x_0[7] x_1[7] multi_finger_inv_14
  Xgate_1_8_0 vdd vss x_0[8] x_1[8] multi_finger_inv_14
  Xgate_1_9_0 vdd vss x_0[9] x_1[9] multi_finger_inv_14
  Xgate_1_10_0 vdd vss x_0[10] x_1[10] multi_finger_inv_14
  Xgate_1_11_0 vdd vss x_0[11] x_1[11] multi_finger_inv_14
  Xgate_1_12_0 vdd vss x_0[12] x_1[12] multi_finger_inv_14
  Xgate_1_13_0 vdd vss x_0[13] x_1[13] multi_finger_inv_14
  Xgate_1_14_0 vdd vss x_0[14] x_1[14] multi_finger_inv_14
  Xgate_1_15_0 vdd vss x_0[15] x_1[15] multi_finger_inv_14
  Xgate_1_16_0 vdd vss x_0[16] x_1[16] multi_finger_inv_14
  Xgate_1_17_0 vdd vss x_0[17] x_1[17] multi_finger_inv_14
  Xgate_1_18_0 vdd vss x_0[18] x_1[18] multi_finger_inv_14
  Xgate_1_19_0 vdd vss x_0[19] x_1[19] multi_finger_inv_14
  Xgate_1_20_0 vdd vss x_0[20] x_1[20] multi_finger_inv_14
  Xgate_1_21_0 vdd vss x_0[21] x_1[21] multi_finger_inv_14
  Xgate_1_22_0 vdd vss x_0[22] x_1[22] multi_finger_inv_14
  Xgate_1_23_0 vdd vss x_0[23] x_1[23] multi_finger_inv_14
  Xgate_1_24_0 vdd vss x_0[24] x_1[24] multi_finger_inv_14
  Xgate_1_25_0 vdd vss x_0[25] x_1[25] multi_finger_inv_14
  Xgate_1_26_0 vdd vss x_0[26] x_1[26] multi_finger_inv_14
  Xgate_1_27_0 vdd vss x_0[27] x_1[27] multi_finger_inv_14
  Xgate_1_28_0 vdd vss x_0[28] x_1[28] multi_finger_inv_14
  Xgate_1_29_0 vdd vss x_0[29] x_1[29] multi_finger_inv_14
  Xgate_1_30_0 vdd vss x_0[30] x_1[30] multi_finger_inv_14
  Xgate_1_31_0 vdd vss x_0[31] x_1[31] multi_finger_inv_14
  Xgate_1_32_0 vdd vss x_0[32] x_1[32] multi_finger_inv_14
  Xgate_1_33_0 vdd vss x_0[33] x_1[33] multi_finger_inv_14
  Xgate_1_34_0 vdd vss x_0[34] x_1[34] multi_finger_inv_14
  Xgate_1_35_0 vdd vss x_0[35] x_1[35] multi_finger_inv_14
  Xgate_1_36_0 vdd vss x_0[36] x_1[36] multi_finger_inv_14
  Xgate_1_37_0 vdd vss x_0[37] x_1[37] multi_finger_inv_14
  Xgate_1_38_0 vdd vss x_0[38] x_1[38] multi_finger_inv_14
  Xgate_1_39_0 vdd vss x_0[39] x_1[39] multi_finger_inv_14
  Xgate_1_40_0 vdd vss x_0[40] x_1[40] multi_finger_inv_14
  Xgate_1_41_0 vdd vss x_0[41] x_1[41] multi_finger_inv_14
  Xgate_1_42_0 vdd vss x_0[42] x_1[42] multi_finger_inv_14
  Xgate_1_43_0 vdd vss x_0[43] x_1[43] multi_finger_inv_14
  Xgate_1_44_0 vdd vss x_0[44] x_1[44] multi_finger_inv_14
  Xgate_1_45_0 vdd vss x_0[45] x_1[45] multi_finger_inv_14
  Xgate_1_46_0 vdd vss x_0[46] x_1[46] multi_finger_inv_14
  Xgate_1_47_0 vdd vss x_0[47] x_1[47] multi_finger_inv_14
  Xgate_1_48_0 vdd vss x_0[48] x_1[48] multi_finger_inv_14
  Xgate_1_49_0 vdd vss x_0[49] x_1[49] multi_finger_inv_14
  Xgate_1_50_0 vdd vss x_0[50] x_1[50] multi_finger_inv_14
  Xgate_1_51_0 vdd vss x_0[51] x_1[51] multi_finger_inv_14
  Xgate_1_52_0 vdd vss x_0[52] x_1[52] multi_finger_inv_14
  Xgate_1_53_0 vdd vss x_0[53] x_1[53] multi_finger_inv_14
  Xgate_1_54_0 vdd vss x_0[54] x_1[54] multi_finger_inv_14
  Xgate_1_55_0 vdd vss x_0[55] x_1[55] multi_finger_inv_14
  Xgate_1_56_0 vdd vss x_0[56] x_1[56] multi_finger_inv_14
  Xgate_1_57_0 vdd vss x_0[57] x_1[57] multi_finger_inv_14
  Xgate_1_58_0 vdd vss x_0[58] x_1[58] multi_finger_inv_14
  Xgate_1_59_0 vdd vss x_0[59] x_1[59] multi_finger_inv_14
  Xgate_1_60_0 vdd vss x_0[60] x_1[60] multi_finger_inv_14
  Xgate_1_61_0 vdd vss x_0[61] x_1[61] multi_finger_inv_14
  Xgate_1_62_0 vdd vss x_0[62] x_1[62] multi_finger_inv_14
  Xgate_1_63_0 vdd vss x_0[63] x_1[63] multi_finger_inv_14
  Xgate_2_0_0 vdd vss x_1[0] x_2[0] multi_finger_inv_15
  Xgate_2_1_0 vdd vss x_1[1] x_2[1] multi_finger_inv_15
  Xgate_2_2_0 vdd vss x_1[2] x_2[2] multi_finger_inv_15
  Xgate_2_3_0 vdd vss x_1[3] x_2[3] multi_finger_inv_15
  Xgate_2_4_0 vdd vss x_1[4] x_2[4] multi_finger_inv_15
  Xgate_2_5_0 vdd vss x_1[5] x_2[5] multi_finger_inv_15
  Xgate_2_6_0 vdd vss x_1[6] x_2[6] multi_finger_inv_15
  Xgate_2_7_0 vdd vss x_1[7] x_2[7] multi_finger_inv_15
  Xgate_2_8_0 vdd vss x_1[8] x_2[8] multi_finger_inv_15
  Xgate_2_9_0 vdd vss x_1[9] x_2[9] multi_finger_inv_15
  Xgate_2_10_0 vdd vss x_1[10] x_2[10] multi_finger_inv_15
  Xgate_2_11_0 vdd vss x_1[11] x_2[11] multi_finger_inv_15
  Xgate_2_12_0 vdd vss x_1[12] x_2[12] multi_finger_inv_15
  Xgate_2_13_0 vdd vss x_1[13] x_2[13] multi_finger_inv_15
  Xgate_2_14_0 vdd vss x_1[14] x_2[14] multi_finger_inv_15
  Xgate_2_15_0 vdd vss x_1[15] x_2[15] multi_finger_inv_15
  Xgate_2_16_0 vdd vss x_1[16] x_2[16] multi_finger_inv_15
  Xgate_2_17_0 vdd vss x_1[17] x_2[17] multi_finger_inv_15
  Xgate_2_18_0 vdd vss x_1[18] x_2[18] multi_finger_inv_15
  Xgate_2_19_0 vdd vss x_1[19] x_2[19] multi_finger_inv_15
  Xgate_2_20_0 vdd vss x_1[20] x_2[20] multi_finger_inv_15
  Xgate_2_21_0 vdd vss x_1[21] x_2[21] multi_finger_inv_15
  Xgate_2_22_0 vdd vss x_1[22] x_2[22] multi_finger_inv_15
  Xgate_2_23_0 vdd vss x_1[23] x_2[23] multi_finger_inv_15
  Xgate_2_24_0 vdd vss x_1[24] x_2[24] multi_finger_inv_15
  Xgate_2_25_0 vdd vss x_1[25] x_2[25] multi_finger_inv_15
  Xgate_2_26_0 vdd vss x_1[26] x_2[26] multi_finger_inv_15
  Xgate_2_27_0 vdd vss x_1[27] x_2[27] multi_finger_inv_15
  Xgate_2_28_0 vdd vss x_1[28] x_2[28] multi_finger_inv_15
  Xgate_2_29_0 vdd vss x_1[29] x_2[29] multi_finger_inv_15
  Xgate_2_30_0 vdd vss x_1[30] x_2[30] multi_finger_inv_15
  Xgate_2_31_0 vdd vss x_1[31] x_2[31] multi_finger_inv_15
  Xgate_2_32_0 vdd vss x_1[32] x_2[32] multi_finger_inv_15
  Xgate_2_33_0 vdd vss x_1[33] x_2[33] multi_finger_inv_15
  Xgate_2_34_0 vdd vss x_1[34] x_2[34] multi_finger_inv_15
  Xgate_2_35_0 vdd vss x_1[35] x_2[35] multi_finger_inv_15
  Xgate_2_36_0 vdd vss x_1[36] x_2[36] multi_finger_inv_15
  Xgate_2_37_0 vdd vss x_1[37] x_2[37] multi_finger_inv_15
  Xgate_2_38_0 vdd vss x_1[38] x_2[38] multi_finger_inv_15
  Xgate_2_39_0 vdd vss x_1[39] x_2[39] multi_finger_inv_15
  Xgate_2_40_0 vdd vss x_1[40] x_2[40] multi_finger_inv_15
  Xgate_2_41_0 vdd vss x_1[41] x_2[41] multi_finger_inv_15
  Xgate_2_42_0 vdd vss x_1[42] x_2[42] multi_finger_inv_15
  Xgate_2_43_0 vdd vss x_1[43] x_2[43] multi_finger_inv_15
  Xgate_2_44_0 vdd vss x_1[44] x_2[44] multi_finger_inv_15
  Xgate_2_45_0 vdd vss x_1[45] x_2[45] multi_finger_inv_15
  Xgate_2_46_0 vdd vss x_1[46] x_2[46] multi_finger_inv_15
  Xgate_2_47_0 vdd vss x_1[47] x_2[47] multi_finger_inv_15
  Xgate_2_48_0 vdd vss x_1[48] x_2[48] multi_finger_inv_15
  Xgate_2_49_0 vdd vss x_1[49] x_2[49] multi_finger_inv_15
  Xgate_2_50_0 vdd vss x_1[50] x_2[50] multi_finger_inv_15
  Xgate_2_51_0 vdd vss x_1[51] x_2[51] multi_finger_inv_15
  Xgate_2_52_0 vdd vss x_1[52] x_2[52] multi_finger_inv_15
  Xgate_2_53_0 vdd vss x_1[53] x_2[53] multi_finger_inv_15
  Xgate_2_54_0 vdd vss x_1[54] x_2[54] multi_finger_inv_15
  Xgate_2_55_0 vdd vss x_1[55] x_2[55] multi_finger_inv_15
  Xgate_2_56_0 vdd vss x_1[56] x_2[56] multi_finger_inv_15
  Xgate_2_57_0 vdd vss x_1[57] x_2[57] multi_finger_inv_15
  Xgate_2_58_0 vdd vss x_1[58] x_2[58] multi_finger_inv_15
  Xgate_2_59_0 vdd vss x_1[59] x_2[59] multi_finger_inv_15
  Xgate_2_60_0 vdd vss x_1[60] x_2[60] multi_finger_inv_15
  Xgate_2_61_0 vdd vss x_1[61] x_2[61] multi_finger_inv_15
  Xgate_2_62_0 vdd vss x_1[62] x_2[62] multi_finger_inv_15
  Xgate_2_63_0 vdd vss x_1[63] x_2[63] multi_finger_inv_15
  Xgate_3_0_0 vdd vss x_2[0] y_b[0] multi_finger_inv_16
  Xgate_3_1_0 vdd vss x_2[1] y_b[1] multi_finger_inv_16
  Xgate_3_2_0 vdd vss x_2[2] y_b[2] multi_finger_inv_16
  Xgate_3_3_0 vdd vss x_2[3] y_b[3] multi_finger_inv_16
  Xgate_3_4_0 vdd vss x_2[4] y_b[4] multi_finger_inv_16
  Xgate_3_5_0 vdd vss x_2[5] y_b[5] multi_finger_inv_16
  Xgate_3_6_0 vdd vss x_2[6] y_b[6] multi_finger_inv_16
  Xgate_3_7_0 vdd vss x_2[7] y_b[7] multi_finger_inv_16
  Xgate_3_8_0 vdd vss x_2[8] y_b[8] multi_finger_inv_16
  Xgate_3_9_0 vdd vss x_2[9] y_b[9] multi_finger_inv_16
  Xgate_3_10_0 vdd vss x_2[10] y_b[10] multi_finger_inv_16
  Xgate_3_11_0 vdd vss x_2[11] y_b[11] multi_finger_inv_16
  Xgate_3_12_0 vdd vss x_2[12] y_b[12] multi_finger_inv_16
  Xgate_3_13_0 vdd vss x_2[13] y_b[13] multi_finger_inv_16
  Xgate_3_14_0 vdd vss x_2[14] y_b[14] multi_finger_inv_16
  Xgate_3_15_0 vdd vss x_2[15] y_b[15] multi_finger_inv_16
  Xgate_3_16_0 vdd vss x_2[16] y_b[16] multi_finger_inv_16
  Xgate_3_17_0 vdd vss x_2[17] y_b[17] multi_finger_inv_16
  Xgate_3_18_0 vdd vss x_2[18] y_b[18] multi_finger_inv_16
  Xgate_3_19_0 vdd vss x_2[19] y_b[19] multi_finger_inv_16
  Xgate_3_20_0 vdd vss x_2[20] y_b[20] multi_finger_inv_16
  Xgate_3_21_0 vdd vss x_2[21] y_b[21] multi_finger_inv_16
  Xgate_3_22_0 vdd vss x_2[22] y_b[22] multi_finger_inv_16
  Xgate_3_23_0 vdd vss x_2[23] y_b[23] multi_finger_inv_16
  Xgate_3_24_0 vdd vss x_2[24] y_b[24] multi_finger_inv_16
  Xgate_3_25_0 vdd vss x_2[25] y_b[25] multi_finger_inv_16
  Xgate_3_26_0 vdd vss x_2[26] y_b[26] multi_finger_inv_16
  Xgate_3_27_0 vdd vss x_2[27] y_b[27] multi_finger_inv_16
  Xgate_3_28_0 vdd vss x_2[28] y_b[28] multi_finger_inv_16
  Xgate_3_29_0 vdd vss x_2[29] y_b[29] multi_finger_inv_16
  Xgate_3_30_0 vdd vss x_2[30] y_b[30] multi_finger_inv_16
  Xgate_3_31_0 vdd vss x_2[31] y_b[31] multi_finger_inv_16
  Xgate_3_32_0 vdd vss x_2[32] y_b[32] multi_finger_inv_16
  Xgate_3_33_0 vdd vss x_2[33] y_b[33] multi_finger_inv_16
  Xgate_3_34_0 vdd vss x_2[34] y_b[34] multi_finger_inv_16
  Xgate_3_35_0 vdd vss x_2[35] y_b[35] multi_finger_inv_16
  Xgate_3_36_0 vdd vss x_2[36] y_b[36] multi_finger_inv_16
  Xgate_3_37_0 vdd vss x_2[37] y_b[37] multi_finger_inv_16
  Xgate_3_38_0 vdd vss x_2[38] y_b[38] multi_finger_inv_16
  Xgate_3_39_0 vdd vss x_2[39] y_b[39] multi_finger_inv_16
  Xgate_3_40_0 vdd vss x_2[40] y_b[40] multi_finger_inv_16
  Xgate_3_41_0 vdd vss x_2[41] y_b[41] multi_finger_inv_16
  Xgate_3_42_0 vdd vss x_2[42] y_b[42] multi_finger_inv_16
  Xgate_3_43_0 vdd vss x_2[43] y_b[43] multi_finger_inv_16
  Xgate_3_44_0 vdd vss x_2[44] y_b[44] multi_finger_inv_16
  Xgate_3_45_0 vdd vss x_2[45] y_b[45] multi_finger_inv_16
  Xgate_3_46_0 vdd vss x_2[46] y_b[46] multi_finger_inv_16
  Xgate_3_47_0 vdd vss x_2[47] y_b[47] multi_finger_inv_16
  Xgate_3_48_0 vdd vss x_2[48] y_b[48] multi_finger_inv_16
  Xgate_3_49_0 vdd vss x_2[49] y_b[49] multi_finger_inv_16
  Xgate_3_50_0 vdd vss x_2[50] y_b[50] multi_finger_inv_16
  Xgate_3_51_0 vdd vss x_2[51] y_b[51] multi_finger_inv_16
  Xgate_3_52_0 vdd vss x_2[52] y_b[52] multi_finger_inv_16
  Xgate_3_53_0 vdd vss x_2[53] y_b[53] multi_finger_inv_16
  Xgate_3_54_0 vdd vss x_2[54] y_b[54] multi_finger_inv_16
  Xgate_3_55_0 vdd vss x_2[55] y_b[55] multi_finger_inv_16
  Xgate_3_56_0 vdd vss x_2[56] y_b[56] multi_finger_inv_16
  Xgate_3_57_0 vdd vss x_2[57] y_b[57] multi_finger_inv_16
  Xgate_3_58_0 vdd vss x_2[58] y_b[58] multi_finger_inv_16
  Xgate_3_59_0 vdd vss x_2[59] y_b[59] multi_finger_inv_16
  Xgate_3_60_0 vdd vss x_2[60] y_b[60] multi_finger_inv_16
  Xgate_3_61_0 vdd vss x_2[61] y_b[61] multi_finger_inv_16
  Xgate_3_62_0 vdd vss x_2[62] y_b[62] multi_finger_inv_16
  Xgate_3_63_0 vdd vss x_2[63] y_b[63] multi_finger_inv_16
  Xgate_4_0_0 vdd vss y_b[0] y[0] multi_finger_inv_17
  Xgate_4_1_0 vdd vss y_b[1] y[1] multi_finger_inv_17
  Xgate_4_2_0 vdd vss y_b[2] y[2] multi_finger_inv_17
  Xgate_4_3_0 vdd vss y_b[3] y[3] multi_finger_inv_17
  Xgate_4_4_0 vdd vss y_b[4] y[4] multi_finger_inv_17
  Xgate_4_5_0 vdd vss y_b[5] y[5] multi_finger_inv_17
  Xgate_4_6_0 vdd vss y_b[6] y[6] multi_finger_inv_17
  Xgate_4_7_0 vdd vss y_b[7] y[7] multi_finger_inv_17
  Xgate_4_8_0 vdd vss y_b[8] y[8] multi_finger_inv_17
  Xgate_4_9_0 vdd vss y_b[9] y[9] multi_finger_inv_17
  Xgate_4_10_0 vdd vss y_b[10] y[10] multi_finger_inv_17
  Xgate_4_11_0 vdd vss y_b[11] y[11] multi_finger_inv_17
  Xgate_4_12_0 vdd vss y_b[12] y[12] multi_finger_inv_17
  Xgate_4_13_0 vdd vss y_b[13] y[13] multi_finger_inv_17
  Xgate_4_14_0 vdd vss y_b[14] y[14] multi_finger_inv_17
  Xgate_4_15_0 vdd vss y_b[15] y[15] multi_finger_inv_17
  Xgate_4_16_0 vdd vss y_b[16] y[16] multi_finger_inv_17
  Xgate_4_17_0 vdd vss y_b[17] y[17] multi_finger_inv_17
  Xgate_4_18_0 vdd vss y_b[18] y[18] multi_finger_inv_17
  Xgate_4_19_0 vdd vss y_b[19] y[19] multi_finger_inv_17
  Xgate_4_20_0 vdd vss y_b[20] y[20] multi_finger_inv_17
  Xgate_4_21_0 vdd vss y_b[21] y[21] multi_finger_inv_17
  Xgate_4_22_0 vdd vss y_b[22] y[22] multi_finger_inv_17
  Xgate_4_23_0 vdd vss y_b[23] y[23] multi_finger_inv_17
  Xgate_4_24_0 vdd vss y_b[24] y[24] multi_finger_inv_17
  Xgate_4_25_0 vdd vss y_b[25] y[25] multi_finger_inv_17
  Xgate_4_26_0 vdd vss y_b[26] y[26] multi_finger_inv_17
  Xgate_4_27_0 vdd vss y_b[27] y[27] multi_finger_inv_17
  Xgate_4_28_0 vdd vss y_b[28] y[28] multi_finger_inv_17
  Xgate_4_29_0 vdd vss y_b[29] y[29] multi_finger_inv_17
  Xgate_4_30_0 vdd vss y_b[30] y[30] multi_finger_inv_17
  Xgate_4_31_0 vdd vss y_b[31] y[31] multi_finger_inv_17
  Xgate_4_32_0 vdd vss y_b[32] y[32] multi_finger_inv_17
  Xgate_4_33_0 vdd vss y_b[33] y[33] multi_finger_inv_17
  Xgate_4_34_0 vdd vss y_b[34] y[34] multi_finger_inv_17
  Xgate_4_35_0 vdd vss y_b[35] y[35] multi_finger_inv_17
  Xgate_4_36_0 vdd vss y_b[36] y[36] multi_finger_inv_17
  Xgate_4_37_0 vdd vss y_b[37] y[37] multi_finger_inv_17
  Xgate_4_38_0 vdd vss y_b[38] y[38] multi_finger_inv_17
  Xgate_4_39_0 vdd vss y_b[39] y[39] multi_finger_inv_17
  Xgate_4_40_0 vdd vss y_b[40] y[40] multi_finger_inv_17
  Xgate_4_41_0 vdd vss y_b[41] y[41] multi_finger_inv_17
  Xgate_4_42_0 vdd vss y_b[42] y[42] multi_finger_inv_17
  Xgate_4_43_0 vdd vss y_b[43] y[43] multi_finger_inv_17
  Xgate_4_44_0 vdd vss y_b[44] y[44] multi_finger_inv_17
  Xgate_4_45_0 vdd vss y_b[45] y[45] multi_finger_inv_17
  Xgate_4_46_0 vdd vss y_b[46] y[46] multi_finger_inv_17
  Xgate_4_47_0 vdd vss y_b[47] y[47] multi_finger_inv_17
  Xgate_4_48_0 vdd vss y_b[48] y[48] multi_finger_inv_17
  Xgate_4_49_0 vdd vss y_b[49] y[49] multi_finger_inv_17
  Xgate_4_50_0 vdd vss y_b[50] y[50] multi_finger_inv_17
  Xgate_4_51_0 vdd vss y_b[51] y[51] multi_finger_inv_17
  Xgate_4_52_0 vdd vss y_b[52] y[52] multi_finger_inv_17
  Xgate_4_53_0 vdd vss y_b[53] y[53] multi_finger_inv_17
  Xgate_4_54_0 vdd vss y_b[54] y[54] multi_finger_inv_17
  Xgate_4_55_0 vdd vss y_b[55] y[55] multi_finger_inv_17
  Xgate_4_56_0 vdd vss y_b[56] y[56] multi_finger_inv_17
  Xgate_4_57_0 vdd vss y_b[57] y[57] multi_finger_inv_17
  Xgate_4_58_0 vdd vss y_b[58] y[58] multi_finger_inv_17
  Xgate_4_59_0 vdd vss y_b[59] y[59] multi_finger_inv_17
  Xgate_4_60_0 vdd vss y_b[60] y[60] multi_finger_inv_17
  Xgate_4_61_0 vdd vss y_b[61] y[61] multi_finger_inv_17
  Xgate_4_62_0 vdd vss y_b[62] y[62] multi_finger_inv_17
  Xgate_4_63_0 vdd vss y_b[63] y[63] multi_finger_inv_17

.ENDS decoder_stage_5

.SUBCKT decoder vdd vss y[0] y[1] y[2] y[3] y[4] y[5] y[6] y[7] y[8] y[9] y[10] y[11] y[12] y[13] y[14] y[15] y[16] y[17] y[18] y[19] y[20] y[21] y[22] y[23] y[24] y[25] y[26] y[27] y[28] y[29] y[30] y[31] y[32] y[33] y[34] y[35] y[36] y[37] y[38] y[39] y[40] y[41] y[42] y[43] y[44] y[45] y[46] y[47] y[48] y[49] y[50] y[51] y[52] y[53] y[54] y[55] y[56] y[57] y[58] y[59] y[60] y[61] y[62] y[63] y_b[0] y_b[1] y_b[2] y_b[3] y_b[4] y_b[5] y_b[6] y_b[7] y_b[8] y_b[9] y_b[10] y_b[11] y_b[12] y_b[13] y_b[14] y_b[15] y_b[16] y_b[17] y_b[18] y_b[19] y_b[20] y_b[21] y_b[22] y_b[23] y_b[24] y_b[25] y_b[26] y_b[27] y_b[28] y_b[29] y_b[30] y_b[31] y_b[32] y_b[33] y_b[34] y_b[35] y_b[36] y_b[37] y_b[38] y_b[39] y_b[40] y_b[41] y_b[42] y_b[43] y_b[44] y_b[45] y_b[46] y_b[47] y_b[48] y_b[49] y_b[50] y_b[51] y_b[52] y_b[53] y_b[54] y_b[55] y_b[56] y_b[57] y_b[58] y_b[59] y_b[60] y_b[61] y_b[62] y_b[63] predecode_0_0 predecode_0_1 predecode_1_0 predecode_1_1 predecode_2_0 predecode_2_1 predecode_3_0 predecode_3_1 predecode_4_0 predecode_4_1 predecode_5_0 predecode_5_1

  X0 vdd vss child_conn_0[0] child_conn_0[1] child_conn_0[2] child_conn_0[3] child_conn_0[4] child_conn_0[5] child_conn_0[6] child_conn_0[7] child_noconn_0[0] child_noconn_0[1] child_noconn_0[2] child_noconn_0[3] child_noconn_0[4] child_noconn_0[5] child_noconn_0[6] child_noconn_0[7] predecode_0_0 predecode_0_1 predecode_1_0 predecode_1_1 predecode_2_0 predecode_2_1 decoder_2
  X0_1 vdd vss child_conn_1[0] child_conn_1[1] child_conn_1[2] child_conn_1[3] child_conn_1[4] child_conn_1[5] child_conn_1[6] child_conn_1[7] child_noconn_1[0] child_noconn_1[1] child_noconn_1[2] child_noconn_1[3] child_noconn_1[4] child_noconn_1[5] child_noconn_1[6] child_noconn_1[7] predecode_3_0 predecode_3_1 predecode_4_0 predecode_4_1 predecode_5_0 predecode_5_1 decoder_2
  X0_2 vdd vss y[0] y[1] y[2] y[3] y[4] y[5] y[6] y[7] y[8] y[9] y[10] y[11] y[12] y[13] y[14] y[15] y[16] y[17] y[18] y[19] y[20] y[21] y[22] y[23] y[24] y[25] y[26] y[27] y[28] y[29] y[30] y[31] y[32] y[33] y[34] y[35] y[36] y[37] y[38] y[39] y[40] y[41] y[42] y[43] y[44] y[45] y[46] y[47] y[48] y[49] y[50] y[51] y[52] y[53] y[54] y[55] y[56] y[57] y[58] y[59] y[60] y[61] y[62] y[63] y_b[0] y_b[1] y_b[2] y_b[3] y_b[4] y_b[5] y_b[6] y_b[7] y_b[8] y_b[9] y_b[10] y_b[11] y_b[12] y_b[13] y_b[14] y_b[15] y_b[16] y_b[17] y_b[18] y_b[19] y_b[20] y_b[21] y_b[22] y_b[23] y_b[24] y_b[25] y_b[26] y_b[27] y_b[28] y_b[29] y_b[30] y_b[31] y_b[32] y_b[33] y_b[34] y_b[35] y_b[36] y_b[37] y_b[38] y_b[39] y_b[40] y_b[41] y_b[42] y_b[43] y_b[44] y_b[45] y_b[46] y_b[47] y_b[48] y_b[49] y_b[50] y_b[51] y_b[52] y_b[53] y_b[54] y_b[55] y_b[56] y_b[57] y_b[58] y_b[59] y_b[60] y_b[61] y_b[62] y_b[63] child_conn_0[0] child_conn_0[1] child_conn_0[2] child_conn_0[3] child_conn_0[4] child_conn_0[5] child_conn_0[6] child_conn_0[7] child_conn_1[0] child_conn_1[1] child_conn_1[2] child_conn_1[3] child_conn_1[4] child_conn_1[5] child_conn_1[6] child_conn_1[7] decoder_stage_5

.ENDS decoder

.SUBCKT nand2_1 vdd vss a b y

  Xn1 x a vss vss mos_w2000_l150_m1_nf1_id0
  Xn2 y b x vss mos_w2000_l150_m1_nf1_id0
  Xp1 y a vdd vdd mos_w2500_l150_m1_nf1_id1
  Xp2 y b vdd vdd mos_w2500_l150_m1_nf1_id1

.ENDS nand2_1

.SUBCKT multi_finger_inv_18 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP8 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN3 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_18

.SUBCKT multi_finger_inv_19 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_19

.SUBCKT multi_finger_inv_20 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP8 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP9 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP10 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP11 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP12 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN3 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN4 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_20

.SUBCKT multi_finger_inv_21 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP8 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP9 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP10 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP11 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP12 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP13 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP14 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP15 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP16 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP17 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP18 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP19 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP20 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP21 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP22 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP23 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP24 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP25 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP26 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP27 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP28 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP29 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP30 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP31 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP32 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP33 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN3 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN4 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN5 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN6 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN7 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN8 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN9 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN10 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN11 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN12 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN13 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_21

.SUBCKT multi_finger_inv_22 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP8 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP9 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP10 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP11 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP12 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP13 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP14 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP15 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP16 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP17 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP18 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP19 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP20 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP21 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP22 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP23 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP24 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP25 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP26 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP27 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP28 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP29 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP30 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP31 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP32 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP33 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP34 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP35 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP36 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP37 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP38 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP39 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP40 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP41 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP42 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP43 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP44 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP45 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP46 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP47 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP48 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP49 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP50 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP51 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP52 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP53 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP54 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP55 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP56 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP57 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP58 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP59 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP60 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP61 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP62 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP63 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP64 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP65 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP66 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP67 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP68 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP69 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP70 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP71 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP72 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP73 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP74 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP75 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP76 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP77 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP78 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP79 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP80 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP81 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP82 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP83 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP84 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP85 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP86 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP87 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP88 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP89 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP90 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN3 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN4 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN5 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN6 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN7 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN8 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN9 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN10 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN11 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN12 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN13 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN14 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN15 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN16 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN17 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN18 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN19 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN20 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN21 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN22 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN23 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN24 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN25 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN26 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN27 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN28 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN29 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN30 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN31 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN32 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN33 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN34 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN35 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_22

.SUBCKT decoder_stage_6 vdd vss y[0] y[1] y[2] y[3] y_b[0] y_b[1] y_b[2] y_b[3] predecode_0_0 predecode_0_1 predecode_1_0 predecode_1_1

  Xgate_0_0_0 vdd vss predecode_0_0 predecode_1_0 x_0[0] nand2_1
  Xgate_0_1_0 vdd vss predecode_0_1 predecode_1_0 x_0[1] nand2_1
  Xgate_0_2_0 vdd vss predecode_0_0 predecode_1_1 x_0[2] nand2_1
  Xgate_0_3_0 vdd vss predecode_0_1 predecode_1_1 x_0[3] nand2_1
  Xgate_1_0_0 vdd vss x_0[0] x_1[0] multi_finger_inv_18
  Xgate_1_1_0 vdd vss x_0[1] x_1[1] multi_finger_inv_18
  Xgate_1_2_0 vdd vss x_0[2] x_1[2] multi_finger_inv_18
  Xgate_1_3_0 vdd vss x_0[3] x_1[3] multi_finger_inv_18
  Xgate_2_0_0 vdd vss x_1[0] x_2[0] multi_finger_inv_19
  Xgate_2_0_1 vdd vss x_1[0] x_2[0] multi_finger_inv_19
  Xgate_2_0_2 vdd vss x_1[0] x_2[0] multi_finger_inv_19
  Xgate_2_1_0 vdd vss x_1[1] x_2[1] multi_finger_inv_19
  Xgate_2_1_1 vdd vss x_1[1] x_2[1] multi_finger_inv_19
  Xgate_2_1_2 vdd vss x_1[1] x_2[1] multi_finger_inv_19
  Xgate_2_2_0 vdd vss x_1[2] x_2[2] multi_finger_inv_19
  Xgate_2_2_1 vdd vss x_1[2] x_2[2] multi_finger_inv_19
  Xgate_2_2_2 vdd vss x_1[2] x_2[2] multi_finger_inv_19
  Xgate_2_3_0 vdd vss x_1[3] x_2[3] multi_finger_inv_19
  Xgate_2_3_1 vdd vss x_1[3] x_2[3] multi_finger_inv_19
  Xgate_2_3_2 vdd vss x_1[3] x_2[3] multi_finger_inv_19
  Xgate_3_0_0 vdd vss x_2[0] x_3[0] multi_finger_inv_20
  Xgate_3_0_1 vdd vss x_2[0] x_3[0] multi_finger_inv_20
  Xgate_3_0_2 vdd vss x_2[0] x_3[0] multi_finger_inv_20
  Xgate_3_0_3 vdd vss x_2[0] x_3[0] multi_finger_inv_20
  Xgate_3_0_4 vdd vss x_2[0] x_3[0] multi_finger_inv_20
  Xgate_3_1_0 vdd vss x_2[1] x_3[1] multi_finger_inv_20
  Xgate_3_1_1 vdd vss x_2[1] x_3[1] multi_finger_inv_20
  Xgate_3_1_2 vdd vss x_2[1] x_3[1] multi_finger_inv_20
  Xgate_3_1_3 vdd vss x_2[1] x_3[1] multi_finger_inv_20
  Xgate_3_1_4 vdd vss x_2[1] x_3[1] multi_finger_inv_20
  Xgate_3_2_0 vdd vss x_2[2] x_3[2] multi_finger_inv_20
  Xgate_3_2_1 vdd vss x_2[2] x_3[2] multi_finger_inv_20
  Xgate_3_2_2 vdd vss x_2[2] x_3[2] multi_finger_inv_20
  Xgate_3_2_3 vdd vss x_2[2] x_3[2] multi_finger_inv_20
  Xgate_3_2_4 vdd vss x_2[2] x_3[2] multi_finger_inv_20
  Xgate_3_3_0 vdd vss x_2[3] x_3[3] multi_finger_inv_20
  Xgate_3_3_1 vdd vss x_2[3] x_3[3] multi_finger_inv_20
  Xgate_3_3_2 vdd vss x_2[3] x_3[3] multi_finger_inv_20
  Xgate_3_3_3 vdd vss x_2[3] x_3[3] multi_finger_inv_20
  Xgate_3_3_4 vdd vss x_2[3] x_3[3] multi_finger_inv_20
  Xgate_4_0_0 vdd vss x_3[0] y_b[0] multi_finger_inv_21
  Xgate_4_0_1 vdd vss x_3[0] y_b[0] multi_finger_inv_21
  Xgate_4_0_2 vdd vss x_3[0] y_b[0] multi_finger_inv_21
  Xgate_4_0_3 vdd vss x_3[0] y_b[0] multi_finger_inv_21
  Xgate_4_0_4 vdd vss x_3[0] y_b[0] multi_finger_inv_21
  Xgate_4_1_0 vdd vss x_3[1] y_b[1] multi_finger_inv_21
  Xgate_4_1_1 vdd vss x_3[1] y_b[1] multi_finger_inv_21
  Xgate_4_1_2 vdd vss x_3[1] y_b[1] multi_finger_inv_21
  Xgate_4_1_3 vdd vss x_3[1] y_b[1] multi_finger_inv_21
  Xgate_4_1_4 vdd vss x_3[1] y_b[1] multi_finger_inv_21
  Xgate_4_2_0 vdd vss x_3[2] y_b[2] multi_finger_inv_21
  Xgate_4_2_1 vdd vss x_3[2] y_b[2] multi_finger_inv_21
  Xgate_4_2_2 vdd vss x_3[2] y_b[2] multi_finger_inv_21
  Xgate_4_2_3 vdd vss x_3[2] y_b[2] multi_finger_inv_21
  Xgate_4_2_4 vdd vss x_3[2] y_b[2] multi_finger_inv_21
  Xgate_4_3_0 vdd vss x_3[3] y_b[3] multi_finger_inv_21
  Xgate_4_3_1 vdd vss x_3[3] y_b[3] multi_finger_inv_21
  Xgate_4_3_2 vdd vss x_3[3] y_b[3] multi_finger_inv_21
  Xgate_4_3_3 vdd vss x_3[3] y_b[3] multi_finger_inv_21
  Xgate_4_3_4 vdd vss x_3[3] y_b[3] multi_finger_inv_21
  Xgate_5_0_0 vdd vss y_b[0] y[0] multi_finger_inv_22
  Xgate_5_0_1 vdd vss y_b[0] y[0] multi_finger_inv_22
  Xgate_5_0_2 vdd vss y_b[0] y[0] multi_finger_inv_22
  Xgate_5_0_3 vdd vss y_b[0] y[0] multi_finger_inv_22
  Xgate_5_0_4 vdd vss y_b[0] y[0] multi_finger_inv_22
  Xgate_5_1_0 vdd vss y_b[1] y[1] multi_finger_inv_22
  Xgate_5_1_1 vdd vss y_b[1] y[1] multi_finger_inv_22
  Xgate_5_1_2 vdd vss y_b[1] y[1] multi_finger_inv_22
  Xgate_5_1_3 vdd vss y_b[1] y[1] multi_finger_inv_22
  Xgate_5_1_4 vdd vss y_b[1] y[1] multi_finger_inv_22
  Xgate_5_2_0 vdd vss y_b[2] y[2] multi_finger_inv_22
  Xgate_5_2_1 vdd vss y_b[2] y[2] multi_finger_inv_22
  Xgate_5_2_2 vdd vss y_b[2] y[2] multi_finger_inv_22
  Xgate_5_2_3 vdd vss y_b[2] y[2] multi_finger_inv_22
  Xgate_5_2_4 vdd vss y_b[2] y[2] multi_finger_inv_22
  Xgate_5_3_0 vdd vss y_b[3] y[3] multi_finger_inv_22
  Xgate_5_3_1 vdd vss y_b[3] y[3] multi_finger_inv_22
  Xgate_5_3_2 vdd vss y_b[3] y[3] multi_finger_inv_22
  Xgate_5_3_3 vdd vss y_b[3] y[3] multi_finger_inv_22
  Xgate_5_3_4 vdd vss y_b[3] y[3] multi_finger_inv_22

.ENDS decoder_stage_6

.SUBCKT decoder_1 vdd vss y[0] y[1] y[2] y[3] y_b[0] y_b[1] y_b[2] y_b[3] predecode_0_0 predecode_0_1 predecode_1_0 predecode_1_1

  X0 vdd vss y[0] y[1] y[2] y[3] y_b[0] y_b[1] y_b[2] y_b[3] predecode_0_0 predecode_0_1 predecode_1_0 predecode_1_1 decoder_stage_6

.ENDS decoder_1

.SUBCKT sky130_fd_sc_hs__inv_16 A VGND VNB VPB VPWR Y

  X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X1 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X2 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X5 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X7 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X9 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X10 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X11 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X12 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X13 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X14 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X15 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X16 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X17 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X18 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X19 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X20 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X21 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X22 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X23 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X24 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X25 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X26 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X27 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X28 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X29 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X30 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X31 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120


.ENDS sky130_fd_sc_hs__inv_16

.SUBCKT sky130_fd_sc_hs__inv_16_wrapper A VGND VNB VPB VPWR Y

  X0 A VGND VNB VPB VPWR Y sky130_fd_sc_hs__inv_16

.ENDS sky130_fd_sc_hs__inv_16_wrapper

.SUBCKT sky130_fd_sc_hs__inv_2_wrapper A VGND VNB VPB VPWR Y

  X0 A VGND VNB VPB VPWR Y sky130_fd_sc_hs__inv_2

.ENDS sky130_fd_sc_hs__inv_2_wrapper

.SUBCKT sky130_fd_sc_hs__inv_4 A VGND VNB VPB VPWR Y

  X0 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X2 VPWR A Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X3 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X4 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X7 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740


.ENDS sky130_fd_sc_hs__inv_4

.SUBCKT sky130_fd_sc_hs__inv_4_wrapper A VGND VNB VPB VPWR Y

  X0 A VGND VNB VPB VPWR Y sky130_fd_sc_hs__inv_4

.ENDS sky130_fd_sc_hs__inv_4_wrapper

.SUBCKT inv_chain_12 din dout vdd vss

  Xinv0 din vss vss vdd vdd x[0] sky130_fd_sc_hs__inv_2_wrapper
  Xinv1 x[0] vss vss vdd vdd x[1] sky130_fd_sc_hs__inv_2_wrapper
  Xinv2 x[1] vss vss vdd vdd x[2] sky130_fd_sc_hs__inv_2_wrapper
  Xinv3 x[2] vss vss vdd vdd x[3] sky130_fd_sc_hs__inv_2_wrapper
  Xinv4 x[3] vss vss vdd vdd x[4] sky130_fd_sc_hs__inv_2_wrapper
  Xinv5 x[4] vss vss vdd vdd x[5] sky130_fd_sc_hs__inv_2_wrapper
  Xinv6 x[5] vss vss vdd vdd x[6] sky130_fd_sc_hs__inv_2_wrapper
  Xinv7 x[6] vss vss vdd vdd x[7] sky130_fd_sc_hs__inv_2_wrapper
  Xinv8 x[7] vss vss vdd vdd x[8] sky130_fd_sc_hs__inv_2_wrapper
  Xinv9 x[8] vss vss vdd vdd x[9] sky130_fd_sc_hs__inv_2_wrapper
  Xinv10 x[9] vss vss vdd vdd x[10] sky130_fd_sc_hs__inv_2_wrapper
  Xinv11 x[10] vss vss vdd vdd dout sky130_fd_sc_hs__inv_4_wrapper

.ENDS inv_chain_12

.SUBCKT sky130_fd_sc_hs__and2_2 A B VGND VNB VPB VPWR X

  X0 a_31_74# B VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X1 X a_31_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X2 X a_31_74# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X3 a_118_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X4 a_31_74# A a_118_74# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X5 VPWR A a_31_74# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X6 VPWR a_31_74# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X7 VGND a_31_74# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740


.ENDS sky130_fd_sc_hs__and2_2

.SUBCKT sky130_fd_sc_hs__and2_2_wrapper A B VGND VNB VPB VPWR X

  X0 A B VGND VNB VPB VPWR X sky130_fd_sc_hs__and2_2

.ENDS sky130_fd_sc_hs__and2_2_wrapper

.SUBCKT inv_chain_9 din dout vdd vss

  Xinv0 din vss vss vdd vdd x[0] sky130_fd_sc_hs__inv_2_wrapper
  Xinv1 x[0] vss vss vdd vdd x[1] sky130_fd_sc_hs__inv_2_wrapper
  Xinv2 x[1] vss vss vdd vdd x[2] sky130_fd_sc_hs__inv_2_wrapper
  Xinv3 x[2] vss vss vdd vdd x[3] sky130_fd_sc_hs__inv_2_wrapper
  Xinv4 x[3] vss vss vdd vdd x[4] sky130_fd_sc_hs__inv_2_wrapper
  Xinv5 x[4] vss vss vdd vdd x[5] sky130_fd_sc_hs__inv_2_wrapper
  Xinv6 x[5] vss vss vdd vdd x[6] sky130_fd_sc_hs__inv_2_wrapper
  Xinv7 x[6] vss vss vdd vdd x[7] sky130_fd_sc_hs__inv_2_wrapper
  Xinv8 x[7] vss vss vdd vdd dout sky130_fd_sc_hs__inv_4_wrapper

.ENDS inv_chain_9

.SUBCKT edge_detector din dout vdd vss

  Xdelay_chain din delayed vdd vss inv_chain_9
  Xand din delayed vss vss vdd vdd dout sky130_fd_sc_hs__and2_4_wrapper

.ENDS edge_detector

.SUBCKT sky130_fd_sc_hs__buf_16 A VGND VNB VPB VPWR X

  X0 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X1 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X2 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X3 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X4 VPWR A a_83_260# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X5 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X6 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X7 VPWR A a_83_260# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X8 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X9 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X10 VPWR A a_83_260# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X11 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X12 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X13 a_83_260# A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X14 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X15 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X16 VGND A a_83_260# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X17 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X18 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X19 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X20 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X21 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X22 VGND A a_83_260# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X23 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X24 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X25 a_83_260# A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X26 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X27 a_83_260# A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X28 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X29 a_83_260# A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X30 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X31 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X32 a_83_260# A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X33 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X34 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X35 a_83_260# A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X36 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X37 VGND A a_83_260# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X38 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X39 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X40 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X41 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X42 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X43 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740


.ENDS sky130_fd_sc_hs__buf_16

.SUBCKT sky130_fd_sc_hs__buf_16_wrapper A VGND VNB VPB VPWR X

  X0 A VGND VNB VPB VPWR X sky130_fd_sc_hs__buf_16

.ENDS sky130_fd_sc_hs__buf_16_wrapper

.SUBCKT inv_chain_3 din dout vdd vss

  Xinv0 din vss vss vdd vdd x[0] sky130_fd_sc_hs__inv_2_wrapper
  Xinv1 x[0] vss vss vdd vdd x[1] sky130_fd_sc_hs__inv_2_wrapper
  Xinv2 x[1] vss vss vdd vdd dout sky130_fd_sc_hs__inv_4_wrapper

.ENDS inv_chain_3

.SUBCKT inv_chain_27 din dout vdd vss

  Xinv0 din vss vss vdd vdd x[0] sky130_fd_sc_hs__inv_2_wrapper
  Xinv1 x[0] vss vss vdd vdd x[1] sky130_fd_sc_hs__inv_2_wrapper
  Xinv2 x[1] vss vss vdd vdd x[2] sky130_fd_sc_hs__inv_2_wrapper
  Xinv3 x[2] vss vss vdd vdd x[3] sky130_fd_sc_hs__inv_2_wrapper
  Xinv4 x[3] vss vss vdd vdd x[4] sky130_fd_sc_hs__inv_2_wrapper
  Xinv5 x[4] vss vss vdd vdd x[5] sky130_fd_sc_hs__inv_2_wrapper
  Xinv6 x[5] vss vss vdd vdd x[6] sky130_fd_sc_hs__inv_2_wrapper
  Xinv7 x[6] vss vss vdd vdd x[7] sky130_fd_sc_hs__inv_2_wrapper
  Xinv8 x[7] vss vss vdd vdd x[8] sky130_fd_sc_hs__inv_2_wrapper
  Xinv9 x[8] vss vss vdd vdd x[9] sky130_fd_sc_hs__inv_2_wrapper
  Xinv10 x[9] vss vss vdd vdd x[10] sky130_fd_sc_hs__inv_2_wrapper
  Xinv11 x[10] vss vss vdd vdd x[11] sky130_fd_sc_hs__inv_2_wrapper
  Xinv12 x[11] vss vss vdd vdd x[12] sky130_fd_sc_hs__inv_2_wrapper
  Xinv13 x[12] vss vss vdd vdd x[13] sky130_fd_sc_hs__inv_2_wrapper
  Xinv14 x[13] vss vss vdd vdd x[14] sky130_fd_sc_hs__inv_2_wrapper
  Xinv15 x[14] vss vss vdd vdd x[15] sky130_fd_sc_hs__inv_2_wrapper
  Xinv16 x[15] vss vss vdd vdd x[16] sky130_fd_sc_hs__inv_2_wrapper
  Xinv17 x[16] vss vss vdd vdd x[17] sky130_fd_sc_hs__inv_2_wrapper
  Xinv18 x[17] vss vss vdd vdd x[18] sky130_fd_sc_hs__inv_2_wrapper
  Xinv19 x[18] vss vss vdd vdd x[19] sky130_fd_sc_hs__inv_2_wrapper
  Xinv20 x[19] vss vss vdd vdd x[20] sky130_fd_sc_hs__inv_2_wrapper
  Xinv21 x[20] vss vss vdd vdd x[21] sky130_fd_sc_hs__inv_2_wrapper
  Xinv22 x[21] vss vss vdd vdd x[22] sky130_fd_sc_hs__inv_2_wrapper
  Xinv23 x[22] vss vss vdd vdd x[23] sky130_fd_sc_hs__inv_2_wrapper
  Xinv24 x[23] vss vss vdd vdd x[24] sky130_fd_sc_hs__inv_2_wrapper
  Xinv25 x[24] vss vss vdd vdd x[25] sky130_fd_sc_hs__inv_2_wrapper
  Xinv26 x[25] vss vss vdd vdd dout sky130_fd_sc_hs__inv_4_wrapper

.ENDS inv_chain_27

.SUBCKT sky130_fd_sc_hs__mux2_4 A0 A1 S VGND VNB VPB VPWR X

  X0 a_27_368# S VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X1 a_722_391# A0 a_193_241# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X2 a_722_391# S VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X3 VGND a_27_368# a_937_119# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X4 a_193_241# A1 a_936_391# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X5 a_709_119# S VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X6 a_709_119# A1 a_193_241# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X7 X a_193_241# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X8 X a_193_241# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X9 VPWR a_27_368# a_936_391# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X10 X a_193_241# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X11 a_193_241# A0 a_722_391# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X12 a_937_119# A0 a_193_241# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X13 a_936_391# a_27_368# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X14 VGND a_193_241# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X15 VPWR a_193_241# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X16 VPWR S a_722_391# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X17 a_936_391# A1 a_193_241# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.000

  X18 a_193_241# A0 a_937_119# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X19 a_193_241# A1 a_709_119# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X20 X a_193_241# VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X21 VGND a_193_241# X VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X22 a_27_368# S VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X23 a_937_119# a_27_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640

  X24 VPWR a_193_241# X VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X25 VGND S a_709_119# VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.640


.ENDS sky130_fd_sc_hs__mux2_4

.SUBCKT sky130_fd_sc_hs__mux2_4_wrapper A0 A1 S VGND VNB VPB VPWR X

  X0 A0 A1 S VGND VNB VPB VPWR X sky130_fd_sc_hs__mux2_4

.ENDS sky130_fd_sc_hs__mux2_4_wrapper

.SUBCKT inv_chain_18 din dout vdd vss

  Xinv0 din vss vss vdd vdd x[0] sky130_fd_sc_hs__inv_2_wrapper
  Xinv1 x[0] vss vss vdd vdd x[1] sky130_fd_sc_hs__inv_2_wrapper
  Xinv2 x[1] vss vss vdd vdd x[2] sky130_fd_sc_hs__inv_2_wrapper
  Xinv3 x[2] vss vss vdd vdd x[3] sky130_fd_sc_hs__inv_2_wrapper
  Xinv4 x[3] vss vss vdd vdd x[4] sky130_fd_sc_hs__inv_2_wrapper
  Xinv5 x[4] vss vss vdd vdd x[5] sky130_fd_sc_hs__inv_2_wrapper
  Xinv6 x[5] vss vss vdd vdd x[6] sky130_fd_sc_hs__inv_2_wrapper
  Xinv7 x[6] vss vss vdd vdd x[7] sky130_fd_sc_hs__inv_2_wrapper
  Xinv8 x[7] vss vss vdd vdd x[8] sky130_fd_sc_hs__inv_2_wrapper
  Xinv9 x[8] vss vss vdd vdd x[9] sky130_fd_sc_hs__inv_2_wrapper
  Xinv10 x[9] vss vss vdd vdd x[10] sky130_fd_sc_hs__inv_2_wrapper
  Xinv11 x[10] vss vss vdd vdd x[11] sky130_fd_sc_hs__inv_2_wrapper
  Xinv12 x[11] vss vss vdd vdd x[12] sky130_fd_sc_hs__inv_2_wrapper
  Xinv13 x[12] vss vss vdd vdd x[13] sky130_fd_sc_hs__inv_2_wrapper
  Xinv14 x[13] vss vss vdd vdd x[14] sky130_fd_sc_hs__inv_2_wrapper
  Xinv15 x[14] vss vss vdd vdd x[15] sky130_fd_sc_hs__inv_2_wrapper
  Xinv16 x[15] vss vss vdd vdd x[16] sky130_fd_sc_hs__inv_2_wrapper
  Xinv17 x[16] vss vss vdd vdd dout sky130_fd_sc_hs__inv_4_wrapper

.ENDS inv_chain_18

.SUBCKT sky130_fd_sc_hs__nor2_4 A B VGND VNB VPB VPWR Y

  X0 a_27_368# A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X1 a_27_368# B Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X2 VGND B Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X3 a_27_368# A VPWR VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X4 Y B a_27_368# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X5 a_27_368# B Y VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X6 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X7 VPWR A a_27_368# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X8 VPWR A a_27_368# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120

  X9 Y A VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X10 Y B VGND VNB sky130_fd_pr__nfet_01v8_lvt l=0.150 nf=1 w=0.740

  X11 Y B a_27_368# VPB sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.120


.ENDS sky130_fd_sc_hs__nor2_4

.SUBCKT sky130_fd_sc_hs__nor2_4_wrapper A B VGND VNB VPB VPWR Y

  X0 A B VGND VNB VPB VPWR Y sky130_fd_sc_hs__nor2_4

.ENDS sky130_fd_sc_hs__nor2_4_wrapper

.SUBCKT sr_latch sb rb q qb vdd vss

  Xnand_set q0b sb vss vss vdd vdd q0 sky130_fd_sc_hs__nand2_8_wrapper
  Xnand_reset q0 rb vss vss vdd vdd q0b sky130_fd_sc_hs__nand2_8_wrapper
  Xqb_inv q0 vss vss vdd vdd qb sky130_fd_sc_hs__inv_2_wrapper
  Xq_inv q0b vss vss vdd vdd q sky130_fd_sc_hs__inv_2_wrapper

.ENDS sr_latch

.SUBCKT inv_chain_2 din dout vdd vss

  Xinv0 din vss vss vdd vdd x sky130_fd_sc_hs__inv_2_wrapper
  Xinv1 x vss vss vdd vdd dout sky130_fd_sc_hs__inv_4_wrapper

.ENDS inv_chain_2

.SUBCKT control_logic_replica_v2 clk ce we rstb rbl saen pc_b rwl wlen wrdrven vdd vss

  Xreset_inv rstb vss vss vdd vdd reset sky130_fd_sc_hs__inv_16_wrapper
  Xclk_delay clk clkd vdd vss inv_chain_12
  Xclk_gate clkd ce vss vss vdd vdd clk_buf sky130_fd_sc_hs__and2_2_wrapper
  Xclk_pulse clk_buf clkp0 vdd vss edge_detector
  Xclk_pulse_buf clkp0 vss vss vdd vdd clkp sky130_fd_sc_hs__buf_16_wrapper
  Xclk_pulse_inv clkp vss vss vdd vdd clkp_b sky130_fd_sc_hs__inv_16_wrapper
  Xclkp_delay clkp_b clkpd vdd vss inv_chain_3
  Xclkpd_inv clkpd vss vss vdd vdd clkpd_b sky130_fd_sc_hs__inv_2_wrapper
  Xclkpd_delay clkpd_b clkpdd vdd vss inv_chain_27
  Xmux_wlen_rst rbl_b clkpdd we vss vss vdd vdd decrepstart sky130_fd_sc_hs__mux2_4_wrapper
  Xdecoder_replica decrepstart decrepend vdd vss svt_inv_chain_22
  Xdecoder_replica_delay decrepend wlen_rst_decoderd vdd vss inv_chain_18
  Xinv_we we vss vss vdd vdd we_b sky130_fd_sc_hs__inv_2_wrapper
  Xinv_rbl rbl vss vss vdd vdd rbl_b sky130_fd_sc_hs__inv_2_wrapper
  Xwlen_grst decrepstart reset vss vss vdd vdd wlen_grst_b sky130_fd_sc_hs__nor2_4_wrapper
  Xpc_set wlen_rst_decoderd reset vss vss vdd vdd pc_set_b sky130_fd_sc_hs__nor2_4_wrapper
  Xwrdrven_grst decrepend reset vss vss vdd vdd wrdrven_grst_b sky130_fd_sc_hs__nor2_4_wrapper
  Xclkp_grst clkp reset vss vss vdd vdd clkp_grst_b sky130_fd_sc_hs__nor2_4_wrapper
  Xnand_sense_en we_b decrepend vss vss vdd vdd saen_set_b sky130_fd_sc_hs__nand2_4_wrapper
  Xnand_wlendb_web rbl_b we_b vss vss vdd vdd wlend sky130_fd_sc_hs__nand2_4_wrapper
  Xand_wlen wlen_q wlend vss vss vdd vdd wlen sky130_fd_sc_hs__and2_4_wrapper
  Xrwl_buf wlen_q vss vss vdd vdd rwl sky130_fd_sc_hs__buf_16_wrapper
  Xwl_ctl clkpd_b wlen_grst_b wlen_q wlen_b vdd vss sr_latch
  Xsaen_ctl saen_set_b clkp_grst_b saen saen_b vdd vss sr_latch
  Xpc_ctl pc_set_b clkp_b pc pc_b0 vdd vss sr_latch
  Xpc_b_buf pc_b0 vss vss vdd vdd pc_b sky130_fd_sc_hs__buf_16_wrapper
  Xwrdrven_set clkpd we vss vss vdd vdd wrdrven_set_b0 sky130_fd_sc_hs__nand2_4_wrapper
  Xwrdrven_set_delay wrdrven_set_b0 wrdrven_set_b vdd vss inv_chain_2
  Xwrdrven_ctl wrdrven_set_b wrdrven_grst_b wrdrven wrdrven_b vdd vss sr_latch

.ENDS control_logic_replica_v2

.SUBCKT mos_w1250_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.250


.ENDS mos_w1250_l150_m1_nf1_id1

.SUBCKT mos_w500_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.500


.ENDS mos_w500_l150_m1_nf1_id0

.SUBCKT folded_inv vdd vss a y

  XMP0 y a vdd vdd mos_w1250_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w500_l150_m1_nf1_id0
  XMP1 y a vdd vdd mos_w1250_l150_m1_nf1_id1
  XMN1 y a vss vss mos_w500_l150_m1_nf1_id0

.ENDS folded_inv

.SUBCKT multi_finger_inv vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP8 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP9 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP10 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN3 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv

.SUBCKT multi_finger_inv_1 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_1

.SUBCKT multi_finger_inv_2 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_2

.SUBCKT multi_finger_inv_3 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP8 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP9 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP10 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP11 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP12 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP13 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP14 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP15 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP16 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP17 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN3 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN4 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN5 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN6 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_3

.SUBCKT decoder_stage_1 vdd vss y y_b predecode_0_0

  Xgate_0_0_0 vdd vss predecode_0_0 x_0 folded_inv
  Xgate_1_0_0 vdd vss x_0 x_1 multi_finger_inv
  Xgate_2_0_0 vdd vss x_1 x_2 multi_finger_inv_1
  Xgate_2_0_1 vdd vss x_1 x_2 multi_finger_inv_1
  Xgate_2_0_2 vdd vss x_1 x_2 multi_finger_inv_1
  Xgate_2_0_3 vdd vss x_1 x_2 multi_finger_inv_1
  Xgate_3_0_0 vdd vss x_2 x_3 multi_finger_inv_2
  Xgate_3_0_1 vdd vss x_2 x_3 multi_finger_inv_2
  Xgate_3_0_2 vdd vss x_2 x_3 multi_finger_inv_2
  Xgate_3_0_3 vdd vss x_2 x_3 multi_finger_inv_2
  Xgate_3_0_4 vdd vss x_2 x_3 multi_finger_inv_2
  Xgate_3_0_5 vdd vss x_2 x_3 multi_finger_inv_2
  Xgate_3_0_6 vdd vss x_2 x_3 multi_finger_inv_2
  Xgate_3_0_7 vdd vss x_2 x_3 multi_finger_inv_2
  Xgate_3_0_8 vdd vss x_2 x_3 multi_finger_inv_2
  Xgate_3_0_9 vdd vss x_2 x_3 multi_finger_inv_2
  Xgate_3_0_10 vdd vss x_2 x_3 multi_finger_inv_2
  Xgate_3_0_11 vdd vss x_2 x_3 multi_finger_inv_2
  Xgate_3_0_12 vdd vss x_2 x_3 multi_finger_inv_2
  Xgate_3_0_13 vdd vss x_2 x_3 multi_finger_inv_2
  Xgate_4_0_0 vdd vss x_3 y_b multi_finger_inv_3
  Xgate_4_0_1 vdd vss x_3 y_b multi_finger_inv_3
  Xgate_4_0_2 vdd vss x_3 y_b multi_finger_inv_3
  Xgate_4_0_3 vdd vss x_3 y_b multi_finger_inv_3
  Xgate_4_0_4 vdd vss x_3 y_b multi_finger_inv_3
  Xgate_4_0_5 vdd vss x_3 y_b multi_finger_inv_3
  Xgate_4_0_6 vdd vss x_3 y_b multi_finger_inv_3
  Xgate_4_0_7 vdd vss x_3 y_b multi_finger_inv_3
  Xgate_4_0_8 vdd vss x_3 y_b multi_finger_inv_3
  Xgate_4_0_9 vdd vss x_3 y_b multi_finger_inv_3
  Xgate_4_0_10 vdd vss x_3 y_b multi_finger_inv_3
  Xgate_4_0_11 vdd vss x_3 y_b multi_finger_inv_3
  Xgate_4_0_12 vdd vss x_3 y_b multi_finger_inv_3
  Xgate_4_0_13 vdd vss x_3 y_b multi_finger_inv_3
  Xgate_4_0_14 vdd vss x_3 y_b multi_finger_inv_3
  Xgate_5_0_0 vdd vss y_b y multi_finger_inv_4
  Xgate_5_0_1 vdd vss y_b y multi_finger_inv_4
  Xgate_5_0_2 vdd vss y_b y multi_finger_inv_4
  Xgate_5_0_3 vdd vss y_b y multi_finger_inv_4
  Xgate_5_0_4 vdd vss y_b y multi_finger_inv_4
  Xgate_5_0_5 vdd vss y_b y multi_finger_inv_4
  Xgate_5_0_6 vdd vss y_b y multi_finger_inv_4
  Xgate_5_0_7 vdd vss y_b y multi_finger_inv_4
  Xgate_5_0_8 vdd vss y_b y multi_finger_inv_4
  Xgate_5_0_9 vdd vss y_b y multi_finger_inv_4
  Xgate_5_0_10 vdd vss y_b y multi_finger_inv_4
  Xgate_5_0_11 vdd vss y_b y multi_finger_inv_4
  Xgate_5_0_12 vdd vss y_b y multi_finger_inv_4
  Xgate_5_0_13 vdd vss y_b y multi_finger_inv_4
  Xgate_5_0_14 vdd vss y_b y multi_finger_inv_4

.ENDS decoder_stage_1

.SUBCKT multi_finger_inv_5 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_5

.SUBCKT decoder_stage_2 vdd vss y y_b predecode_0_0

  Xgate_0_0_0 vdd vss predecode_0_0 y_b folded_inv
  Xgate_1_0_0 vdd vss y_b y multi_finger_inv_5
  Xgate_1_0_1 vdd vss y_b y multi_finger_inv_5

.ENDS decoder_stage_2

.SUBCKT multi_finger_inv_6 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP8 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_6

.SUBCKT multi_finger_inv_7 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP8 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP9 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN3 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_7

.SUBCKT multi_finger_inv_8 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP8 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP9 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP10 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP11 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP12 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP13 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP14 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP15 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP16 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP17 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP18 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP19 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP20 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP21 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP22 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP23 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN3 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN4 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN5 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN6 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN7 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN8 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN9 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_8

.SUBCKT decoder_stage_3 vdd vss y y_b predecode_0_0

  Xgate_0_0_0 vdd vss predecode_0_0 x_0 folded_inv
  Xgate_1_0_0 vdd vss x_0 x_1 multi_finger_inv_6
  Xgate_2_0_0 vdd vss x_1 y_b multi_finger_inv_7
  Xgate_2_0_1 vdd vss x_1 y_b multi_finger_inv_7
  Xgate_3_0_0 vdd vss y_b y multi_finger_inv_8
  Xgate_3_0_1 vdd vss y_b y multi_finger_inv_8

.ENDS decoder_stage_3

.SUBCKT multi_finger_inv_9 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP8 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP9 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN3 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_9

.SUBCKT multi_finger_inv_10 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_10

.SUBCKT multi_finger_inv_11 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_11

.SUBCKT multi_finger_inv_12 vdd vss a y

  XMP0 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP1 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP2 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP3 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP4 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP5 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP6 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP7 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP8 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP9 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP10 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP11 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP12 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP13 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP14 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP15 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP16 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP17 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP18 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMP19 y a vdd vdd mos_w700_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN1 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN2 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN3 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN4 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN5 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN6 y a vss vss mos_w700_l150_m1_nf1_id0
  XMN7 y a vss vss mos_w700_l150_m1_nf1_id0

.ENDS multi_finger_inv_12

.SUBCKT decoder_stage_4 vdd vss y y_b predecode_0_0

  Xgate_0_0_0 vdd vss predecode_0_0 x_0 folded_inv
  Xgate_1_0_0 vdd vss x_0 x_1 multi_finger_inv_9
  Xgate_2_0_0 vdd vss x_1 x_2 multi_finger_inv_10
  Xgate_2_0_1 vdd vss x_1 x_2 multi_finger_inv_10
  Xgate_2_0_2 vdd vss x_1 x_2 multi_finger_inv_10
  Xgate_3_0_0 vdd vss x_2 x_3 multi_finger_inv_11
  Xgate_3_0_1 vdd vss x_2 x_3 multi_finger_inv_11
  Xgate_3_0_2 vdd vss x_2 x_3 multi_finger_inv_11
  Xgate_3_0_3 vdd vss x_2 x_3 multi_finger_inv_11
  Xgate_3_0_4 vdd vss x_2 x_3 multi_finger_inv_11
  Xgate_3_0_5 vdd vss x_2 x_3 multi_finger_inv_11
  Xgate_3_0_6 vdd vss x_2 x_3 multi_finger_inv_11
  Xgate_3_0_7 vdd vss x_2 x_3 multi_finger_inv_11
  Xgate_3_0_8 vdd vss x_2 x_3 multi_finger_inv_11
  Xgate_4_0_0 vdd vss x_3 y_b multi_finger_inv_12
  Xgate_4_0_1 vdd vss x_3 y_b multi_finger_inv_12
  Xgate_4_0_2 vdd vss x_3 y_b multi_finger_inv_12
  Xgate_4_0_3 vdd vss x_3 y_b multi_finger_inv_12
  Xgate_4_0_4 vdd vss x_3 y_b multi_finger_inv_12
  Xgate_4_0_5 vdd vss x_3 y_b multi_finger_inv_12
  Xgate_4_0_6 vdd vss x_3 y_b multi_finger_inv_12
  Xgate_4_0_7 vdd vss x_3 y_b multi_finger_inv_12
  Xgate_4_0_8 vdd vss x_3 y_b multi_finger_inv_12
  Xgate_5_0_0 vdd vss y_b y multi_finger_inv_13
  Xgate_5_0_1 vdd vss y_b y multi_finger_inv_13
  Xgate_5_0_2 vdd vss y_b y multi_finger_inv_13
  Xgate_5_0_3 vdd vss y_b y multi_finger_inv_13
  Xgate_5_0_4 vdd vss y_b y multi_finger_inv_13
  Xgate_5_0_5 vdd vss y_b y multi_finger_inv_13
  Xgate_5_0_6 vdd vss y_b y multi_finger_inv_13
  Xgate_5_0_7 vdd vss y_b y multi_finger_inv_13
  Xgate_5_0_8 vdd vss y_b y multi_finger_inv_13

.ENDS decoder_stage_4

.SUBCKT dff_array_10 vdd vss clk rb d[0] d[1] d[2] d[3] d[4] d[5] d[6] d[7] d[8] d[9] q[0] q[1] q[2] q[3] q[4] q[5] q[6] q[7] q[8] q[9] qn[0] qn[1] qn[2] qn[3] qn[4] qn[5] qn[6] qn[7] qn[8] qn[9]

  Xdff_0 clk d[0] rb vss vss vdd vdd q[0] qn[0] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_1 clk d[1] rb vss vss vdd vdd q[1] qn[1] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_2 clk d[2] rb vss vss vdd vdd q[2] qn[2] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_3 clk d[3] rb vss vss vdd vdd q[3] qn[3] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_4 clk d[4] rb vss vss vdd vdd q[4] qn[4] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_5 clk d[5] rb vss vss vdd vdd q[5] qn[5] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_6 clk d[6] rb vss vss vdd vdd q[6] qn[6] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_7 clk d[7] rb vss vss vdd vdd q[7] qn[7] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_8 clk d[8] rb vss vss vdd vdd q[8] qn[8] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_9 clk d[9] rb vss vss vdd vdd q[9] qn[9] sky130_fd_sc_hs__dfrbp_2_wrapper

.ENDS dff_array_10

.SUBCKT sram_sp_cell BL BR VDD VSS WL VNB VPB

  X0 QB WL BR VNB sky130_fd_pr__special_nfet_pass l=0.150 nf=1 w=0.140

  X1 Q QB VSS VNB sky130_fd_pr__special_nfet_latch l=0.150 nf=1 w=0.210

  X2 BL WL Q VNB sky130_fd_pr__special_nfet_pass l=0.150 nf=1 w=0.140

  X3 Q WL Q VPB sky130_fd_pr__special_pfet_pass l=0.025 nf=1 w=0.140

  X4 QB WL QB VPB sky130_fd_pr__special_pfet_pass l=0.025 nf=1 w=0.140

  X5 VDD Q QB VPB sky130_fd_pr__special_pfet_pass l=0.150 nf=1 w=0.140

  X6 Q QB VDD VPB sky130_fd_pr__special_pfet_pass l=0.150 nf=1 w=0.140

  X7 VSS Q QB VNB sky130_fd_pr__special_nfet_latch l=0.150 nf=1 w=0.210


.ENDS sram_sp_cell

.SUBCKT sram_sp_cell_wrapper BL BR VDD VSS WL VNB VPB

  X0 BL BR VDD VSS WL VNB VPB sram_sp_cell

.ENDS sram_sp_cell_wrapper

.SUBCKT sram_sp_colend BR VDD VSS BL VNB VPB

  X0 BR VNB BR VNB sky130_fd_pr__special_nfet_pass l=0.140 nf=1 w=0.140


.ENDS sram_sp_colend

.SUBCKT sram_sp_colend_wrapper BR VDD VSS BL VNB VPB

  X0 BR VDD VSS BL VNB VPB sram_sp_colend

.ENDS sram_sp_colend_wrapper

.SUBCKT sram_sp_hstrap BR VDD VSS BL VNB VPB

  X0 BL VNB BL VNB sky130_fd_pr__special_nfet_pass l=0.140 nf=1 w=0.140

  X1 BL VNB BL VNB sky130_fd_pr__special_nfet_pass l=0.140 nf=1 w=0.140


.ENDS sram_sp_hstrap

.SUBCKT sram_sp_hstrap_wrapper BR VDD VSS BL VNB VPB

  X0 BR VDD VSS BL VNB VPB sram_sp_hstrap

.ENDS sram_sp_hstrap_wrapper

.SUBCKT sram_sp_horiz_wlstrap_p2 VSS VNB

  X0 VSS VSS VSS VNB sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.420


.ENDS sram_sp_horiz_wlstrap_p2

.SUBCKT sram_sp_horiz_wlstrap_p2_wrapper VSS VNB

  X0 VSS VNB sram_sp_horiz_wlstrap_p2

.ENDS sram_sp_horiz_wlstrap_p2_wrapper

.SUBCKT sp_cell_array vdd vss dummy_bl dummy_br bl[0] bl[1] bl[2] bl[3] bl[4] bl[5] bl[6] bl[7] bl[8] bl[9] bl[10] bl[11] bl[12] bl[13] bl[14] bl[15] bl[16] bl[17] bl[18] bl[19] bl[20] bl[21] bl[22] bl[23] bl[24] bl[25] bl[26] bl[27] bl[28] bl[29] bl[30] bl[31] bl[32] bl[33] bl[34] bl[35] bl[36] bl[37] bl[38] bl[39] bl[40] bl[41] bl[42] bl[43] bl[44] bl[45] bl[46] bl[47] bl[48] bl[49] bl[50] bl[51] bl[52] bl[53] bl[54] bl[55] bl[56] bl[57] bl[58] bl[59] bl[60] bl[61] bl[62] bl[63] bl[64] bl[65] bl[66] bl[67] bl[68] bl[69] bl[70] bl[71] bl[72] bl[73] bl[74] bl[75] bl[76] bl[77] bl[78] bl[79] bl[80] bl[81] bl[82] bl[83] bl[84] bl[85] bl[86] bl[87] bl[88] bl[89] bl[90] bl[91] bl[92] bl[93] bl[94] bl[95] bl[96] bl[97] bl[98] bl[99] bl[100] bl[101] bl[102] bl[103] bl[104] bl[105] bl[106] bl[107] bl[108] bl[109] bl[110] bl[111] bl[112] bl[113] bl[114] bl[115] bl[116] bl[117] bl[118] bl[119] bl[120] bl[121] bl[122] bl[123] bl[124] bl[125] bl[126] bl[127] bl[128] bl[129] bl[130] bl[131] bl[132] bl[133] bl[134] bl[135] bl[136] bl[137] bl[138] bl[139] bl[140] bl[141] bl[142] bl[143] bl[144] bl[145] bl[146] bl[147] bl[148] bl[149] bl[150] bl[151] bl[152] bl[153] bl[154] bl[155] bl[156] bl[157] bl[158] bl[159] bl[160] bl[161] bl[162] bl[163] bl[164] bl[165] bl[166] bl[167] bl[168] bl[169] bl[170] bl[171] bl[172] bl[173] bl[174] bl[175] bl[176] bl[177] bl[178] bl[179] bl[180] bl[181] bl[182] bl[183] bl[184] bl[185] bl[186] bl[187] bl[188] bl[189] bl[190] bl[191] bl[192] bl[193] bl[194] bl[195] bl[196] bl[197] bl[198] bl[199] bl[200] bl[201] bl[202] bl[203] bl[204] bl[205] bl[206] bl[207] bl[208] bl[209] bl[210] bl[211] bl[212] bl[213] bl[214] bl[215] bl[216] bl[217] bl[218] bl[219] bl[220] bl[221] bl[222] bl[223] bl[224] bl[225] bl[226] bl[227] bl[228] bl[229] bl[230] bl[231] bl[232] bl[233] bl[234] bl[235] bl[236] bl[237] bl[238] bl[239] bl[240] bl[241] bl[242] bl[243] bl[244] bl[245] bl[246] bl[247] bl[248] bl[249] bl[250] bl[251] bl[252] bl[253] bl[254] bl[255] bl[256] bl[257] bl[258] bl[259] bl[260] bl[261] bl[262] bl[263] bl[264] bl[265] bl[266] bl[267] bl[268] bl[269] bl[270] bl[271] bl[272] bl[273] bl[274] bl[275] bl[276] bl[277] bl[278] bl[279] bl[280] bl[281] bl[282] bl[283] bl[284] bl[285] bl[286] bl[287] bl[288] bl[289] bl[290] bl[291] bl[292] bl[293] bl[294] bl[295] bl[296] bl[297] bl[298] bl[299] bl[300] bl[301] bl[302] bl[303] bl[304] bl[305] bl[306] bl[307] bl[308] bl[309] bl[310] bl[311] bl[312] bl[313] bl[314] bl[315] bl[316] bl[317] bl[318] bl[319] bl[320] bl[321] bl[322] bl[323] bl[324] bl[325] bl[326] bl[327] bl[328] bl[329] bl[330] bl[331] bl[332] bl[333] bl[334] bl[335] bl[336] bl[337] bl[338] bl[339] bl[340] bl[341] bl[342] bl[343] bl[344] bl[345] bl[346] bl[347] bl[348] bl[349] bl[350] bl[351] bl[352] bl[353] bl[354] bl[355] bl[356] bl[357] bl[358] bl[359] bl[360] bl[361] bl[362] bl[363] bl[364] bl[365] bl[366] bl[367] bl[368] bl[369] bl[370] bl[371] bl[372] bl[373] bl[374] bl[375] bl[376] bl[377] bl[378] bl[379] bl[380] bl[381] bl[382] bl[383] bl[384] bl[385] bl[386] bl[387] bl[388] bl[389] bl[390] bl[391] bl[392] bl[393] bl[394] bl[395] bl[396] bl[397] bl[398] bl[399] bl[400] bl[401] bl[402] bl[403] bl[404] bl[405] bl[406] bl[407] bl[408] bl[409] bl[410] bl[411] bl[412] bl[413] bl[414] bl[415] bl[416] bl[417] bl[418] bl[419] bl[420] bl[421] bl[422] bl[423] bl[424] bl[425] bl[426] bl[427] bl[428] bl[429] bl[430] bl[431] bl[432] bl[433] bl[434] bl[435] bl[436] bl[437] bl[438] bl[439] bl[440] bl[441] bl[442] bl[443] bl[444] bl[445] bl[446] bl[447] bl[448] bl[449] bl[450] bl[451] bl[452] bl[453] bl[454] bl[455] bl[456] bl[457] bl[458] bl[459] bl[460] bl[461] bl[462] bl[463] bl[464] bl[465] bl[466] bl[467] bl[468] bl[469] bl[470] bl[471] bl[472] bl[473] bl[474] bl[475] bl[476] bl[477] bl[478] bl[479] bl[480] bl[481] bl[482] bl[483] bl[484] bl[485] bl[486] bl[487] bl[488] bl[489] bl[490] bl[491] bl[492] bl[493] bl[494] bl[495] bl[496] bl[497] bl[498] bl[499] bl[500] bl[501] bl[502] bl[503] bl[504] bl[505] bl[506] bl[507] bl[508] bl[509] bl[510] bl[511] br[0] br[1] br[2] br[3] br[4] br[5] br[6] br[7] br[8] br[9] br[10] br[11] br[12] br[13] br[14] br[15] br[16] br[17] br[18] br[19] br[20] br[21] br[22] br[23] br[24] br[25] br[26] br[27] br[28] br[29] br[30] br[31] br[32] br[33] br[34] br[35] br[36] br[37] br[38] br[39] br[40] br[41] br[42] br[43] br[44] br[45] br[46] br[47] br[48] br[49] br[50] br[51] br[52] br[53] br[54] br[55] br[56] br[57] br[58] br[59] br[60] br[61] br[62] br[63] br[64] br[65] br[66] br[67] br[68] br[69] br[70] br[71] br[72] br[73] br[74] br[75] br[76] br[77] br[78] br[79] br[80] br[81] br[82] br[83] br[84] br[85] br[86] br[87] br[88] br[89] br[90] br[91] br[92] br[93] br[94] br[95] br[96] br[97] br[98] br[99] br[100] br[101] br[102] br[103] br[104] br[105] br[106] br[107] br[108] br[109] br[110] br[111] br[112] br[113] br[114] br[115] br[116] br[117] br[118] br[119] br[120] br[121] br[122] br[123] br[124] br[125] br[126] br[127] br[128] br[129] br[130] br[131] br[132] br[133] br[134] br[135] br[136] br[137] br[138] br[139] br[140] br[141] br[142] br[143] br[144] br[145] br[146] br[147] br[148] br[149] br[150] br[151] br[152] br[153] br[154] br[155] br[156] br[157] br[158] br[159] br[160] br[161] br[162] br[163] br[164] br[165] br[166] br[167] br[168] br[169] br[170] br[171] br[172] br[173] br[174] br[175] br[176] br[177] br[178] br[179] br[180] br[181] br[182] br[183] br[184] br[185] br[186] br[187] br[188] br[189] br[190] br[191] br[192] br[193] br[194] br[195] br[196] br[197] br[198] br[199] br[200] br[201] br[202] br[203] br[204] br[205] br[206] br[207] br[208] br[209] br[210] br[211] br[212] br[213] br[214] br[215] br[216] br[217] br[218] br[219] br[220] br[221] br[222] br[223] br[224] br[225] br[226] br[227] br[228] br[229] br[230] br[231] br[232] br[233] br[234] br[235] br[236] br[237] br[238] br[239] br[240] br[241] br[242] br[243] br[244] br[245] br[246] br[247] br[248] br[249] br[250] br[251] br[252] br[253] br[254] br[255] br[256] br[257] br[258] br[259] br[260] br[261] br[262] br[263] br[264] br[265] br[266] br[267] br[268] br[269] br[270] br[271] br[272] br[273] br[274] br[275] br[276] br[277] br[278] br[279] br[280] br[281] br[282] br[283] br[284] br[285] br[286] br[287] br[288] br[289] br[290] br[291] br[292] br[293] br[294] br[295] br[296] br[297] br[298] br[299] br[300] br[301] br[302] br[303] br[304] br[305] br[306] br[307] br[308] br[309] br[310] br[311] br[312] br[313] br[314] br[315] br[316] br[317] br[318] br[319] br[320] br[321] br[322] br[323] br[324] br[325] br[326] br[327] br[328] br[329] br[330] br[331] br[332] br[333] br[334] br[335] br[336] br[337] br[338] br[339] br[340] br[341] br[342] br[343] br[344] br[345] br[346] br[347] br[348] br[349] br[350] br[351] br[352] br[353] br[354] br[355] br[356] br[357] br[358] br[359] br[360] br[361] br[362] br[363] br[364] br[365] br[366] br[367] br[368] br[369] br[370] br[371] br[372] br[373] br[374] br[375] br[376] br[377] br[378] br[379] br[380] br[381] br[382] br[383] br[384] br[385] br[386] br[387] br[388] br[389] br[390] br[391] br[392] br[393] br[394] br[395] br[396] br[397] br[398] br[399] br[400] br[401] br[402] br[403] br[404] br[405] br[406] br[407] br[408] br[409] br[410] br[411] br[412] br[413] br[414] br[415] br[416] br[417] br[418] br[419] br[420] br[421] br[422] br[423] br[424] br[425] br[426] br[427] br[428] br[429] br[430] br[431] br[432] br[433] br[434] br[435] br[436] br[437] br[438] br[439] br[440] br[441] br[442] br[443] br[444] br[445] br[446] br[447] br[448] br[449] br[450] br[451] br[452] br[453] br[454] br[455] br[456] br[457] br[458] br[459] br[460] br[461] br[462] br[463] br[464] br[465] br[466] br[467] br[468] br[469] br[470] br[471] br[472] br[473] br[474] br[475] br[476] br[477] br[478] br[479] br[480] br[481] br[482] br[483] br[484] br[485] br[486] br[487] br[488] br[489] br[490] br[491] br[492] br[493] br[494] br[495] br[496] br[497] br[498] br[499] br[500] br[501] br[502] br[503] br[504] br[505] br[506] br[507] br[508] br[509] br[510] br[511] wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63]

  Xcell_0_0 bl[0] br[0] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_1 bl[1] br[1] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_2 bl[2] br[2] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_3 bl[3] br[3] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_4 bl[4] br[4] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_5 bl[5] br[5] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_6 bl[6] br[6] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_7 bl[7] br[7] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_8 bl[8] br[8] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_9 bl[9] br[9] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_10 bl[10] br[10] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_11 bl[11] br[11] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_12 bl[12] br[12] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_13 bl[13] br[13] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_14 bl[14] br[14] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_15 bl[15] br[15] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_16 bl[16] br[16] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_17 bl[17] br[17] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_18 bl[18] br[18] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_19 bl[19] br[19] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_20 bl[20] br[20] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_21 bl[21] br[21] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_22 bl[22] br[22] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_23 bl[23] br[23] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_24 bl[24] br[24] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_25 bl[25] br[25] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_26 bl[26] br[26] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_27 bl[27] br[27] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_28 bl[28] br[28] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_29 bl[29] br[29] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_30 bl[30] br[30] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_31 bl[31] br[31] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_32 bl[32] br[32] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_33 bl[33] br[33] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_34 bl[34] br[34] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_35 bl[35] br[35] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_36 bl[36] br[36] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_37 bl[37] br[37] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_38 bl[38] br[38] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_39 bl[39] br[39] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_40 bl[40] br[40] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_41 bl[41] br[41] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_42 bl[42] br[42] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_43 bl[43] br[43] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_44 bl[44] br[44] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_45 bl[45] br[45] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_46 bl[46] br[46] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_47 bl[47] br[47] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_48 bl[48] br[48] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_49 bl[49] br[49] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_50 bl[50] br[50] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_51 bl[51] br[51] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_52 bl[52] br[52] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_53 bl[53] br[53] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_54 bl[54] br[54] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_55 bl[55] br[55] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_56 bl[56] br[56] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_57 bl[57] br[57] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_58 bl[58] br[58] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_59 bl[59] br[59] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_60 bl[60] br[60] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_61 bl[61] br[61] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_62 bl[62] br[62] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_63 bl[63] br[63] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_64 bl[64] br[64] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_65 bl[65] br[65] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_66 bl[66] br[66] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_67 bl[67] br[67] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_68 bl[68] br[68] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_69 bl[69] br[69] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_70 bl[70] br[70] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_71 bl[71] br[71] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_72 bl[72] br[72] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_73 bl[73] br[73] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_74 bl[74] br[74] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_75 bl[75] br[75] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_76 bl[76] br[76] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_77 bl[77] br[77] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_78 bl[78] br[78] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_79 bl[79] br[79] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_80 bl[80] br[80] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_81 bl[81] br[81] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_82 bl[82] br[82] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_83 bl[83] br[83] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_84 bl[84] br[84] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_85 bl[85] br[85] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_86 bl[86] br[86] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_87 bl[87] br[87] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_88 bl[88] br[88] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_89 bl[89] br[89] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_90 bl[90] br[90] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_91 bl[91] br[91] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_92 bl[92] br[92] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_93 bl[93] br[93] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_94 bl[94] br[94] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_95 bl[95] br[95] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_96 bl[96] br[96] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_97 bl[97] br[97] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_98 bl[98] br[98] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_99 bl[99] br[99] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_100 bl[100] br[100] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_101 bl[101] br[101] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_102 bl[102] br[102] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_103 bl[103] br[103] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_104 bl[104] br[104] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_105 bl[105] br[105] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_106 bl[106] br[106] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_107 bl[107] br[107] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_108 bl[108] br[108] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_109 bl[109] br[109] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_110 bl[110] br[110] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_111 bl[111] br[111] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_112 bl[112] br[112] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_113 bl[113] br[113] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_114 bl[114] br[114] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_115 bl[115] br[115] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_116 bl[116] br[116] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_117 bl[117] br[117] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_118 bl[118] br[118] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_119 bl[119] br[119] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_120 bl[120] br[120] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_121 bl[121] br[121] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_122 bl[122] br[122] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_123 bl[123] br[123] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_124 bl[124] br[124] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_125 bl[125] br[125] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_126 bl[126] br[126] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_127 bl[127] br[127] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_128 bl[128] br[128] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_129 bl[129] br[129] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_130 bl[130] br[130] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_131 bl[131] br[131] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_132 bl[132] br[132] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_133 bl[133] br[133] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_134 bl[134] br[134] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_135 bl[135] br[135] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_136 bl[136] br[136] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_137 bl[137] br[137] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_138 bl[138] br[138] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_139 bl[139] br[139] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_140 bl[140] br[140] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_141 bl[141] br[141] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_142 bl[142] br[142] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_143 bl[143] br[143] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_144 bl[144] br[144] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_145 bl[145] br[145] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_146 bl[146] br[146] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_147 bl[147] br[147] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_148 bl[148] br[148] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_149 bl[149] br[149] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_150 bl[150] br[150] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_151 bl[151] br[151] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_152 bl[152] br[152] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_153 bl[153] br[153] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_154 bl[154] br[154] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_155 bl[155] br[155] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_156 bl[156] br[156] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_157 bl[157] br[157] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_158 bl[158] br[158] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_159 bl[159] br[159] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_160 bl[160] br[160] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_161 bl[161] br[161] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_162 bl[162] br[162] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_163 bl[163] br[163] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_164 bl[164] br[164] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_165 bl[165] br[165] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_166 bl[166] br[166] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_167 bl[167] br[167] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_168 bl[168] br[168] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_169 bl[169] br[169] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_170 bl[170] br[170] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_171 bl[171] br[171] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_172 bl[172] br[172] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_173 bl[173] br[173] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_174 bl[174] br[174] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_175 bl[175] br[175] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_176 bl[176] br[176] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_177 bl[177] br[177] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_178 bl[178] br[178] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_179 bl[179] br[179] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_180 bl[180] br[180] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_181 bl[181] br[181] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_182 bl[182] br[182] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_183 bl[183] br[183] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_184 bl[184] br[184] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_185 bl[185] br[185] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_186 bl[186] br[186] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_187 bl[187] br[187] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_188 bl[188] br[188] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_189 bl[189] br[189] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_190 bl[190] br[190] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_191 bl[191] br[191] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_192 bl[192] br[192] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_193 bl[193] br[193] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_194 bl[194] br[194] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_195 bl[195] br[195] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_196 bl[196] br[196] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_197 bl[197] br[197] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_198 bl[198] br[198] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_199 bl[199] br[199] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_200 bl[200] br[200] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_201 bl[201] br[201] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_202 bl[202] br[202] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_203 bl[203] br[203] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_204 bl[204] br[204] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_205 bl[205] br[205] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_206 bl[206] br[206] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_207 bl[207] br[207] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_208 bl[208] br[208] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_209 bl[209] br[209] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_210 bl[210] br[210] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_211 bl[211] br[211] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_212 bl[212] br[212] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_213 bl[213] br[213] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_214 bl[214] br[214] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_215 bl[215] br[215] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_216 bl[216] br[216] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_217 bl[217] br[217] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_218 bl[218] br[218] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_219 bl[219] br[219] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_220 bl[220] br[220] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_221 bl[221] br[221] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_222 bl[222] br[222] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_223 bl[223] br[223] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_224 bl[224] br[224] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_225 bl[225] br[225] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_226 bl[226] br[226] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_227 bl[227] br[227] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_228 bl[228] br[228] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_229 bl[229] br[229] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_230 bl[230] br[230] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_231 bl[231] br[231] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_232 bl[232] br[232] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_233 bl[233] br[233] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_234 bl[234] br[234] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_235 bl[235] br[235] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_236 bl[236] br[236] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_237 bl[237] br[237] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_238 bl[238] br[238] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_239 bl[239] br[239] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_240 bl[240] br[240] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_241 bl[241] br[241] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_242 bl[242] br[242] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_243 bl[243] br[243] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_244 bl[244] br[244] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_245 bl[245] br[245] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_246 bl[246] br[246] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_247 bl[247] br[247] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_248 bl[248] br[248] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_249 bl[249] br[249] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_250 bl[250] br[250] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_251 bl[251] br[251] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_252 bl[252] br[252] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_253 bl[253] br[253] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_254 bl[254] br[254] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_255 bl[255] br[255] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_256 bl[256] br[256] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_257 bl[257] br[257] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_258 bl[258] br[258] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_259 bl[259] br[259] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_260 bl[260] br[260] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_261 bl[261] br[261] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_262 bl[262] br[262] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_263 bl[263] br[263] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_264 bl[264] br[264] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_265 bl[265] br[265] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_266 bl[266] br[266] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_267 bl[267] br[267] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_268 bl[268] br[268] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_269 bl[269] br[269] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_270 bl[270] br[270] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_271 bl[271] br[271] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_272 bl[272] br[272] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_273 bl[273] br[273] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_274 bl[274] br[274] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_275 bl[275] br[275] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_276 bl[276] br[276] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_277 bl[277] br[277] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_278 bl[278] br[278] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_279 bl[279] br[279] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_280 bl[280] br[280] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_281 bl[281] br[281] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_282 bl[282] br[282] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_283 bl[283] br[283] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_284 bl[284] br[284] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_285 bl[285] br[285] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_286 bl[286] br[286] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_287 bl[287] br[287] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_288 bl[288] br[288] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_289 bl[289] br[289] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_290 bl[290] br[290] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_291 bl[291] br[291] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_292 bl[292] br[292] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_293 bl[293] br[293] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_294 bl[294] br[294] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_295 bl[295] br[295] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_296 bl[296] br[296] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_297 bl[297] br[297] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_298 bl[298] br[298] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_299 bl[299] br[299] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_300 bl[300] br[300] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_301 bl[301] br[301] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_302 bl[302] br[302] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_303 bl[303] br[303] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_304 bl[304] br[304] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_305 bl[305] br[305] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_306 bl[306] br[306] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_307 bl[307] br[307] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_308 bl[308] br[308] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_309 bl[309] br[309] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_310 bl[310] br[310] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_311 bl[311] br[311] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_312 bl[312] br[312] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_313 bl[313] br[313] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_314 bl[314] br[314] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_315 bl[315] br[315] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_316 bl[316] br[316] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_317 bl[317] br[317] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_318 bl[318] br[318] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_319 bl[319] br[319] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_320 bl[320] br[320] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_321 bl[321] br[321] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_322 bl[322] br[322] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_323 bl[323] br[323] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_324 bl[324] br[324] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_325 bl[325] br[325] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_326 bl[326] br[326] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_327 bl[327] br[327] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_328 bl[328] br[328] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_329 bl[329] br[329] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_330 bl[330] br[330] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_331 bl[331] br[331] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_332 bl[332] br[332] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_333 bl[333] br[333] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_334 bl[334] br[334] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_335 bl[335] br[335] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_336 bl[336] br[336] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_337 bl[337] br[337] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_338 bl[338] br[338] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_339 bl[339] br[339] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_340 bl[340] br[340] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_341 bl[341] br[341] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_342 bl[342] br[342] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_343 bl[343] br[343] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_344 bl[344] br[344] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_345 bl[345] br[345] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_346 bl[346] br[346] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_347 bl[347] br[347] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_348 bl[348] br[348] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_349 bl[349] br[349] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_350 bl[350] br[350] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_351 bl[351] br[351] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_352 bl[352] br[352] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_353 bl[353] br[353] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_354 bl[354] br[354] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_355 bl[355] br[355] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_356 bl[356] br[356] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_357 bl[357] br[357] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_358 bl[358] br[358] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_359 bl[359] br[359] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_360 bl[360] br[360] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_361 bl[361] br[361] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_362 bl[362] br[362] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_363 bl[363] br[363] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_364 bl[364] br[364] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_365 bl[365] br[365] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_366 bl[366] br[366] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_367 bl[367] br[367] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_368 bl[368] br[368] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_369 bl[369] br[369] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_370 bl[370] br[370] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_371 bl[371] br[371] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_372 bl[372] br[372] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_373 bl[373] br[373] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_374 bl[374] br[374] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_375 bl[375] br[375] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_376 bl[376] br[376] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_377 bl[377] br[377] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_378 bl[378] br[378] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_379 bl[379] br[379] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_380 bl[380] br[380] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_381 bl[381] br[381] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_382 bl[382] br[382] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_383 bl[383] br[383] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_384 bl[384] br[384] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_385 bl[385] br[385] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_386 bl[386] br[386] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_387 bl[387] br[387] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_388 bl[388] br[388] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_389 bl[389] br[389] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_390 bl[390] br[390] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_391 bl[391] br[391] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_392 bl[392] br[392] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_393 bl[393] br[393] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_394 bl[394] br[394] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_395 bl[395] br[395] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_396 bl[396] br[396] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_397 bl[397] br[397] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_398 bl[398] br[398] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_399 bl[399] br[399] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_400 bl[400] br[400] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_401 bl[401] br[401] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_402 bl[402] br[402] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_403 bl[403] br[403] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_404 bl[404] br[404] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_405 bl[405] br[405] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_406 bl[406] br[406] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_407 bl[407] br[407] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_408 bl[408] br[408] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_409 bl[409] br[409] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_410 bl[410] br[410] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_411 bl[411] br[411] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_412 bl[412] br[412] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_413 bl[413] br[413] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_414 bl[414] br[414] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_415 bl[415] br[415] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_416 bl[416] br[416] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_417 bl[417] br[417] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_418 bl[418] br[418] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_419 bl[419] br[419] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_420 bl[420] br[420] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_421 bl[421] br[421] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_422 bl[422] br[422] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_423 bl[423] br[423] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_424 bl[424] br[424] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_425 bl[425] br[425] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_426 bl[426] br[426] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_427 bl[427] br[427] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_428 bl[428] br[428] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_429 bl[429] br[429] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_430 bl[430] br[430] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_431 bl[431] br[431] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_432 bl[432] br[432] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_433 bl[433] br[433] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_434 bl[434] br[434] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_435 bl[435] br[435] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_436 bl[436] br[436] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_437 bl[437] br[437] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_438 bl[438] br[438] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_439 bl[439] br[439] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_440 bl[440] br[440] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_441 bl[441] br[441] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_442 bl[442] br[442] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_443 bl[443] br[443] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_444 bl[444] br[444] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_445 bl[445] br[445] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_446 bl[446] br[446] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_447 bl[447] br[447] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_448 bl[448] br[448] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_449 bl[449] br[449] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_450 bl[450] br[450] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_451 bl[451] br[451] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_452 bl[452] br[452] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_453 bl[453] br[453] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_454 bl[454] br[454] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_455 bl[455] br[455] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_456 bl[456] br[456] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_457 bl[457] br[457] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_458 bl[458] br[458] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_459 bl[459] br[459] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_460 bl[460] br[460] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_461 bl[461] br[461] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_462 bl[462] br[462] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_463 bl[463] br[463] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_464 bl[464] br[464] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_465 bl[465] br[465] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_466 bl[466] br[466] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_467 bl[467] br[467] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_468 bl[468] br[468] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_469 bl[469] br[469] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_470 bl[470] br[470] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_471 bl[471] br[471] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_472 bl[472] br[472] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_473 bl[473] br[473] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_474 bl[474] br[474] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_475 bl[475] br[475] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_476 bl[476] br[476] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_477 bl[477] br[477] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_478 bl[478] br[478] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_479 bl[479] br[479] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_480 bl[480] br[480] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_481 bl[481] br[481] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_482 bl[482] br[482] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_483 bl[483] br[483] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_484 bl[484] br[484] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_485 bl[485] br[485] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_486 bl[486] br[486] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_487 bl[487] br[487] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_488 bl[488] br[488] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_489 bl[489] br[489] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_490 bl[490] br[490] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_491 bl[491] br[491] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_492 bl[492] br[492] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_493 bl[493] br[493] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_494 bl[494] br[494] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_495 bl[495] br[495] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_496 bl[496] br[496] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_497 bl[497] br[497] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_498 bl[498] br[498] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_499 bl[499] br[499] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_500 bl[500] br[500] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_501 bl[501] br[501] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_502 bl[502] br[502] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_503 bl[503] br[503] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_504 bl[504] br[504] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_505 bl[505] br[505] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_506 bl[506] br[506] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_507 bl[507] br[507] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_508 bl[508] br[508] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_509 bl[509] br[509] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_510 bl[510] br[510] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_0_511 bl[511] br[511] vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xcell_1_0 bl[0] br[0] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_1 bl[1] br[1] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_2 bl[2] br[2] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_3 bl[3] br[3] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_4 bl[4] br[4] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_5 bl[5] br[5] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_6 bl[6] br[6] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_7 bl[7] br[7] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_8 bl[8] br[8] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_9 bl[9] br[9] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_10 bl[10] br[10] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_11 bl[11] br[11] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_12 bl[12] br[12] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_13 bl[13] br[13] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_14 bl[14] br[14] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_15 bl[15] br[15] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_16 bl[16] br[16] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_17 bl[17] br[17] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_18 bl[18] br[18] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_19 bl[19] br[19] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_20 bl[20] br[20] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_21 bl[21] br[21] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_22 bl[22] br[22] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_23 bl[23] br[23] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_24 bl[24] br[24] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_25 bl[25] br[25] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_26 bl[26] br[26] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_27 bl[27] br[27] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_28 bl[28] br[28] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_29 bl[29] br[29] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_30 bl[30] br[30] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_31 bl[31] br[31] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_32 bl[32] br[32] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_33 bl[33] br[33] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_34 bl[34] br[34] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_35 bl[35] br[35] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_36 bl[36] br[36] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_37 bl[37] br[37] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_38 bl[38] br[38] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_39 bl[39] br[39] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_40 bl[40] br[40] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_41 bl[41] br[41] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_42 bl[42] br[42] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_43 bl[43] br[43] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_44 bl[44] br[44] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_45 bl[45] br[45] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_46 bl[46] br[46] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_47 bl[47] br[47] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_48 bl[48] br[48] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_49 bl[49] br[49] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_50 bl[50] br[50] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_51 bl[51] br[51] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_52 bl[52] br[52] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_53 bl[53] br[53] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_54 bl[54] br[54] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_55 bl[55] br[55] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_56 bl[56] br[56] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_57 bl[57] br[57] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_58 bl[58] br[58] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_59 bl[59] br[59] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_60 bl[60] br[60] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_61 bl[61] br[61] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_62 bl[62] br[62] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_63 bl[63] br[63] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_64 bl[64] br[64] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_65 bl[65] br[65] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_66 bl[66] br[66] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_67 bl[67] br[67] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_68 bl[68] br[68] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_69 bl[69] br[69] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_70 bl[70] br[70] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_71 bl[71] br[71] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_72 bl[72] br[72] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_73 bl[73] br[73] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_74 bl[74] br[74] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_75 bl[75] br[75] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_76 bl[76] br[76] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_77 bl[77] br[77] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_78 bl[78] br[78] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_79 bl[79] br[79] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_80 bl[80] br[80] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_81 bl[81] br[81] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_82 bl[82] br[82] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_83 bl[83] br[83] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_84 bl[84] br[84] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_85 bl[85] br[85] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_86 bl[86] br[86] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_87 bl[87] br[87] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_88 bl[88] br[88] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_89 bl[89] br[89] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_90 bl[90] br[90] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_91 bl[91] br[91] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_92 bl[92] br[92] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_93 bl[93] br[93] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_94 bl[94] br[94] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_95 bl[95] br[95] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_96 bl[96] br[96] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_97 bl[97] br[97] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_98 bl[98] br[98] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_99 bl[99] br[99] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_100 bl[100] br[100] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_101 bl[101] br[101] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_102 bl[102] br[102] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_103 bl[103] br[103] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_104 bl[104] br[104] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_105 bl[105] br[105] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_106 bl[106] br[106] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_107 bl[107] br[107] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_108 bl[108] br[108] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_109 bl[109] br[109] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_110 bl[110] br[110] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_111 bl[111] br[111] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_112 bl[112] br[112] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_113 bl[113] br[113] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_114 bl[114] br[114] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_115 bl[115] br[115] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_116 bl[116] br[116] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_117 bl[117] br[117] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_118 bl[118] br[118] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_119 bl[119] br[119] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_120 bl[120] br[120] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_121 bl[121] br[121] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_122 bl[122] br[122] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_123 bl[123] br[123] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_124 bl[124] br[124] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_125 bl[125] br[125] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_126 bl[126] br[126] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_127 bl[127] br[127] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_128 bl[128] br[128] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_129 bl[129] br[129] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_130 bl[130] br[130] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_131 bl[131] br[131] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_132 bl[132] br[132] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_133 bl[133] br[133] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_134 bl[134] br[134] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_135 bl[135] br[135] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_136 bl[136] br[136] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_137 bl[137] br[137] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_138 bl[138] br[138] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_139 bl[139] br[139] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_140 bl[140] br[140] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_141 bl[141] br[141] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_142 bl[142] br[142] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_143 bl[143] br[143] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_144 bl[144] br[144] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_145 bl[145] br[145] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_146 bl[146] br[146] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_147 bl[147] br[147] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_148 bl[148] br[148] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_149 bl[149] br[149] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_150 bl[150] br[150] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_151 bl[151] br[151] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_152 bl[152] br[152] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_153 bl[153] br[153] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_154 bl[154] br[154] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_155 bl[155] br[155] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_156 bl[156] br[156] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_157 bl[157] br[157] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_158 bl[158] br[158] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_159 bl[159] br[159] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_160 bl[160] br[160] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_161 bl[161] br[161] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_162 bl[162] br[162] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_163 bl[163] br[163] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_164 bl[164] br[164] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_165 bl[165] br[165] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_166 bl[166] br[166] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_167 bl[167] br[167] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_168 bl[168] br[168] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_169 bl[169] br[169] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_170 bl[170] br[170] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_171 bl[171] br[171] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_172 bl[172] br[172] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_173 bl[173] br[173] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_174 bl[174] br[174] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_175 bl[175] br[175] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_176 bl[176] br[176] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_177 bl[177] br[177] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_178 bl[178] br[178] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_179 bl[179] br[179] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_180 bl[180] br[180] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_181 bl[181] br[181] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_182 bl[182] br[182] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_183 bl[183] br[183] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_184 bl[184] br[184] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_185 bl[185] br[185] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_186 bl[186] br[186] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_187 bl[187] br[187] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_188 bl[188] br[188] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_189 bl[189] br[189] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_190 bl[190] br[190] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_191 bl[191] br[191] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_192 bl[192] br[192] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_193 bl[193] br[193] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_194 bl[194] br[194] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_195 bl[195] br[195] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_196 bl[196] br[196] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_197 bl[197] br[197] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_198 bl[198] br[198] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_199 bl[199] br[199] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_200 bl[200] br[200] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_201 bl[201] br[201] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_202 bl[202] br[202] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_203 bl[203] br[203] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_204 bl[204] br[204] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_205 bl[205] br[205] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_206 bl[206] br[206] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_207 bl[207] br[207] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_208 bl[208] br[208] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_209 bl[209] br[209] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_210 bl[210] br[210] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_211 bl[211] br[211] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_212 bl[212] br[212] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_213 bl[213] br[213] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_214 bl[214] br[214] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_215 bl[215] br[215] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_216 bl[216] br[216] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_217 bl[217] br[217] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_218 bl[218] br[218] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_219 bl[219] br[219] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_220 bl[220] br[220] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_221 bl[221] br[221] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_222 bl[222] br[222] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_223 bl[223] br[223] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_224 bl[224] br[224] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_225 bl[225] br[225] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_226 bl[226] br[226] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_227 bl[227] br[227] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_228 bl[228] br[228] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_229 bl[229] br[229] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_230 bl[230] br[230] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_231 bl[231] br[231] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_232 bl[232] br[232] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_233 bl[233] br[233] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_234 bl[234] br[234] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_235 bl[235] br[235] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_236 bl[236] br[236] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_237 bl[237] br[237] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_238 bl[238] br[238] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_239 bl[239] br[239] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_240 bl[240] br[240] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_241 bl[241] br[241] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_242 bl[242] br[242] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_243 bl[243] br[243] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_244 bl[244] br[244] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_245 bl[245] br[245] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_246 bl[246] br[246] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_247 bl[247] br[247] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_248 bl[248] br[248] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_249 bl[249] br[249] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_250 bl[250] br[250] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_251 bl[251] br[251] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_252 bl[252] br[252] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_253 bl[253] br[253] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_254 bl[254] br[254] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_255 bl[255] br[255] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_256 bl[256] br[256] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_257 bl[257] br[257] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_258 bl[258] br[258] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_259 bl[259] br[259] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_260 bl[260] br[260] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_261 bl[261] br[261] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_262 bl[262] br[262] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_263 bl[263] br[263] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_264 bl[264] br[264] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_265 bl[265] br[265] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_266 bl[266] br[266] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_267 bl[267] br[267] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_268 bl[268] br[268] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_269 bl[269] br[269] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_270 bl[270] br[270] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_271 bl[271] br[271] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_272 bl[272] br[272] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_273 bl[273] br[273] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_274 bl[274] br[274] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_275 bl[275] br[275] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_276 bl[276] br[276] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_277 bl[277] br[277] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_278 bl[278] br[278] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_279 bl[279] br[279] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_280 bl[280] br[280] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_281 bl[281] br[281] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_282 bl[282] br[282] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_283 bl[283] br[283] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_284 bl[284] br[284] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_285 bl[285] br[285] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_286 bl[286] br[286] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_287 bl[287] br[287] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_288 bl[288] br[288] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_289 bl[289] br[289] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_290 bl[290] br[290] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_291 bl[291] br[291] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_292 bl[292] br[292] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_293 bl[293] br[293] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_294 bl[294] br[294] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_295 bl[295] br[295] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_296 bl[296] br[296] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_297 bl[297] br[297] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_298 bl[298] br[298] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_299 bl[299] br[299] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_300 bl[300] br[300] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_301 bl[301] br[301] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_302 bl[302] br[302] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_303 bl[303] br[303] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_304 bl[304] br[304] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_305 bl[305] br[305] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_306 bl[306] br[306] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_307 bl[307] br[307] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_308 bl[308] br[308] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_309 bl[309] br[309] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_310 bl[310] br[310] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_311 bl[311] br[311] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_312 bl[312] br[312] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_313 bl[313] br[313] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_314 bl[314] br[314] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_315 bl[315] br[315] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_316 bl[316] br[316] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_317 bl[317] br[317] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_318 bl[318] br[318] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_319 bl[319] br[319] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_320 bl[320] br[320] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_321 bl[321] br[321] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_322 bl[322] br[322] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_323 bl[323] br[323] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_324 bl[324] br[324] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_325 bl[325] br[325] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_326 bl[326] br[326] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_327 bl[327] br[327] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_328 bl[328] br[328] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_329 bl[329] br[329] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_330 bl[330] br[330] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_331 bl[331] br[331] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_332 bl[332] br[332] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_333 bl[333] br[333] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_334 bl[334] br[334] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_335 bl[335] br[335] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_336 bl[336] br[336] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_337 bl[337] br[337] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_338 bl[338] br[338] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_339 bl[339] br[339] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_340 bl[340] br[340] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_341 bl[341] br[341] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_342 bl[342] br[342] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_343 bl[343] br[343] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_344 bl[344] br[344] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_345 bl[345] br[345] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_346 bl[346] br[346] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_347 bl[347] br[347] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_348 bl[348] br[348] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_349 bl[349] br[349] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_350 bl[350] br[350] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_351 bl[351] br[351] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_352 bl[352] br[352] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_353 bl[353] br[353] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_354 bl[354] br[354] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_355 bl[355] br[355] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_356 bl[356] br[356] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_357 bl[357] br[357] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_358 bl[358] br[358] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_359 bl[359] br[359] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_360 bl[360] br[360] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_361 bl[361] br[361] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_362 bl[362] br[362] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_363 bl[363] br[363] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_364 bl[364] br[364] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_365 bl[365] br[365] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_366 bl[366] br[366] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_367 bl[367] br[367] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_368 bl[368] br[368] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_369 bl[369] br[369] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_370 bl[370] br[370] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_371 bl[371] br[371] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_372 bl[372] br[372] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_373 bl[373] br[373] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_374 bl[374] br[374] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_375 bl[375] br[375] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_376 bl[376] br[376] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_377 bl[377] br[377] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_378 bl[378] br[378] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_379 bl[379] br[379] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_380 bl[380] br[380] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_381 bl[381] br[381] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_382 bl[382] br[382] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_383 bl[383] br[383] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_384 bl[384] br[384] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_385 bl[385] br[385] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_386 bl[386] br[386] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_387 bl[387] br[387] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_388 bl[388] br[388] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_389 bl[389] br[389] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_390 bl[390] br[390] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_391 bl[391] br[391] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_392 bl[392] br[392] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_393 bl[393] br[393] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_394 bl[394] br[394] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_395 bl[395] br[395] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_396 bl[396] br[396] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_397 bl[397] br[397] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_398 bl[398] br[398] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_399 bl[399] br[399] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_400 bl[400] br[400] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_401 bl[401] br[401] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_402 bl[402] br[402] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_403 bl[403] br[403] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_404 bl[404] br[404] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_405 bl[405] br[405] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_406 bl[406] br[406] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_407 bl[407] br[407] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_408 bl[408] br[408] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_409 bl[409] br[409] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_410 bl[410] br[410] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_411 bl[411] br[411] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_412 bl[412] br[412] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_413 bl[413] br[413] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_414 bl[414] br[414] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_415 bl[415] br[415] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_416 bl[416] br[416] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_417 bl[417] br[417] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_418 bl[418] br[418] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_419 bl[419] br[419] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_420 bl[420] br[420] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_421 bl[421] br[421] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_422 bl[422] br[422] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_423 bl[423] br[423] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_424 bl[424] br[424] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_425 bl[425] br[425] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_426 bl[426] br[426] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_427 bl[427] br[427] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_428 bl[428] br[428] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_429 bl[429] br[429] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_430 bl[430] br[430] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_431 bl[431] br[431] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_432 bl[432] br[432] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_433 bl[433] br[433] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_434 bl[434] br[434] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_435 bl[435] br[435] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_436 bl[436] br[436] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_437 bl[437] br[437] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_438 bl[438] br[438] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_439 bl[439] br[439] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_440 bl[440] br[440] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_441 bl[441] br[441] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_442 bl[442] br[442] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_443 bl[443] br[443] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_444 bl[444] br[444] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_445 bl[445] br[445] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_446 bl[446] br[446] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_447 bl[447] br[447] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_448 bl[448] br[448] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_449 bl[449] br[449] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_450 bl[450] br[450] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_451 bl[451] br[451] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_452 bl[452] br[452] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_453 bl[453] br[453] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_454 bl[454] br[454] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_455 bl[455] br[455] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_456 bl[456] br[456] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_457 bl[457] br[457] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_458 bl[458] br[458] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_459 bl[459] br[459] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_460 bl[460] br[460] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_461 bl[461] br[461] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_462 bl[462] br[462] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_463 bl[463] br[463] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_464 bl[464] br[464] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_465 bl[465] br[465] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_466 bl[466] br[466] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_467 bl[467] br[467] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_468 bl[468] br[468] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_469 bl[469] br[469] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_470 bl[470] br[470] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_471 bl[471] br[471] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_472 bl[472] br[472] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_473 bl[473] br[473] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_474 bl[474] br[474] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_475 bl[475] br[475] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_476 bl[476] br[476] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_477 bl[477] br[477] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_478 bl[478] br[478] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_479 bl[479] br[479] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_480 bl[480] br[480] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_481 bl[481] br[481] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_482 bl[482] br[482] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_483 bl[483] br[483] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_484 bl[484] br[484] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_485 bl[485] br[485] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_486 bl[486] br[486] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_487 bl[487] br[487] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_488 bl[488] br[488] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_489 bl[489] br[489] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_490 bl[490] br[490] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_491 bl[491] br[491] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_492 bl[492] br[492] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_493 bl[493] br[493] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_494 bl[494] br[494] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_495 bl[495] br[495] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_496 bl[496] br[496] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_497 bl[497] br[497] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_498 bl[498] br[498] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_499 bl[499] br[499] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_500 bl[500] br[500] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_501 bl[501] br[501] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_502 bl[502] br[502] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_503 bl[503] br[503] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_504 bl[504] br[504] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_505 bl[505] br[505] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_506 bl[506] br[506] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_507 bl[507] br[507] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_508 bl[508] br[508] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_509 bl[509] br[509] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_510 bl[510] br[510] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_1_511 bl[511] br[511] vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xcell_2_0 bl[0] br[0] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_1 bl[1] br[1] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_2 bl[2] br[2] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_3 bl[3] br[3] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_4 bl[4] br[4] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_5 bl[5] br[5] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_6 bl[6] br[6] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_7 bl[7] br[7] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_8 bl[8] br[8] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_9 bl[9] br[9] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_10 bl[10] br[10] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_11 bl[11] br[11] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_12 bl[12] br[12] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_13 bl[13] br[13] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_14 bl[14] br[14] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_15 bl[15] br[15] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_16 bl[16] br[16] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_17 bl[17] br[17] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_18 bl[18] br[18] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_19 bl[19] br[19] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_20 bl[20] br[20] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_21 bl[21] br[21] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_22 bl[22] br[22] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_23 bl[23] br[23] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_24 bl[24] br[24] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_25 bl[25] br[25] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_26 bl[26] br[26] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_27 bl[27] br[27] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_28 bl[28] br[28] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_29 bl[29] br[29] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_30 bl[30] br[30] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_31 bl[31] br[31] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_32 bl[32] br[32] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_33 bl[33] br[33] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_34 bl[34] br[34] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_35 bl[35] br[35] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_36 bl[36] br[36] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_37 bl[37] br[37] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_38 bl[38] br[38] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_39 bl[39] br[39] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_40 bl[40] br[40] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_41 bl[41] br[41] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_42 bl[42] br[42] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_43 bl[43] br[43] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_44 bl[44] br[44] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_45 bl[45] br[45] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_46 bl[46] br[46] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_47 bl[47] br[47] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_48 bl[48] br[48] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_49 bl[49] br[49] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_50 bl[50] br[50] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_51 bl[51] br[51] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_52 bl[52] br[52] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_53 bl[53] br[53] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_54 bl[54] br[54] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_55 bl[55] br[55] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_56 bl[56] br[56] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_57 bl[57] br[57] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_58 bl[58] br[58] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_59 bl[59] br[59] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_60 bl[60] br[60] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_61 bl[61] br[61] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_62 bl[62] br[62] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_63 bl[63] br[63] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_64 bl[64] br[64] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_65 bl[65] br[65] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_66 bl[66] br[66] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_67 bl[67] br[67] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_68 bl[68] br[68] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_69 bl[69] br[69] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_70 bl[70] br[70] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_71 bl[71] br[71] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_72 bl[72] br[72] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_73 bl[73] br[73] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_74 bl[74] br[74] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_75 bl[75] br[75] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_76 bl[76] br[76] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_77 bl[77] br[77] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_78 bl[78] br[78] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_79 bl[79] br[79] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_80 bl[80] br[80] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_81 bl[81] br[81] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_82 bl[82] br[82] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_83 bl[83] br[83] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_84 bl[84] br[84] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_85 bl[85] br[85] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_86 bl[86] br[86] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_87 bl[87] br[87] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_88 bl[88] br[88] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_89 bl[89] br[89] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_90 bl[90] br[90] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_91 bl[91] br[91] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_92 bl[92] br[92] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_93 bl[93] br[93] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_94 bl[94] br[94] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_95 bl[95] br[95] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_96 bl[96] br[96] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_97 bl[97] br[97] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_98 bl[98] br[98] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_99 bl[99] br[99] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_100 bl[100] br[100] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_101 bl[101] br[101] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_102 bl[102] br[102] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_103 bl[103] br[103] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_104 bl[104] br[104] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_105 bl[105] br[105] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_106 bl[106] br[106] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_107 bl[107] br[107] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_108 bl[108] br[108] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_109 bl[109] br[109] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_110 bl[110] br[110] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_111 bl[111] br[111] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_112 bl[112] br[112] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_113 bl[113] br[113] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_114 bl[114] br[114] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_115 bl[115] br[115] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_116 bl[116] br[116] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_117 bl[117] br[117] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_118 bl[118] br[118] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_119 bl[119] br[119] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_120 bl[120] br[120] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_121 bl[121] br[121] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_122 bl[122] br[122] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_123 bl[123] br[123] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_124 bl[124] br[124] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_125 bl[125] br[125] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_126 bl[126] br[126] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_127 bl[127] br[127] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_128 bl[128] br[128] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_129 bl[129] br[129] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_130 bl[130] br[130] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_131 bl[131] br[131] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_132 bl[132] br[132] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_133 bl[133] br[133] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_134 bl[134] br[134] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_135 bl[135] br[135] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_136 bl[136] br[136] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_137 bl[137] br[137] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_138 bl[138] br[138] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_139 bl[139] br[139] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_140 bl[140] br[140] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_141 bl[141] br[141] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_142 bl[142] br[142] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_143 bl[143] br[143] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_144 bl[144] br[144] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_145 bl[145] br[145] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_146 bl[146] br[146] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_147 bl[147] br[147] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_148 bl[148] br[148] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_149 bl[149] br[149] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_150 bl[150] br[150] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_151 bl[151] br[151] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_152 bl[152] br[152] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_153 bl[153] br[153] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_154 bl[154] br[154] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_155 bl[155] br[155] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_156 bl[156] br[156] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_157 bl[157] br[157] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_158 bl[158] br[158] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_159 bl[159] br[159] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_160 bl[160] br[160] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_161 bl[161] br[161] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_162 bl[162] br[162] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_163 bl[163] br[163] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_164 bl[164] br[164] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_165 bl[165] br[165] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_166 bl[166] br[166] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_167 bl[167] br[167] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_168 bl[168] br[168] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_169 bl[169] br[169] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_170 bl[170] br[170] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_171 bl[171] br[171] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_172 bl[172] br[172] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_173 bl[173] br[173] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_174 bl[174] br[174] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_175 bl[175] br[175] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_176 bl[176] br[176] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_177 bl[177] br[177] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_178 bl[178] br[178] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_179 bl[179] br[179] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_180 bl[180] br[180] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_181 bl[181] br[181] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_182 bl[182] br[182] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_183 bl[183] br[183] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_184 bl[184] br[184] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_185 bl[185] br[185] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_186 bl[186] br[186] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_187 bl[187] br[187] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_188 bl[188] br[188] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_189 bl[189] br[189] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_190 bl[190] br[190] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_191 bl[191] br[191] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_192 bl[192] br[192] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_193 bl[193] br[193] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_194 bl[194] br[194] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_195 bl[195] br[195] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_196 bl[196] br[196] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_197 bl[197] br[197] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_198 bl[198] br[198] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_199 bl[199] br[199] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_200 bl[200] br[200] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_201 bl[201] br[201] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_202 bl[202] br[202] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_203 bl[203] br[203] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_204 bl[204] br[204] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_205 bl[205] br[205] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_206 bl[206] br[206] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_207 bl[207] br[207] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_208 bl[208] br[208] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_209 bl[209] br[209] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_210 bl[210] br[210] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_211 bl[211] br[211] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_212 bl[212] br[212] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_213 bl[213] br[213] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_214 bl[214] br[214] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_215 bl[215] br[215] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_216 bl[216] br[216] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_217 bl[217] br[217] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_218 bl[218] br[218] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_219 bl[219] br[219] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_220 bl[220] br[220] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_221 bl[221] br[221] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_222 bl[222] br[222] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_223 bl[223] br[223] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_224 bl[224] br[224] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_225 bl[225] br[225] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_226 bl[226] br[226] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_227 bl[227] br[227] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_228 bl[228] br[228] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_229 bl[229] br[229] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_230 bl[230] br[230] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_231 bl[231] br[231] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_232 bl[232] br[232] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_233 bl[233] br[233] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_234 bl[234] br[234] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_235 bl[235] br[235] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_236 bl[236] br[236] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_237 bl[237] br[237] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_238 bl[238] br[238] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_239 bl[239] br[239] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_240 bl[240] br[240] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_241 bl[241] br[241] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_242 bl[242] br[242] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_243 bl[243] br[243] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_244 bl[244] br[244] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_245 bl[245] br[245] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_246 bl[246] br[246] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_247 bl[247] br[247] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_248 bl[248] br[248] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_249 bl[249] br[249] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_250 bl[250] br[250] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_251 bl[251] br[251] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_252 bl[252] br[252] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_253 bl[253] br[253] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_254 bl[254] br[254] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_255 bl[255] br[255] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_256 bl[256] br[256] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_257 bl[257] br[257] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_258 bl[258] br[258] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_259 bl[259] br[259] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_260 bl[260] br[260] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_261 bl[261] br[261] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_262 bl[262] br[262] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_263 bl[263] br[263] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_264 bl[264] br[264] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_265 bl[265] br[265] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_266 bl[266] br[266] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_267 bl[267] br[267] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_268 bl[268] br[268] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_269 bl[269] br[269] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_270 bl[270] br[270] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_271 bl[271] br[271] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_272 bl[272] br[272] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_273 bl[273] br[273] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_274 bl[274] br[274] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_275 bl[275] br[275] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_276 bl[276] br[276] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_277 bl[277] br[277] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_278 bl[278] br[278] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_279 bl[279] br[279] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_280 bl[280] br[280] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_281 bl[281] br[281] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_282 bl[282] br[282] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_283 bl[283] br[283] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_284 bl[284] br[284] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_285 bl[285] br[285] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_286 bl[286] br[286] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_287 bl[287] br[287] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_288 bl[288] br[288] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_289 bl[289] br[289] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_290 bl[290] br[290] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_291 bl[291] br[291] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_292 bl[292] br[292] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_293 bl[293] br[293] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_294 bl[294] br[294] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_295 bl[295] br[295] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_296 bl[296] br[296] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_297 bl[297] br[297] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_298 bl[298] br[298] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_299 bl[299] br[299] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_300 bl[300] br[300] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_301 bl[301] br[301] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_302 bl[302] br[302] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_303 bl[303] br[303] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_304 bl[304] br[304] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_305 bl[305] br[305] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_306 bl[306] br[306] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_307 bl[307] br[307] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_308 bl[308] br[308] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_309 bl[309] br[309] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_310 bl[310] br[310] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_311 bl[311] br[311] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_312 bl[312] br[312] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_313 bl[313] br[313] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_314 bl[314] br[314] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_315 bl[315] br[315] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_316 bl[316] br[316] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_317 bl[317] br[317] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_318 bl[318] br[318] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_319 bl[319] br[319] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_320 bl[320] br[320] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_321 bl[321] br[321] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_322 bl[322] br[322] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_323 bl[323] br[323] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_324 bl[324] br[324] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_325 bl[325] br[325] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_326 bl[326] br[326] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_327 bl[327] br[327] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_328 bl[328] br[328] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_329 bl[329] br[329] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_330 bl[330] br[330] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_331 bl[331] br[331] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_332 bl[332] br[332] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_333 bl[333] br[333] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_334 bl[334] br[334] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_335 bl[335] br[335] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_336 bl[336] br[336] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_337 bl[337] br[337] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_338 bl[338] br[338] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_339 bl[339] br[339] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_340 bl[340] br[340] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_341 bl[341] br[341] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_342 bl[342] br[342] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_343 bl[343] br[343] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_344 bl[344] br[344] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_345 bl[345] br[345] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_346 bl[346] br[346] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_347 bl[347] br[347] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_348 bl[348] br[348] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_349 bl[349] br[349] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_350 bl[350] br[350] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_351 bl[351] br[351] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_352 bl[352] br[352] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_353 bl[353] br[353] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_354 bl[354] br[354] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_355 bl[355] br[355] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_356 bl[356] br[356] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_357 bl[357] br[357] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_358 bl[358] br[358] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_359 bl[359] br[359] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_360 bl[360] br[360] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_361 bl[361] br[361] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_362 bl[362] br[362] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_363 bl[363] br[363] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_364 bl[364] br[364] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_365 bl[365] br[365] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_366 bl[366] br[366] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_367 bl[367] br[367] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_368 bl[368] br[368] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_369 bl[369] br[369] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_370 bl[370] br[370] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_371 bl[371] br[371] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_372 bl[372] br[372] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_373 bl[373] br[373] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_374 bl[374] br[374] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_375 bl[375] br[375] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_376 bl[376] br[376] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_377 bl[377] br[377] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_378 bl[378] br[378] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_379 bl[379] br[379] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_380 bl[380] br[380] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_381 bl[381] br[381] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_382 bl[382] br[382] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_383 bl[383] br[383] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_384 bl[384] br[384] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_385 bl[385] br[385] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_386 bl[386] br[386] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_387 bl[387] br[387] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_388 bl[388] br[388] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_389 bl[389] br[389] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_390 bl[390] br[390] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_391 bl[391] br[391] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_392 bl[392] br[392] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_393 bl[393] br[393] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_394 bl[394] br[394] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_395 bl[395] br[395] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_396 bl[396] br[396] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_397 bl[397] br[397] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_398 bl[398] br[398] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_399 bl[399] br[399] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_400 bl[400] br[400] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_401 bl[401] br[401] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_402 bl[402] br[402] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_403 bl[403] br[403] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_404 bl[404] br[404] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_405 bl[405] br[405] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_406 bl[406] br[406] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_407 bl[407] br[407] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_408 bl[408] br[408] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_409 bl[409] br[409] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_410 bl[410] br[410] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_411 bl[411] br[411] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_412 bl[412] br[412] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_413 bl[413] br[413] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_414 bl[414] br[414] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_415 bl[415] br[415] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_416 bl[416] br[416] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_417 bl[417] br[417] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_418 bl[418] br[418] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_419 bl[419] br[419] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_420 bl[420] br[420] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_421 bl[421] br[421] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_422 bl[422] br[422] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_423 bl[423] br[423] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_424 bl[424] br[424] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_425 bl[425] br[425] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_426 bl[426] br[426] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_427 bl[427] br[427] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_428 bl[428] br[428] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_429 bl[429] br[429] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_430 bl[430] br[430] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_431 bl[431] br[431] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_432 bl[432] br[432] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_433 bl[433] br[433] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_434 bl[434] br[434] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_435 bl[435] br[435] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_436 bl[436] br[436] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_437 bl[437] br[437] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_438 bl[438] br[438] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_439 bl[439] br[439] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_440 bl[440] br[440] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_441 bl[441] br[441] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_442 bl[442] br[442] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_443 bl[443] br[443] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_444 bl[444] br[444] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_445 bl[445] br[445] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_446 bl[446] br[446] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_447 bl[447] br[447] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_448 bl[448] br[448] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_449 bl[449] br[449] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_450 bl[450] br[450] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_451 bl[451] br[451] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_452 bl[452] br[452] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_453 bl[453] br[453] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_454 bl[454] br[454] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_455 bl[455] br[455] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_456 bl[456] br[456] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_457 bl[457] br[457] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_458 bl[458] br[458] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_459 bl[459] br[459] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_460 bl[460] br[460] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_461 bl[461] br[461] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_462 bl[462] br[462] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_463 bl[463] br[463] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_464 bl[464] br[464] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_465 bl[465] br[465] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_466 bl[466] br[466] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_467 bl[467] br[467] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_468 bl[468] br[468] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_469 bl[469] br[469] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_470 bl[470] br[470] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_471 bl[471] br[471] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_472 bl[472] br[472] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_473 bl[473] br[473] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_474 bl[474] br[474] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_475 bl[475] br[475] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_476 bl[476] br[476] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_477 bl[477] br[477] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_478 bl[478] br[478] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_479 bl[479] br[479] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_480 bl[480] br[480] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_481 bl[481] br[481] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_482 bl[482] br[482] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_483 bl[483] br[483] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_484 bl[484] br[484] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_485 bl[485] br[485] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_486 bl[486] br[486] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_487 bl[487] br[487] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_488 bl[488] br[488] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_489 bl[489] br[489] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_490 bl[490] br[490] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_491 bl[491] br[491] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_492 bl[492] br[492] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_493 bl[493] br[493] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_494 bl[494] br[494] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_495 bl[495] br[495] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_496 bl[496] br[496] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_497 bl[497] br[497] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_498 bl[498] br[498] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_499 bl[499] br[499] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_500 bl[500] br[500] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_501 bl[501] br[501] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_502 bl[502] br[502] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_503 bl[503] br[503] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_504 bl[504] br[504] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_505 bl[505] br[505] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_506 bl[506] br[506] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_507 bl[507] br[507] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_508 bl[508] br[508] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_509 bl[509] br[509] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_510 bl[510] br[510] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_2_511 bl[511] br[511] vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xcell_3_0 bl[0] br[0] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_1 bl[1] br[1] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_2 bl[2] br[2] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_3 bl[3] br[3] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_4 bl[4] br[4] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_5 bl[5] br[5] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_6 bl[6] br[6] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_7 bl[7] br[7] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_8 bl[8] br[8] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_9 bl[9] br[9] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_10 bl[10] br[10] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_11 bl[11] br[11] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_12 bl[12] br[12] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_13 bl[13] br[13] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_14 bl[14] br[14] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_15 bl[15] br[15] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_16 bl[16] br[16] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_17 bl[17] br[17] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_18 bl[18] br[18] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_19 bl[19] br[19] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_20 bl[20] br[20] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_21 bl[21] br[21] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_22 bl[22] br[22] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_23 bl[23] br[23] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_24 bl[24] br[24] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_25 bl[25] br[25] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_26 bl[26] br[26] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_27 bl[27] br[27] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_28 bl[28] br[28] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_29 bl[29] br[29] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_30 bl[30] br[30] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_31 bl[31] br[31] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_32 bl[32] br[32] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_33 bl[33] br[33] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_34 bl[34] br[34] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_35 bl[35] br[35] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_36 bl[36] br[36] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_37 bl[37] br[37] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_38 bl[38] br[38] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_39 bl[39] br[39] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_40 bl[40] br[40] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_41 bl[41] br[41] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_42 bl[42] br[42] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_43 bl[43] br[43] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_44 bl[44] br[44] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_45 bl[45] br[45] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_46 bl[46] br[46] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_47 bl[47] br[47] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_48 bl[48] br[48] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_49 bl[49] br[49] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_50 bl[50] br[50] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_51 bl[51] br[51] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_52 bl[52] br[52] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_53 bl[53] br[53] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_54 bl[54] br[54] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_55 bl[55] br[55] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_56 bl[56] br[56] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_57 bl[57] br[57] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_58 bl[58] br[58] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_59 bl[59] br[59] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_60 bl[60] br[60] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_61 bl[61] br[61] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_62 bl[62] br[62] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_63 bl[63] br[63] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_64 bl[64] br[64] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_65 bl[65] br[65] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_66 bl[66] br[66] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_67 bl[67] br[67] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_68 bl[68] br[68] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_69 bl[69] br[69] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_70 bl[70] br[70] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_71 bl[71] br[71] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_72 bl[72] br[72] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_73 bl[73] br[73] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_74 bl[74] br[74] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_75 bl[75] br[75] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_76 bl[76] br[76] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_77 bl[77] br[77] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_78 bl[78] br[78] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_79 bl[79] br[79] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_80 bl[80] br[80] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_81 bl[81] br[81] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_82 bl[82] br[82] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_83 bl[83] br[83] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_84 bl[84] br[84] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_85 bl[85] br[85] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_86 bl[86] br[86] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_87 bl[87] br[87] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_88 bl[88] br[88] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_89 bl[89] br[89] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_90 bl[90] br[90] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_91 bl[91] br[91] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_92 bl[92] br[92] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_93 bl[93] br[93] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_94 bl[94] br[94] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_95 bl[95] br[95] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_96 bl[96] br[96] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_97 bl[97] br[97] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_98 bl[98] br[98] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_99 bl[99] br[99] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_100 bl[100] br[100] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_101 bl[101] br[101] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_102 bl[102] br[102] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_103 bl[103] br[103] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_104 bl[104] br[104] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_105 bl[105] br[105] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_106 bl[106] br[106] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_107 bl[107] br[107] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_108 bl[108] br[108] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_109 bl[109] br[109] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_110 bl[110] br[110] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_111 bl[111] br[111] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_112 bl[112] br[112] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_113 bl[113] br[113] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_114 bl[114] br[114] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_115 bl[115] br[115] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_116 bl[116] br[116] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_117 bl[117] br[117] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_118 bl[118] br[118] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_119 bl[119] br[119] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_120 bl[120] br[120] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_121 bl[121] br[121] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_122 bl[122] br[122] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_123 bl[123] br[123] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_124 bl[124] br[124] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_125 bl[125] br[125] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_126 bl[126] br[126] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_127 bl[127] br[127] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_128 bl[128] br[128] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_129 bl[129] br[129] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_130 bl[130] br[130] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_131 bl[131] br[131] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_132 bl[132] br[132] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_133 bl[133] br[133] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_134 bl[134] br[134] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_135 bl[135] br[135] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_136 bl[136] br[136] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_137 bl[137] br[137] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_138 bl[138] br[138] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_139 bl[139] br[139] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_140 bl[140] br[140] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_141 bl[141] br[141] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_142 bl[142] br[142] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_143 bl[143] br[143] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_144 bl[144] br[144] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_145 bl[145] br[145] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_146 bl[146] br[146] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_147 bl[147] br[147] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_148 bl[148] br[148] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_149 bl[149] br[149] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_150 bl[150] br[150] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_151 bl[151] br[151] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_152 bl[152] br[152] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_153 bl[153] br[153] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_154 bl[154] br[154] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_155 bl[155] br[155] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_156 bl[156] br[156] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_157 bl[157] br[157] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_158 bl[158] br[158] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_159 bl[159] br[159] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_160 bl[160] br[160] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_161 bl[161] br[161] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_162 bl[162] br[162] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_163 bl[163] br[163] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_164 bl[164] br[164] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_165 bl[165] br[165] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_166 bl[166] br[166] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_167 bl[167] br[167] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_168 bl[168] br[168] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_169 bl[169] br[169] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_170 bl[170] br[170] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_171 bl[171] br[171] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_172 bl[172] br[172] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_173 bl[173] br[173] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_174 bl[174] br[174] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_175 bl[175] br[175] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_176 bl[176] br[176] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_177 bl[177] br[177] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_178 bl[178] br[178] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_179 bl[179] br[179] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_180 bl[180] br[180] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_181 bl[181] br[181] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_182 bl[182] br[182] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_183 bl[183] br[183] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_184 bl[184] br[184] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_185 bl[185] br[185] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_186 bl[186] br[186] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_187 bl[187] br[187] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_188 bl[188] br[188] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_189 bl[189] br[189] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_190 bl[190] br[190] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_191 bl[191] br[191] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_192 bl[192] br[192] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_193 bl[193] br[193] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_194 bl[194] br[194] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_195 bl[195] br[195] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_196 bl[196] br[196] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_197 bl[197] br[197] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_198 bl[198] br[198] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_199 bl[199] br[199] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_200 bl[200] br[200] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_201 bl[201] br[201] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_202 bl[202] br[202] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_203 bl[203] br[203] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_204 bl[204] br[204] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_205 bl[205] br[205] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_206 bl[206] br[206] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_207 bl[207] br[207] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_208 bl[208] br[208] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_209 bl[209] br[209] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_210 bl[210] br[210] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_211 bl[211] br[211] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_212 bl[212] br[212] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_213 bl[213] br[213] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_214 bl[214] br[214] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_215 bl[215] br[215] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_216 bl[216] br[216] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_217 bl[217] br[217] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_218 bl[218] br[218] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_219 bl[219] br[219] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_220 bl[220] br[220] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_221 bl[221] br[221] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_222 bl[222] br[222] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_223 bl[223] br[223] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_224 bl[224] br[224] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_225 bl[225] br[225] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_226 bl[226] br[226] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_227 bl[227] br[227] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_228 bl[228] br[228] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_229 bl[229] br[229] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_230 bl[230] br[230] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_231 bl[231] br[231] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_232 bl[232] br[232] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_233 bl[233] br[233] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_234 bl[234] br[234] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_235 bl[235] br[235] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_236 bl[236] br[236] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_237 bl[237] br[237] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_238 bl[238] br[238] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_239 bl[239] br[239] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_240 bl[240] br[240] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_241 bl[241] br[241] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_242 bl[242] br[242] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_243 bl[243] br[243] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_244 bl[244] br[244] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_245 bl[245] br[245] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_246 bl[246] br[246] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_247 bl[247] br[247] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_248 bl[248] br[248] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_249 bl[249] br[249] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_250 bl[250] br[250] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_251 bl[251] br[251] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_252 bl[252] br[252] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_253 bl[253] br[253] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_254 bl[254] br[254] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_255 bl[255] br[255] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_256 bl[256] br[256] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_257 bl[257] br[257] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_258 bl[258] br[258] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_259 bl[259] br[259] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_260 bl[260] br[260] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_261 bl[261] br[261] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_262 bl[262] br[262] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_263 bl[263] br[263] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_264 bl[264] br[264] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_265 bl[265] br[265] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_266 bl[266] br[266] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_267 bl[267] br[267] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_268 bl[268] br[268] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_269 bl[269] br[269] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_270 bl[270] br[270] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_271 bl[271] br[271] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_272 bl[272] br[272] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_273 bl[273] br[273] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_274 bl[274] br[274] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_275 bl[275] br[275] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_276 bl[276] br[276] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_277 bl[277] br[277] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_278 bl[278] br[278] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_279 bl[279] br[279] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_280 bl[280] br[280] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_281 bl[281] br[281] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_282 bl[282] br[282] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_283 bl[283] br[283] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_284 bl[284] br[284] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_285 bl[285] br[285] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_286 bl[286] br[286] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_287 bl[287] br[287] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_288 bl[288] br[288] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_289 bl[289] br[289] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_290 bl[290] br[290] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_291 bl[291] br[291] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_292 bl[292] br[292] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_293 bl[293] br[293] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_294 bl[294] br[294] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_295 bl[295] br[295] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_296 bl[296] br[296] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_297 bl[297] br[297] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_298 bl[298] br[298] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_299 bl[299] br[299] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_300 bl[300] br[300] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_301 bl[301] br[301] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_302 bl[302] br[302] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_303 bl[303] br[303] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_304 bl[304] br[304] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_305 bl[305] br[305] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_306 bl[306] br[306] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_307 bl[307] br[307] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_308 bl[308] br[308] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_309 bl[309] br[309] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_310 bl[310] br[310] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_311 bl[311] br[311] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_312 bl[312] br[312] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_313 bl[313] br[313] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_314 bl[314] br[314] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_315 bl[315] br[315] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_316 bl[316] br[316] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_317 bl[317] br[317] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_318 bl[318] br[318] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_319 bl[319] br[319] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_320 bl[320] br[320] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_321 bl[321] br[321] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_322 bl[322] br[322] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_323 bl[323] br[323] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_324 bl[324] br[324] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_325 bl[325] br[325] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_326 bl[326] br[326] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_327 bl[327] br[327] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_328 bl[328] br[328] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_329 bl[329] br[329] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_330 bl[330] br[330] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_331 bl[331] br[331] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_332 bl[332] br[332] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_333 bl[333] br[333] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_334 bl[334] br[334] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_335 bl[335] br[335] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_336 bl[336] br[336] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_337 bl[337] br[337] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_338 bl[338] br[338] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_339 bl[339] br[339] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_340 bl[340] br[340] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_341 bl[341] br[341] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_342 bl[342] br[342] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_343 bl[343] br[343] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_344 bl[344] br[344] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_345 bl[345] br[345] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_346 bl[346] br[346] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_347 bl[347] br[347] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_348 bl[348] br[348] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_349 bl[349] br[349] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_350 bl[350] br[350] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_351 bl[351] br[351] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_352 bl[352] br[352] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_353 bl[353] br[353] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_354 bl[354] br[354] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_355 bl[355] br[355] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_356 bl[356] br[356] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_357 bl[357] br[357] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_358 bl[358] br[358] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_359 bl[359] br[359] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_360 bl[360] br[360] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_361 bl[361] br[361] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_362 bl[362] br[362] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_363 bl[363] br[363] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_364 bl[364] br[364] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_365 bl[365] br[365] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_366 bl[366] br[366] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_367 bl[367] br[367] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_368 bl[368] br[368] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_369 bl[369] br[369] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_370 bl[370] br[370] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_371 bl[371] br[371] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_372 bl[372] br[372] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_373 bl[373] br[373] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_374 bl[374] br[374] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_375 bl[375] br[375] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_376 bl[376] br[376] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_377 bl[377] br[377] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_378 bl[378] br[378] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_379 bl[379] br[379] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_380 bl[380] br[380] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_381 bl[381] br[381] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_382 bl[382] br[382] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_383 bl[383] br[383] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_384 bl[384] br[384] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_385 bl[385] br[385] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_386 bl[386] br[386] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_387 bl[387] br[387] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_388 bl[388] br[388] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_389 bl[389] br[389] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_390 bl[390] br[390] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_391 bl[391] br[391] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_392 bl[392] br[392] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_393 bl[393] br[393] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_394 bl[394] br[394] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_395 bl[395] br[395] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_396 bl[396] br[396] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_397 bl[397] br[397] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_398 bl[398] br[398] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_399 bl[399] br[399] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_400 bl[400] br[400] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_401 bl[401] br[401] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_402 bl[402] br[402] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_403 bl[403] br[403] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_404 bl[404] br[404] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_405 bl[405] br[405] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_406 bl[406] br[406] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_407 bl[407] br[407] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_408 bl[408] br[408] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_409 bl[409] br[409] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_410 bl[410] br[410] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_411 bl[411] br[411] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_412 bl[412] br[412] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_413 bl[413] br[413] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_414 bl[414] br[414] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_415 bl[415] br[415] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_416 bl[416] br[416] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_417 bl[417] br[417] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_418 bl[418] br[418] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_419 bl[419] br[419] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_420 bl[420] br[420] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_421 bl[421] br[421] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_422 bl[422] br[422] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_423 bl[423] br[423] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_424 bl[424] br[424] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_425 bl[425] br[425] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_426 bl[426] br[426] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_427 bl[427] br[427] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_428 bl[428] br[428] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_429 bl[429] br[429] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_430 bl[430] br[430] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_431 bl[431] br[431] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_432 bl[432] br[432] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_433 bl[433] br[433] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_434 bl[434] br[434] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_435 bl[435] br[435] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_436 bl[436] br[436] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_437 bl[437] br[437] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_438 bl[438] br[438] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_439 bl[439] br[439] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_440 bl[440] br[440] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_441 bl[441] br[441] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_442 bl[442] br[442] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_443 bl[443] br[443] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_444 bl[444] br[444] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_445 bl[445] br[445] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_446 bl[446] br[446] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_447 bl[447] br[447] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_448 bl[448] br[448] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_449 bl[449] br[449] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_450 bl[450] br[450] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_451 bl[451] br[451] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_452 bl[452] br[452] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_453 bl[453] br[453] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_454 bl[454] br[454] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_455 bl[455] br[455] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_456 bl[456] br[456] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_457 bl[457] br[457] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_458 bl[458] br[458] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_459 bl[459] br[459] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_460 bl[460] br[460] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_461 bl[461] br[461] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_462 bl[462] br[462] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_463 bl[463] br[463] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_464 bl[464] br[464] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_465 bl[465] br[465] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_466 bl[466] br[466] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_467 bl[467] br[467] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_468 bl[468] br[468] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_469 bl[469] br[469] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_470 bl[470] br[470] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_471 bl[471] br[471] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_472 bl[472] br[472] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_473 bl[473] br[473] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_474 bl[474] br[474] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_475 bl[475] br[475] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_476 bl[476] br[476] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_477 bl[477] br[477] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_478 bl[478] br[478] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_479 bl[479] br[479] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_480 bl[480] br[480] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_481 bl[481] br[481] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_482 bl[482] br[482] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_483 bl[483] br[483] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_484 bl[484] br[484] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_485 bl[485] br[485] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_486 bl[486] br[486] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_487 bl[487] br[487] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_488 bl[488] br[488] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_489 bl[489] br[489] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_490 bl[490] br[490] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_491 bl[491] br[491] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_492 bl[492] br[492] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_493 bl[493] br[493] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_494 bl[494] br[494] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_495 bl[495] br[495] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_496 bl[496] br[496] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_497 bl[497] br[497] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_498 bl[498] br[498] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_499 bl[499] br[499] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_500 bl[500] br[500] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_501 bl[501] br[501] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_502 bl[502] br[502] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_503 bl[503] br[503] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_504 bl[504] br[504] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_505 bl[505] br[505] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_506 bl[506] br[506] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_507 bl[507] br[507] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_508 bl[508] br[508] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_509 bl[509] br[509] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_510 bl[510] br[510] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_3_511 bl[511] br[511] vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xcell_4_0 bl[0] br[0] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_1 bl[1] br[1] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_2 bl[2] br[2] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_3 bl[3] br[3] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_4 bl[4] br[4] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_5 bl[5] br[5] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_6 bl[6] br[6] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_7 bl[7] br[7] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_8 bl[8] br[8] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_9 bl[9] br[9] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_10 bl[10] br[10] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_11 bl[11] br[11] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_12 bl[12] br[12] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_13 bl[13] br[13] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_14 bl[14] br[14] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_15 bl[15] br[15] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_16 bl[16] br[16] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_17 bl[17] br[17] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_18 bl[18] br[18] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_19 bl[19] br[19] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_20 bl[20] br[20] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_21 bl[21] br[21] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_22 bl[22] br[22] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_23 bl[23] br[23] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_24 bl[24] br[24] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_25 bl[25] br[25] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_26 bl[26] br[26] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_27 bl[27] br[27] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_28 bl[28] br[28] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_29 bl[29] br[29] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_30 bl[30] br[30] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_31 bl[31] br[31] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_32 bl[32] br[32] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_33 bl[33] br[33] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_34 bl[34] br[34] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_35 bl[35] br[35] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_36 bl[36] br[36] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_37 bl[37] br[37] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_38 bl[38] br[38] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_39 bl[39] br[39] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_40 bl[40] br[40] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_41 bl[41] br[41] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_42 bl[42] br[42] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_43 bl[43] br[43] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_44 bl[44] br[44] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_45 bl[45] br[45] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_46 bl[46] br[46] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_47 bl[47] br[47] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_48 bl[48] br[48] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_49 bl[49] br[49] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_50 bl[50] br[50] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_51 bl[51] br[51] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_52 bl[52] br[52] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_53 bl[53] br[53] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_54 bl[54] br[54] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_55 bl[55] br[55] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_56 bl[56] br[56] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_57 bl[57] br[57] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_58 bl[58] br[58] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_59 bl[59] br[59] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_60 bl[60] br[60] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_61 bl[61] br[61] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_62 bl[62] br[62] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_63 bl[63] br[63] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_64 bl[64] br[64] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_65 bl[65] br[65] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_66 bl[66] br[66] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_67 bl[67] br[67] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_68 bl[68] br[68] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_69 bl[69] br[69] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_70 bl[70] br[70] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_71 bl[71] br[71] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_72 bl[72] br[72] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_73 bl[73] br[73] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_74 bl[74] br[74] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_75 bl[75] br[75] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_76 bl[76] br[76] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_77 bl[77] br[77] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_78 bl[78] br[78] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_79 bl[79] br[79] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_80 bl[80] br[80] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_81 bl[81] br[81] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_82 bl[82] br[82] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_83 bl[83] br[83] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_84 bl[84] br[84] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_85 bl[85] br[85] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_86 bl[86] br[86] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_87 bl[87] br[87] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_88 bl[88] br[88] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_89 bl[89] br[89] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_90 bl[90] br[90] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_91 bl[91] br[91] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_92 bl[92] br[92] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_93 bl[93] br[93] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_94 bl[94] br[94] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_95 bl[95] br[95] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_96 bl[96] br[96] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_97 bl[97] br[97] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_98 bl[98] br[98] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_99 bl[99] br[99] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_100 bl[100] br[100] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_101 bl[101] br[101] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_102 bl[102] br[102] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_103 bl[103] br[103] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_104 bl[104] br[104] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_105 bl[105] br[105] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_106 bl[106] br[106] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_107 bl[107] br[107] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_108 bl[108] br[108] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_109 bl[109] br[109] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_110 bl[110] br[110] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_111 bl[111] br[111] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_112 bl[112] br[112] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_113 bl[113] br[113] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_114 bl[114] br[114] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_115 bl[115] br[115] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_116 bl[116] br[116] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_117 bl[117] br[117] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_118 bl[118] br[118] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_119 bl[119] br[119] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_120 bl[120] br[120] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_121 bl[121] br[121] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_122 bl[122] br[122] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_123 bl[123] br[123] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_124 bl[124] br[124] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_125 bl[125] br[125] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_126 bl[126] br[126] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_127 bl[127] br[127] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_128 bl[128] br[128] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_129 bl[129] br[129] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_130 bl[130] br[130] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_131 bl[131] br[131] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_132 bl[132] br[132] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_133 bl[133] br[133] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_134 bl[134] br[134] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_135 bl[135] br[135] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_136 bl[136] br[136] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_137 bl[137] br[137] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_138 bl[138] br[138] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_139 bl[139] br[139] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_140 bl[140] br[140] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_141 bl[141] br[141] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_142 bl[142] br[142] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_143 bl[143] br[143] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_144 bl[144] br[144] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_145 bl[145] br[145] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_146 bl[146] br[146] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_147 bl[147] br[147] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_148 bl[148] br[148] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_149 bl[149] br[149] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_150 bl[150] br[150] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_151 bl[151] br[151] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_152 bl[152] br[152] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_153 bl[153] br[153] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_154 bl[154] br[154] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_155 bl[155] br[155] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_156 bl[156] br[156] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_157 bl[157] br[157] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_158 bl[158] br[158] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_159 bl[159] br[159] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_160 bl[160] br[160] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_161 bl[161] br[161] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_162 bl[162] br[162] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_163 bl[163] br[163] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_164 bl[164] br[164] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_165 bl[165] br[165] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_166 bl[166] br[166] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_167 bl[167] br[167] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_168 bl[168] br[168] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_169 bl[169] br[169] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_170 bl[170] br[170] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_171 bl[171] br[171] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_172 bl[172] br[172] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_173 bl[173] br[173] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_174 bl[174] br[174] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_175 bl[175] br[175] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_176 bl[176] br[176] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_177 bl[177] br[177] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_178 bl[178] br[178] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_179 bl[179] br[179] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_180 bl[180] br[180] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_181 bl[181] br[181] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_182 bl[182] br[182] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_183 bl[183] br[183] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_184 bl[184] br[184] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_185 bl[185] br[185] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_186 bl[186] br[186] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_187 bl[187] br[187] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_188 bl[188] br[188] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_189 bl[189] br[189] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_190 bl[190] br[190] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_191 bl[191] br[191] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_192 bl[192] br[192] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_193 bl[193] br[193] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_194 bl[194] br[194] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_195 bl[195] br[195] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_196 bl[196] br[196] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_197 bl[197] br[197] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_198 bl[198] br[198] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_199 bl[199] br[199] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_200 bl[200] br[200] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_201 bl[201] br[201] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_202 bl[202] br[202] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_203 bl[203] br[203] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_204 bl[204] br[204] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_205 bl[205] br[205] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_206 bl[206] br[206] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_207 bl[207] br[207] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_208 bl[208] br[208] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_209 bl[209] br[209] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_210 bl[210] br[210] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_211 bl[211] br[211] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_212 bl[212] br[212] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_213 bl[213] br[213] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_214 bl[214] br[214] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_215 bl[215] br[215] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_216 bl[216] br[216] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_217 bl[217] br[217] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_218 bl[218] br[218] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_219 bl[219] br[219] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_220 bl[220] br[220] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_221 bl[221] br[221] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_222 bl[222] br[222] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_223 bl[223] br[223] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_224 bl[224] br[224] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_225 bl[225] br[225] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_226 bl[226] br[226] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_227 bl[227] br[227] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_228 bl[228] br[228] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_229 bl[229] br[229] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_230 bl[230] br[230] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_231 bl[231] br[231] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_232 bl[232] br[232] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_233 bl[233] br[233] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_234 bl[234] br[234] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_235 bl[235] br[235] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_236 bl[236] br[236] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_237 bl[237] br[237] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_238 bl[238] br[238] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_239 bl[239] br[239] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_240 bl[240] br[240] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_241 bl[241] br[241] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_242 bl[242] br[242] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_243 bl[243] br[243] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_244 bl[244] br[244] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_245 bl[245] br[245] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_246 bl[246] br[246] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_247 bl[247] br[247] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_248 bl[248] br[248] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_249 bl[249] br[249] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_250 bl[250] br[250] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_251 bl[251] br[251] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_252 bl[252] br[252] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_253 bl[253] br[253] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_254 bl[254] br[254] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_255 bl[255] br[255] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_256 bl[256] br[256] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_257 bl[257] br[257] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_258 bl[258] br[258] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_259 bl[259] br[259] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_260 bl[260] br[260] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_261 bl[261] br[261] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_262 bl[262] br[262] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_263 bl[263] br[263] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_264 bl[264] br[264] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_265 bl[265] br[265] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_266 bl[266] br[266] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_267 bl[267] br[267] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_268 bl[268] br[268] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_269 bl[269] br[269] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_270 bl[270] br[270] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_271 bl[271] br[271] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_272 bl[272] br[272] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_273 bl[273] br[273] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_274 bl[274] br[274] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_275 bl[275] br[275] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_276 bl[276] br[276] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_277 bl[277] br[277] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_278 bl[278] br[278] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_279 bl[279] br[279] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_280 bl[280] br[280] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_281 bl[281] br[281] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_282 bl[282] br[282] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_283 bl[283] br[283] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_284 bl[284] br[284] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_285 bl[285] br[285] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_286 bl[286] br[286] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_287 bl[287] br[287] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_288 bl[288] br[288] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_289 bl[289] br[289] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_290 bl[290] br[290] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_291 bl[291] br[291] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_292 bl[292] br[292] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_293 bl[293] br[293] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_294 bl[294] br[294] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_295 bl[295] br[295] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_296 bl[296] br[296] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_297 bl[297] br[297] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_298 bl[298] br[298] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_299 bl[299] br[299] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_300 bl[300] br[300] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_301 bl[301] br[301] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_302 bl[302] br[302] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_303 bl[303] br[303] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_304 bl[304] br[304] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_305 bl[305] br[305] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_306 bl[306] br[306] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_307 bl[307] br[307] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_308 bl[308] br[308] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_309 bl[309] br[309] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_310 bl[310] br[310] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_311 bl[311] br[311] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_312 bl[312] br[312] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_313 bl[313] br[313] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_314 bl[314] br[314] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_315 bl[315] br[315] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_316 bl[316] br[316] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_317 bl[317] br[317] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_318 bl[318] br[318] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_319 bl[319] br[319] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_320 bl[320] br[320] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_321 bl[321] br[321] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_322 bl[322] br[322] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_323 bl[323] br[323] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_324 bl[324] br[324] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_325 bl[325] br[325] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_326 bl[326] br[326] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_327 bl[327] br[327] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_328 bl[328] br[328] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_329 bl[329] br[329] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_330 bl[330] br[330] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_331 bl[331] br[331] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_332 bl[332] br[332] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_333 bl[333] br[333] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_334 bl[334] br[334] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_335 bl[335] br[335] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_336 bl[336] br[336] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_337 bl[337] br[337] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_338 bl[338] br[338] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_339 bl[339] br[339] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_340 bl[340] br[340] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_341 bl[341] br[341] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_342 bl[342] br[342] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_343 bl[343] br[343] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_344 bl[344] br[344] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_345 bl[345] br[345] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_346 bl[346] br[346] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_347 bl[347] br[347] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_348 bl[348] br[348] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_349 bl[349] br[349] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_350 bl[350] br[350] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_351 bl[351] br[351] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_352 bl[352] br[352] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_353 bl[353] br[353] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_354 bl[354] br[354] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_355 bl[355] br[355] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_356 bl[356] br[356] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_357 bl[357] br[357] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_358 bl[358] br[358] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_359 bl[359] br[359] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_360 bl[360] br[360] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_361 bl[361] br[361] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_362 bl[362] br[362] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_363 bl[363] br[363] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_364 bl[364] br[364] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_365 bl[365] br[365] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_366 bl[366] br[366] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_367 bl[367] br[367] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_368 bl[368] br[368] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_369 bl[369] br[369] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_370 bl[370] br[370] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_371 bl[371] br[371] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_372 bl[372] br[372] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_373 bl[373] br[373] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_374 bl[374] br[374] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_375 bl[375] br[375] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_376 bl[376] br[376] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_377 bl[377] br[377] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_378 bl[378] br[378] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_379 bl[379] br[379] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_380 bl[380] br[380] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_381 bl[381] br[381] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_382 bl[382] br[382] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_383 bl[383] br[383] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_384 bl[384] br[384] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_385 bl[385] br[385] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_386 bl[386] br[386] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_387 bl[387] br[387] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_388 bl[388] br[388] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_389 bl[389] br[389] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_390 bl[390] br[390] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_391 bl[391] br[391] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_392 bl[392] br[392] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_393 bl[393] br[393] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_394 bl[394] br[394] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_395 bl[395] br[395] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_396 bl[396] br[396] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_397 bl[397] br[397] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_398 bl[398] br[398] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_399 bl[399] br[399] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_400 bl[400] br[400] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_401 bl[401] br[401] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_402 bl[402] br[402] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_403 bl[403] br[403] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_404 bl[404] br[404] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_405 bl[405] br[405] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_406 bl[406] br[406] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_407 bl[407] br[407] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_408 bl[408] br[408] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_409 bl[409] br[409] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_410 bl[410] br[410] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_411 bl[411] br[411] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_412 bl[412] br[412] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_413 bl[413] br[413] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_414 bl[414] br[414] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_415 bl[415] br[415] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_416 bl[416] br[416] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_417 bl[417] br[417] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_418 bl[418] br[418] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_419 bl[419] br[419] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_420 bl[420] br[420] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_421 bl[421] br[421] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_422 bl[422] br[422] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_423 bl[423] br[423] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_424 bl[424] br[424] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_425 bl[425] br[425] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_426 bl[426] br[426] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_427 bl[427] br[427] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_428 bl[428] br[428] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_429 bl[429] br[429] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_430 bl[430] br[430] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_431 bl[431] br[431] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_432 bl[432] br[432] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_433 bl[433] br[433] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_434 bl[434] br[434] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_435 bl[435] br[435] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_436 bl[436] br[436] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_437 bl[437] br[437] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_438 bl[438] br[438] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_439 bl[439] br[439] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_440 bl[440] br[440] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_441 bl[441] br[441] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_442 bl[442] br[442] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_443 bl[443] br[443] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_444 bl[444] br[444] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_445 bl[445] br[445] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_446 bl[446] br[446] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_447 bl[447] br[447] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_448 bl[448] br[448] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_449 bl[449] br[449] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_450 bl[450] br[450] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_451 bl[451] br[451] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_452 bl[452] br[452] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_453 bl[453] br[453] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_454 bl[454] br[454] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_455 bl[455] br[455] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_456 bl[456] br[456] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_457 bl[457] br[457] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_458 bl[458] br[458] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_459 bl[459] br[459] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_460 bl[460] br[460] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_461 bl[461] br[461] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_462 bl[462] br[462] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_463 bl[463] br[463] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_464 bl[464] br[464] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_465 bl[465] br[465] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_466 bl[466] br[466] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_467 bl[467] br[467] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_468 bl[468] br[468] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_469 bl[469] br[469] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_470 bl[470] br[470] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_471 bl[471] br[471] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_472 bl[472] br[472] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_473 bl[473] br[473] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_474 bl[474] br[474] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_475 bl[475] br[475] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_476 bl[476] br[476] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_477 bl[477] br[477] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_478 bl[478] br[478] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_479 bl[479] br[479] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_480 bl[480] br[480] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_481 bl[481] br[481] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_482 bl[482] br[482] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_483 bl[483] br[483] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_484 bl[484] br[484] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_485 bl[485] br[485] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_486 bl[486] br[486] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_487 bl[487] br[487] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_488 bl[488] br[488] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_489 bl[489] br[489] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_490 bl[490] br[490] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_491 bl[491] br[491] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_492 bl[492] br[492] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_493 bl[493] br[493] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_494 bl[494] br[494] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_495 bl[495] br[495] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_496 bl[496] br[496] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_497 bl[497] br[497] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_498 bl[498] br[498] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_499 bl[499] br[499] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_500 bl[500] br[500] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_501 bl[501] br[501] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_502 bl[502] br[502] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_503 bl[503] br[503] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_504 bl[504] br[504] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_505 bl[505] br[505] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_506 bl[506] br[506] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_507 bl[507] br[507] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_508 bl[508] br[508] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_509 bl[509] br[509] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_510 bl[510] br[510] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_4_511 bl[511] br[511] vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xcell_5_0 bl[0] br[0] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_1 bl[1] br[1] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_2 bl[2] br[2] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_3 bl[3] br[3] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_4 bl[4] br[4] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_5 bl[5] br[5] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_6 bl[6] br[6] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_7 bl[7] br[7] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_8 bl[8] br[8] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_9 bl[9] br[9] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_10 bl[10] br[10] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_11 bl[11] br[11] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_12 bl[12] br[12] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_13 bl[13] br[13] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_14 bl[14] br[14] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_15 bl[15] br[15] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_16 bl[16] br[16] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_17 bl[17] br[17] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_18 bl[18] br[18] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_19 bl[19] br[19] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_20 bl[20] br[20] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_21 bl[21] br[21] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_22 bl[22] br[22] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_23 bl[23] br[23] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_24 bl[24] br[24] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_25 bl[25] br[25] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_26 bl[26] br[26] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_27 bl[27] br[27] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_28 bl[28] br[28] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_29 bl[29] br[29] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_30 bl[30] br[30] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_31 bl[31] br[31] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_32 bl[32] br[32] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_33 bl[33] br[33] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_34 bl[34] br[34] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_35 bl[35] br[35] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_36 bl[36] br[36] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_37 bl[37] br[37] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_38 bl[38] br[38] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_39 bl[39] br[39] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_40 bl[40] br[40] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_41 bl[41] br[41] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_42 bl[42] br[42] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_43 bl[43] br[43] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_44 bl[44] br[44] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_45 bl[45] br[45] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_46 bl[46] br[46] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_47 bl[47] br[47] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_48 bl[48] br[48] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_49 bl[49] br[49] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_50 bl[50] br[50] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_51 bl[51] br[51] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_52 bl[52] br[52] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_53 bl[53] br[53] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_54 bl[54] br[54] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_55 bl[55] br[55] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_56 bl[56] br[56] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_57 bl[57] br[57] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_58 bl[58] br[58] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_59 bl[59] br[59] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_60 bl[60] br[60] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_61 bl[61] br[61] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_62 bl[62] br[62] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_63 bl[63] br[63] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_64 bl[64] br[64] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_65 bl[65] br[65] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_66 bl[66] br[66] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_67 bl[67] br[67] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_68 bl[68] br[68] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_69 bl[69] br[69] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_70 bl[70] br[70] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_71 bl[71] br[71] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_72 bl[72] br[72] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_73 bl[73] br[73] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_74 bl[74] br[74] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_75 bl[75] br[75] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_76 bl[76] br[76] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_77 bl[77] br[77] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_78 bl[78] br[78] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_79 bl[79] br[79] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_80 bl[80] br[80] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_81 bl[81] br[81] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_82 bl[82] br[82] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_83 bl[83] br[83] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_84 bl[84] br[84] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_85 bl[85] br[85] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_86 bl[86] br[86] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_87 bl[87] br[87] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_88 bl[88] br[88] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_89 bl[89] br[89] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_90 bl[90] br[90] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_91 bl[91] br[91] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_92 bl[92] br[92] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_93 bl[93] br[93] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_94 bl[94] br[94] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_95 bl[95] br[95] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_96 bl[96] br[96] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_97 bl[97] br[97] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_98 bl[98] br[98] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_99 bl[99] br[99] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_100 bl[100] br[100] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_101 bl[101] br[101] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_102 bl[102] br[102] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_103 bl[103] br[103] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_104 bl[104] br[104] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_105 bl[105] br[105] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_106 bl[106] br[106] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_107 bl[107] br[107] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_108 bl[108] br[108] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_109 bl[109] br[109] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_110 bl[110] br[110] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_111 bl[111] br[111] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_112 bl[112] br[112] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_113 bl[113] br[113] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_114 bl[114] br[114] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_115 bl[115] br[115] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_116 bl[116] br[116] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_117 bl[117] br[117] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_118 bl[118] br[118] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_119 bl[119] br[119] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_120 bl[120] br[120] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_121 bl[121] br[121] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_122 bl[122] br[122] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_123 bl[123] br[123] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_124 bl[124] br[124] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_125 bl[125] br[125] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_126 bl[126] br[126] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_127 bl[127] br[127] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_128 bl[128] br[128] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_129 bl[129] br[129] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_130 bl[130] br[130] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_131 bl[131] br[131] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_132 bl[132] br[132] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_133 bl[133] br[133] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_134 bl[134] br[134] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_135 bl[135] br[135] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_136 bl[136] br[136] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_137 bl[137] br[137] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_138 bl[138] br[138] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_139 bl[139] br[139] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_140 bl[140] br[140] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_141 bl[141] br[141] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_142 bl[142] br[142] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_143 bl[143] br[143] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_144 bl[144] br[144] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_145 bl[145] br[145] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_146 bl[146] br[146] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_147 bl[147] br[147] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_148 bl[148] br[148] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_149 bl[149] br[149] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_150 bl[150] br[150] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_151 bl[151] br[151] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_152 bl[152] br[152] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_153 bl[153] br[153] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_154 bl[154] br[154] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_155 bl[155] br[155] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_156 bl[156] br[156] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_157 bl[157] br[157] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_158 bl[158] br[158] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_159 bl[159] br[159] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_160 bl[160] br[160] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_161 bl[161] br[161] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_162 bl[162] br[162] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_163 bl[163] br[163] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_164 bl[164] br[164] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_165 bl[165] br[165] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_166 bl[166] br[166] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_167 bl[167] br[167] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_168 bl[168] br[168] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_169 bl[169] br[169] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_170 bl[170] br[170] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_171 bl[171] br[171] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_172 bl[172] br[172] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_173 bl[173] br[173] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_174 bl[174] br[174] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_175 bl[175] br[175] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_176 bl[176] br[176] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_177 bl[177] br[177] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_178 bl[178] br[178] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_179 bl[179] br[179] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_180 bl[180] br[180] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_181 bl[181] br[181] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_182 bl[182] br[182] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_183 bl[183] br[183] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_184 bl[184] br[184] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_185 bl[185] br[185] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_186 bl[186] br[186] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_187 bl[187] br[187] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_188 bl[188] br[188] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_189 bl[189] br[189] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_190 bl[190] br[190] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_191 bl[191] br[191] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_192 bl[192] br[192] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_193 bl[193] br[193] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_194 bl[194] br[194] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_195 bl[195] br[195] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_196 bl[196] br[196] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_197 bl[197] br[197] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_198 bl[198] br[198] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_199 bl[199] br[199] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_200 bl[200] br[200] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_201 bl[201] br[201] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_202 bl[202] br[202] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_203 bl[203] br[203] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_204 bl[204] br[204] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_205 bl[205] br[205] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_206 bl[206] br[206] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_207 bl[207] br[207] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_208 bl[208] br[208] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_209 bl[209] br[209] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_210 bl[210] br[210] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_211 bl[211] br[211] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_212 bl[212] br[212] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_213 bl[213] br[213] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_214 bl[214] br[214] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_215 bl[215] br[215] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_216 bl[216] br[216] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_217 bl[217] br[217] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_218 bl[218] br[218] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_219 bl[219] br[219] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_220 bl[220] br[220] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_221 bl[221] br[221] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_222 bl[222] br[222] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_223 bl[223] br[223] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_224 bl[224] br[224] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_225 bl[225] br[225] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_226 bl[226] br[226] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_227 bl[227] br[227] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_228 bl[228] br[228] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_229 bl[229] br[229] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_230 bl[230] br[230] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_231 bl[231] br[231] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_232 bl[232] br[232] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_233 bl[233] br[233] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_234 bl[234] br[234] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_235 bl[235] br[235] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_236 bl[236] br[236] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_237 bl[237] br[237] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_238 bl[238] br[238] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_239 bl[239] br[239] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_240 bl[240] br[240] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_241 bl[241] br[241] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_242 bl[242] br[242] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_243 bl[243] br[243] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_244 bl[244] br[244] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_245 bl[245] br[245] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_246 bl[246] br[246] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_247 bl[247] br[247] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_248 bl[248] br[248] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_249 bl[249] br[249] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_250 bl[250] br[250] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_251 bl[251] br[251] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_252 bl[252] br[252] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_253 bl[253] br[253] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_254 bl[254] br[254] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_255 bl[255] br[255] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_256 bl[256] br[256] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_257 bl[257] br[257] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_258 bl[258] br[258] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_259 bl[259] br[259] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_260 bl[260] br[260] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_261 bl[261] br[261] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_262 bl[262] br[262] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_263 bl[263] br[263] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_264 bl[264] br[264] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_265 bl[265] br[265] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_266 bl[266] br[266] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_267 bl[267] br[267] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_268 bl[268] br[268] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_269 bl[269] br[269] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_270 bl[270] br[270] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_271 bl[271] br[271] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_272 bl[272] br[272] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_273 bl[273] br[273] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_274 bl[274] br[274] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_275 bl[275] br[275] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_276 bl[276] br[276] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_277 bl[277] br[277] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_278 bl[278] br[278] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_279 bl[279] br[279] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_280 bl[280] br[280] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_281 bl[281] br[281] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_282 bl[282] br[282] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_283 bl[283] br[283] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_284 bl[284] br[284] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_285 bl[285] br[285] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_286 bl[286] br[286] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_287 bl[287] br[287] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_288 bl[288] br[288] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_289 bl[289] br[289] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_290 bl[290] br[290] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_291 bl[291] br[291] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_292 bl[292] br[292] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_293 bl[293] br[293] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_294 bl[294] br[294] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_295 bl[295] br[295] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_296 bl[296] br[296] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_297 bl[297] br[297] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_298 bl[298] br[298] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_299 bl[299] br[299] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_300 bl[300] br[300] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_301 bl[301] br[301] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_302 bl[302] br[302] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_303 bl[303] br[303] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_304 bl[304] br[304] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_305 bl[305] br[305] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_306 bl[306] br[306] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_307 bl[307] br[307] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_308 bl[308] br[308] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_309 bl[309] br[309] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_310 bl[310] br[310] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_311 bl[311] br[311] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_312 bl[312] br[312] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_313 bl[313] br[313] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_314 bl[314] br[314] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_315 bl[315] br[315] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_316 bl[316] br[316] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_317 bl[317] br[317] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_318 bl[318] br[318] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_319 bl[319] br[319] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_320 bl[320] br[320] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_321 bl[321] br[321] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_322 bl[322] br[322] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_323 bl[323] br[323] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_324 bl[324] br[324] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_325 bl[325] br[325] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_326 bl[326] br[326] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_327 bl[327] br[327] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_328 bl[328] br[328] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_329 bl[329] br[329] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_330 bl[330] br[330] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_331 bl[331] br[331] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_332 bl[332] br[332] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_333 bl[333] br[333] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_334 bl[334] br[334] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_335 bl[335] br[335] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_336 bl[336] br[336] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_337 bl[337] br[337] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_338 bl[338] br[338] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_339 bl[339] br[339] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_340 bl[340] br[340] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_341 bl[341] br[341] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_342 bl[342] br[342] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_343 bl[343] br[343] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_344 bl[344] br[344] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_345 bl[345] br[345] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_346 bl[346] br[346] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_347 bl[347] br[347] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_348 bl[348] br[348] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_349 bl[349] br[349] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_350 bl[350] br[350] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_351 bl[351] br[351] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_352 bl[352] br[352] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_353 bl[353] br[353] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_354 bl[354] br[354] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_355 bl[355] br[355] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_356 bl[356] br[356] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_357 bl[357] br[357] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_358 bl[358] br[358] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_359 bl[359] br[359] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_360 bl[360] br[360] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_361 bl[361] br[361] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_362 bl[362] br[362] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_363 bl[363] br[363] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_364 bl[364] br[364] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_365 bl[365] br[365] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_366 bl[366] br[366] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_367 bl[367] br[367] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_368 bl[368] br[368] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_369 bl[369] br[369] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_370 bl[370] br[370] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_371 bl[371] br[371] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_372 bl[372] br[372] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_373 bl[373] br[373] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_374 bl[374] br[374] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_375 bl[375] br[375] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_376 bl[376] br[376] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_377 bl[377] br[377] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_378 bl[378] br[378] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_379 bl[379] br[379] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_380 bl[380] br[380] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_381 bl[381] br[381] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_382 bl[382] br[382] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_383 bl[383] br[383] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_384 bl[384] br[384] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_385 bl[385] br[385] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_386 bl[386] br[386] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_387 bl[387] br[387] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_388 bl[388] br[388] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_389 bl[389] br[389] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_390 bl[390] br[390] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_391 bl[391] br[391] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_392 bl[392] br[392] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_393 bl[393] br[393] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_394 bl[394] br[394] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_395 bl[395] br[395] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_396 bl[396] br[396] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_397 bl[397] br[397] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_398 bl[398] br[398] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_399 bl[399] br[399] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_400 bl[400] br[400] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_401 bl[401] br[401] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_402 bl[402] br[402] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_403 bl[403] br[403] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_404 bl[404] br[404] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_405 bl[405] br[405] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_406 bl[406] br[406] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_407 bl[407] br[407] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_408 bl[408] br[408] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_409 bl[409] br[409] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_410 bl[410] br[410] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_411 bl[411] br[411] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_412 bl[412] br[412] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_413 bl[413] br[413] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_414 bl[414] br[414] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_415 bl[415] br[415] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_416 bl[416] br[416] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_417 bl[417] br[417] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_418 bl[418] br[418] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_419 bl[419] br[419] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_420 bl[420] br[420] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_421 bl[421] br[421] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_422 bl[422] br[422] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_423 bl[423] br[423] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_424 bl[424] br[424] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_425 bl[425] br[425] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_426 bl[426] br[426] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_427 bl[427] br[427] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_428 bl[428] br[428] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_429 bl[429] br[429] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_430 bl[430] br[430] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_431 bl[431] br[431] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_432 bl[432] br[432] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_433 bl[433] br[433] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_434 bl[434] br[434] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_435 bl[435] br[435] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_436 bl[436] br[436] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_437 bl[437] br[437] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_438 bl[438] br[438] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_439 bl[439] br[439] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_440 bl[440] br[440] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_441 bl[441] br[441] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_442 bl[442] br[442] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_443 bl[443] br[443] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_444 bl[444] br[444] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_445 bl[445] br[445] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_446 bl[446] br[446] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_447 bl[447] br[447] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_448 bl[448] br[448] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_449 bl[449] br[449] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_450 bl[450] br[450] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_451 bl[451] br[451] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_452 bl[452] br[452] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_453 bl[453] br[453] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_454 bl[454] br[454] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_455 bl[455] br[455] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_456 bl[456] br[456] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_457 bl[457] br[457] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_458 bl[458] br[458] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_459 bl[459] br[459] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_460 bl[460] br[460] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_461 bl[461] br[461] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_462 bl[462] br[462] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_463 bl[463] br[463] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_464 bl[464] br[464] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_465 bl[465] br[465] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_466 bl[466] br[466] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_467 bl[467] br[467] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_468 bl[468] br[468] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_469 bl[469] br[469] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_470 bl[470] br[470] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_471 bl[471] br[471] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_472 bl[472] br[472] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_473 bl[473] br[473] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_474 bl[474] br[474] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_475 bl[475] br[475] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_476 bl[476] br[476] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_477 bl[477] br[477] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_478 bl[478] br[478] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_479 bl[479] br[479] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_480 bl[480] br[480] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_481 bl[481] br[481] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_482 bl[482] br[482] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_483 bl[483] br[483] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_484 bl[484] br[484] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_485 bl[485] br[485] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_486 bl[486] br[486] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_487 bl[487] br[487] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_488 bl[488] br[488] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_489 bl[489] br[489] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_490 bl[490] br[490] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_491 bl[491] br[491] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_492 bl[492] br[492] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_493 bl[493] br[493] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_494 bl[494] br[494] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_495 bl[495] br[495] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_496 bl[496] br[496] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_497 bl[497] br[497] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_498 bl[498] br[498] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_499 bl[499] br[499] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_500 bl[500] br[500] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_501 bl[501] br[501] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_502 bl[502] br[502] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_503 bl[503] br[503] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_504 bl[504] br[504] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_505 bl[505] br[505] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_506 bl[506] br[506] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_507 bl[507] br[507] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_508 bl[508] br[508] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_509 bl[509] br[509] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_510 bl[510] br[510] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_5_511 bl[511] br[511] vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xcell_6_0 bl[0] br[0] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_1 bl[1] br[1] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_2 bl[2] br[2] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_3 bl[3] br[3] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_4 bl[4] br[4] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_5 bl[5] br[5] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_6 bl[6] br[6] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_7 bl[7] br[7] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_8 bl[8] br[8] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_9 bl[9] br[9] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_10 bl[10] br[10] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_11 bl[11] br[11] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_12 bl[12] br[12] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_13 bl[13] br[13] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_14 bl[14] br[14] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_15 bl[15] br[15] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_16 bl[16] br[16] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_17 bl[17] br[17] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_18 bl[18] br[18] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_19 bl[19] br[19] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_20 bl[20] br[20] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_21 bl[21] br[21] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_22 bl[22] br[22] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_23 bl[23] br[23] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_24 bl[24] br[24] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_25 bl[25] br[25] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_26 bl[26] br[26] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_27 bl[27] br[27] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_28 bl[28] br[28] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_29 bl[29] br[29] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_30 bl[30] br[30] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_31 bl[31] br[31] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_32 bl[32] br[32] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_33 bl[33] br[33] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_34 bl[34] br[34] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_35 bl[35] br[35] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_36 bl[36] br[36] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_37 bl[37] br[37] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_38 bl[38] br[38] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_39 bl[39] br[39] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_40 bl[40] br[40] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_41 bl[41] br[41] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_42 bl[42] br[42] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_43 bl[43] br[43] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_44 bl[44] br[44] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_45 bl[45] br[45] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_46 bl[46] br[46] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_47 bl[47] br[47] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_48 bl[48] br[48] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_49 bl[49] br[49] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_50 bl[50] br[50] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_51 bl[51] br[51] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_52 bl[52] br[52] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_53 bl[53] br[53] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_54 bl[54] br[54] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_55 bl[55] br[55] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_56 bl[56] br[56] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_57 bl[57] br[57] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_58 bl[58] br[58] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_59 bl[59] br[59] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_60 bl[60] br[60] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_61 bl[61] br[61] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_62 bl[62] br[62] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_63 bl[63] br[63] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_64 bl[64] br[64] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_65 bl[65] br[65] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_66 bl[66] br[66] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_67 bl[67] br[67] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_68 bl[68] br[68] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_69 bl[69] br[69] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_70 bl[70] br[70] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_71 bl[71] br[71] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_72 bl[72] br[72] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_73 bl[73] br[73] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_74 bl[74] br[74] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_75 bl[75] br[75] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_76 bl[76] br[76] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_77 bl[77] br[77] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_78 bl[78] br[78] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_79 bl[79] br[79] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_80 bl[80] br[80] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_81 bl[81] br[81] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_82 bl[82] br[82] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_83 bl[83] br[83] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_84 bl[84] br[84] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_85 bl[85] br[85] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_86 bl[86] br[86] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_87 bl[87] br[87] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_88 bl[88] br[88] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_89 bl[89] br[89] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_90 bl[90] br[90] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_91 bl[91] br[91] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_92 bl[92] br[92] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_93 bl[93] br[93] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_94 bl[94] br[94] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_95 bl[95] br[95] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_96 bl[96] br[96] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_97 bl[97] br[97] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_98 bl[98] br[98] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_99 bl[99] br[99] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_100 bl[100] br[100] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_101 bl[101] br[101] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_102 bl[102] br[102] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_103 bl[103] br[103] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_104 bl[104] br[104] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_105 bl[105] br[105] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_106 bl[106] br[106] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_107 bl[107] br[107] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_108 bl[108] br[108] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_109 bl[109] br[109] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_110 bl[110] br[110] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_111 bl[111] br[111] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_112 bl[112] br[112] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_113 bl[113] br[113] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_114 bl[114] br[114] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_115 bl[115] br[115] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_116 bl[116] br[116] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_117 bl[117] br[117] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_118 bl[118] br[118] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_119 bl[119] br[119] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_120 bl[120] br[120] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_121 bl[121] br[121] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_122 bl[122] br[122] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_123 bl[123] br[123] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_124 bl[124] br[124] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_125 bl[125] br[125] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_126 bl[126] br[126] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_127 bl[127] br[127] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_128 bl[128] br[128] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_129 bl[129] br[129] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_130 bl[130] br[130] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_131 bl[131] br[131] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_132 bl[132] br[132] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_133 bl[133] br[133] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_134 bl[134] br[134] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_135 bl[135] br[135] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_136 bl[136] br[136] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_137 bl[137] br[137] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_138 bl[138] br[138] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_139 bl[139] br[139] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_140 bl[140] br[140] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_141 bl[141] br[141] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_142 bl[142] br[142] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_143 bl[143] br[143] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_144 bl[144] br[144] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_145 bl[145] br[145] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_146 bl[146] br[146] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_147 bl[147] br[147] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_148 bl[148] br[148] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_149 bl[149] br[149] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_150 bl[150] br[150] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_151 bl[151] br[151] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_152 bl[152] br[152] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_153 bl[153] br[153] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_154 bl[154] br[154] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_155 bl[155] br[155] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_156 bl[156] br[156] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_157 bl[157] br[157] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_158 bl[158] br[158] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_159 bl[159] br[159] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_160 bl[160] br[160] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_161 bl[161] br[161] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_162 bl[162] br[162] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_163 bl[163] br[163] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_164 bl[164] br[164] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_165 bl[165] br[165] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_166 bl[166] br[166] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_167 bl[167] br[167] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_168 bl[168] br[168] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_169 bl[169] br[169] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_170 bl[170] br[170] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_171 bl[171] br[171] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_172 bl[172] br[172] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_173 bl[173] br[173] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_174 bl[174] br[174] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_175 bl[175] br[175] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_176 bl[176] br[176] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_177 bl[177] br[177] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_178 bl[178] br[178] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_179 bl[179] br[179] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_180 bl[180] br[180] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_181 bl[181] br[181] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_182 bl[182] br[182] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_183 bl[183] br[183] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_184 bl[184] br[184] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_185 bl[185] br[185] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_186 bl[186] br[186] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_187 bl[187] br[187] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_188 bl[188] br[188] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_189 bl[189] br[189] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_190 bl[190] br[190] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_191 bl[191] br[191] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_192 bl[192] br[192] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_193 bl[193] br[193] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_194 bl[194] br[194] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_195 bl[195] br[195] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_196 bl[196] br[196] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_197 bl[197] br[197] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_198 bl[198] br[198] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_199 bl[199] br[199] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_200 bl[200] br[200] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_201 bl[201] br[201] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_202 bl[202] br[202] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_203 bl[203] br[203] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_204 bl[204] br[204] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_205 bl[205] br[205] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_206 bl[206] br[206] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_207 bl[207] br[207] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_208 bl[208] br[208] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_209 bl[209] br[209] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_210 bl[210] br[210] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_211 bl[211] br[211] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_212 bl[212] br[212] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_213 bl[213] br[213] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_214 bl[214] br[214] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_215 bl[215] br[215] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_216 bl[216] br[216] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_217 bl[217] br[217] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_218 bl[218] br[218] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_219 bl[219] br[219] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_220 bl[220] br[220] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_221 bl[221] br[221] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_222 bl[222] br[222] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_223 bl[223] br[223] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_224 bl[224] br[224] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_225 bl[225] br[225] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_226 bl[226] br[226] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_227 bl[227] br[227] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_228 bl[228] br[228] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_229 bl[229] br[229] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_230 bl[230] br[230] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_231 bl[231] br[231] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_232 bl[232] br[232] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_233 bl[233] br[233] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_234 bl[234] br[234] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_235 bl[235] br[235] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_236 bl[236] br[236] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_237 bl[237] br[237] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_238 bl[238] br[238] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_239 bl[239] br[239] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_240 bl[240] br[240] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_241 bl[241] br[241] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_242 bl[242] br[242] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_243 bl[243] br[243] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_244 bl[244] br[244] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_245 bl[245] br[245] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_246 bl[246] br[246] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_247 bl[247] br[247] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_248 bl[248] br[248] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_249 bl[249] br[249] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_250 bl[250] br[250] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_251 bl[251] br[251] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_252 bl[252] br[252] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_253 bl[253] br[253] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_254 bl[254] br[254] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_255 bl[255] br[255] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_256 bl[256] br[256] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_257 bl[257] br[257] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_258 bl[258] br[258] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_259 bl[259] br[259] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_260 bl[260] br[260] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_261 bl[261] br[261] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_262 bl[262] br[262] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_263 bl[263] br[263] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_264 bl[264] br[264] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_265 bl[265] br[265] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_266 bl[266] br[266] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_267 bl[267] br[267] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_268 bl[268] br[268] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_269 bl[269] br[269] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_270 bl[270] br[270] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_271 bl[271] br[271] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_272 bl[272] br[272] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_273 bl[273] br[273] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_274 bl[274] br[274] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_275 bl[275] br[275] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_276 bl[276] br[276] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_277 bl[277] br[277] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_278 bl[278] br[278] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_279 bl[279] br[279] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_280 bl[280] br[280] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_281 bl[281] br[281] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_282 bl[282] br[282] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_283 bl[283] br[283] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_284 bl[284] br[284] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_285 bl[285] br[285] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_286 bl[286] br[286] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_287 bl[287] br[287] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_288 bl[288] br[288] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_289 bl[289] br[289] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_290 bl[290] br[290] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_291 bl[291] br[291] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_292 bl[292] br[292] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_293 bl[293] br[293] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_294 bl[294] br[294] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_295 bl[295] br[295] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_296 bl[296] br[296] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_297 bl[297] br[297] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_298 bl[298] br[298] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_299 bl[299] br[299] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_300 bl[300] br[300] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_301 bl[301] br[301] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_302 bl[302] br[302] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_303 bl[303] br[303] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_304 bl[304] br[304] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_305 bl[305] br[305] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_306 bl[306] br[306] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_307 bl[307] br[307] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_308 bl[308] br[308] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_309 bl[309] br[309] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_310 bl[310] br[310] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_311 bl[311] br[311] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_312 bl[312] br[312] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_313 bl[313] br[313] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_314 bl[314] br[314] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_315 bl[315] br[315] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_316 bl[316] br[316] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_317 bl[317] br[317] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_318 bl[318] br[318] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_319 bl[319] br[319] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_320 bl[320] br[320] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_321 bl[321] br[321] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_322 bl[322] br[322] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_323 bl[323] br[323] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_324 bl[324] br[324] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_325 bl[325] br[325] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_326 bl[326] br[326] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_327 bl[327] br[327] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_328 bl[328] br[328] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_329 bl[329] br[329] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_330 bl[330] br[330] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_331 bl[331] br[331] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_332 bl[332] br[332] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_333 bl[333] br[333] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_334 bl[334] br[334] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_335 bl[335] br[335] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_336 bl[336] br[336] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_337 bl[337] br[337] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_338 bl[338] br[338] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_339 bl[339] br[339] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_340 bl[340] br[340] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_341 bl[341] br[341] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_342 bl[342] br[342] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_343 bl[343] br[343] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_344 bl[344] br[344] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_345 bl[345] br[345] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_346 bl[346] br[346] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_347 bl[347] br[347] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_348 bl[348] br[348] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_349 bl[349] br[349] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_350 bl[350] br[350] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_351 bl[351] br[351] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_352 bl[352] br[352] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_353 bl[353] br[353] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_354 bl[354] br[354] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_355 bl[355] br[355] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_356 bl[356] br[356] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_357 bl[357] br[357] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_358 bl[358] br[358] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_359 bl[359] br[359] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_360 bl[360] br[360] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_361 bl[361] br[361] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_362 bl[362] br[362] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_363 bl[363] br[363] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_364 bl[364] br[364] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_365 bl[365] br[365] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_366 bl[366] br[366] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_367 bl[367] br[367] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_368 bl[368] br[368] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_369 bl[369] br[369] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_370 bl[370] br[370] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_371 bl[371] br[371] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_372 bl[372] br[372] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_373 bl[373] br[373] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_374 bl[374] br[374] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_375 bl[375] br[375] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_376 bl[376] br[376] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_377 bl[377] br[377] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_378 bl[378] br[378] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_379 bl[379] br[379] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_380 bl[380] br[380] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_381 bl[381] br[381] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_382 bl[382] br[382] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_383 bl[383] br[383] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_384 bl[384] br[384] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_385 bl[385] br[385] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_386 bl[386] br[386] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_387 bl[387] br[387] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_388 bl[388] br[388] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_389 bl[389] br[389] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_390 bl[390] br[390] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_391 bl[391] br[391] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_392 bl[392] br[392] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_393 bl[393] br[393] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_394 bl[394] br[394] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_395 bl[395] br[395] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_396 bl[396] br[396] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_397 bl[397] br[397] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_398 bl[398] br[398] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_399 bl[399] br[399] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_400 bl[400] br[400] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_401 bl[401] br[401] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_402 bl[402] br[402] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_403 bl[403] br[403] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_404 bl[404] br[404] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_405 bl[405] br[405] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_406 bl[406] br[406] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_407 bl[407] br[407] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_408 bl[408] br[408] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_409 bl[409] br[409] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_410 bl[410] br[410] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_411 bl[411] br[411] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_412 bl[412] br[412] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_413 bl[413] br[413] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_414 bl[414] br[414] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_415 bl[415] br[415] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_416 bl[416] br[416] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_417 bl[417] br[417] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_418 bl[418] br[418] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_419 bl[419] br[419] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_420 bl[420] br[420] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_421 bl[421] br[421] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_422 bl[422] br[422] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_423 bl[423] br[423] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_424 bl[424] br[424] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_425 bl[425] br[425] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_426 bl[426] br[426] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_427 bl[427] br[427] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_428 bl[428] br[428] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_429 bl[429] br[429] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_430 bl[430] br[430] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_431 bl[431] br[431] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_432 bl[432] br[432] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_433 bl[433] br[433] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_434 bl[434] br[434] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_435 bl[435] br[435] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_436 bl[436] br[436] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_437 bl[437] br[437] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_438 bl[438] br[438] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_439 bl[439] br[439] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_440 bl[440] br[440] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_441 bl[441] br[441] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_442 bl[442] br[442] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_443 bl[443] br[443] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_444 bl[444] br[444] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_445 bl[445] br[445] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_446 bl[446] br[446] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_447 bl[447] br[447] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_448 bl[448] br[448] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_449 bl[449] br[449] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_450 bl[450] br[450] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_451 bl[451] br[451] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_452 bl[452] br[452] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_453 bl[453] br[453] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_454 bl[454] br[454] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_455 bl[455] br[455] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_456 bl[456] br[456] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_457 bl[457] br[457] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_458 bl[458] br[458] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_459 bl[459] br[459] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_460 bl[460] br[460] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_461 bl[461] br[461] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_462 bl[462] br[462] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_463 bl[463] br[463] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_464 bl[464] br[464] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_465 bl[465] br[465] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_466 bl[466] br[466] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_467 bl[467] br[467] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_468 bl[468] br[468] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_469 bl[469] br[469] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_470 bl[470] br[470] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_471 bl[471] br[471] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_472 bl[472] br[472] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_473 bl[473] br[473] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_474 bl[474] br[474] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_475 bl[475] br[475] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_476 bl[476] br[476] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_477 bl[477] br[477] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_478 bl[478] br[478] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_479 bl[479] br[479] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_480 bl[480] br[480] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_481 bl[481] br[481] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_482 bl[482] br[482] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_483 bl[483] br[483] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_484 bl[484] br[484] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_485 bl[485] br[485] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_486 bl[486] br[486] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_487 bl[487] br[487] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_488 bl[488] br[488] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_489 bl[489] br[489] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_490 bl[490] br[490] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_491 bl[491] br[491] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_492 bl[492] br[492] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_493 bl[493] br[493] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_494 bl[494] br[494] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_495 bl[495] br[495] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_496 bl[496] br[496] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_497 bl[497] br[497] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_498 bl[498] br[498] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_499 bl[499] br[499] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_500 bl[500] br[500] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_501 bl[501] br[501] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_502 bl[502] br[502] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_503 bl[503] br[503] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_504 bl[504] br[504] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_505 bl[505] br[505] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_506 bl[506] br[506] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_507 bl[507] br[507] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_508 bl[508] br[508] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_509 bl[509] br[509] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_510 bl[510] br[510] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_6_511 bl[511] br[511] vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xcell_7_0 bl[0] br[0] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_1 bl[1] br[1] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_2 bl[2] br[2] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_3 bl[3] br[3] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_4 bl[4] br[4] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_5 bl[5] br[5] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_6 bl[6] br[6] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_7 bl[7] br[7] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_8 bl[8] br[8] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_9 bl[9] br[9] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_10 bl[10] br[10] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_11 bl[11] br[11] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_12 bl[12] br[12] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_13 bl[13] br[13] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_14 bl[14] br[14] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_15 bl[15] br[15] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_16 bl[16] br[16] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_17 bl[17] br[17] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_18 bl[18] br[18] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_19 bl[19] br[19] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_20 bl[20] br[20] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_21 bl[21] br[21] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_22 bl[22] br[22] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_23 bl[23] br[23] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_24 bl[24] br[24] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_25 bl[25] br[25] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_26 bl[26] br[26] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_27 bl[27] br[27] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_28 bl[28] br[28] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_29 bl[29] br[29] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_30 bl[30] br[30] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_31 bl[31] br[31] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_32 bl[32] br[32] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_33 bl[33] br[33] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_34 bl[34] br[34] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_35 bl[35] br[35] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_36 bl[36] br[36] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_37 bl[37] br[37] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_38 bl[38] br[38] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_39 bl[39] br[39] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_40 bl[40] br[40] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_41 bl[41] br[41] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_42 bl[42] br[42] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_43 bl[43] br[43] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_44 bl[44] br[44] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_45 bl[45] br[45] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_46 bl[46] br[46] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_47 bl[47] br[47] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_48 bl[48] br[48] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_49 bl[49] br[49] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_50 bl[50] br[50] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_51 bl[51] br[51] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_52 bl[52] br[52] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_53 bl[53] br[53] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_54 bl[54] br[54] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_55 bl[55] br[55] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_56 bl[56] br[56] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_57 bl[57] br[57] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_58 bl[58] br[58] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_59 bl[59] br[59] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_60 bl[60] br[60] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_61 bl[61] br[61] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_62 bl[62] br[62] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_63 bl[63] br[63] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_64 bl[64] br[64] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_65 bl[65] br[65] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_66 bl[66] br[66] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_67 bl[67] br[67] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_68 bl[68] br[68] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_69 bl[69] br[69] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_70 bl[70] br[70] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_71 bl[71] br[71] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_72 bl[72] br[72] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_73 bl[73] br[73] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_74 bl[74] br[74] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_75 bl[75] br[75] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_76 bl[76] br[76] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_77 bl[77] br[77] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_78 bl[78] br[78] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_79 bl[79] br[79] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_80 bl[80] br[80] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_81 bl[81] br[81] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_82 bl[82] br[82] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_83 bl[83] br[83] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_84 bl[84] br[84] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_85 bl[85] br[85] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_86 bl[86] br[86] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_87 bl[87] br[87] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_88 bl[88] br[88] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_89 bl[89] br[89] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_90 bl[90] br[90] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_91 bl[91] br[91] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_92 bl[92] br[92] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_93 bl[93] br[93] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_94 bl[94] br[94] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_95 bl[95] br[95] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_96 bl[96] br[96] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_97 bl[97] br[97] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_98 bl[98] br[98] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_99 bl[99] br[99] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_100 bl[100] br[100] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_101 bl[101] br[101] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_102 bl[102] br[102] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_103 bl[103] br[103] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_104 bl[104] br[104] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_105 bl[105] br[105] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_106 bl[106] br[106] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_107 bl[107] br[107] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_108 bl[108] br[108] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_109 bl[109] br[109] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_110 bl[110] br[110] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_111 bl[111] br[111] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_112 bl[112] br[112] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_113 bl[113] br[113] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_114 bl[114] br[114] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_115 bl[115] br[115] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_116 bl[116] br[116] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_117 bl[117] br[117] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_118 bl[118] br[118] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_119 bl[119] br[119] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_120 bl[120] br[120] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_121 bl[121] br[121] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_122 bl[122] br[122] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_123 bl[123] br[123] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_124 bl[124] br[124] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_125 bl[125] br[125] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_126 bl[126] br[126] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_127 bl[127] br[127] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_128 bl[128] br[128] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_129 bl[129] br[129] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_130 bl[130] br[130] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_131 bl[131] br[131] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_132 bl[132] br[132] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_133 bl[133] br[133] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_134 bl[134] br[134] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_135 bl[135] br[135] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_136 bl[136] br[136] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_137 bl[137] br[137] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_138 bl[138] br[138] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_139 bl[139] br[139] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_140 bl[140] br[140] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_141 bl[141] br[141] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_142 bl[142] br[142] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_143 bl[143] br[143] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_144 bl[144] br[144] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_145 bl[145] br[145] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_146 bl[146] br[146] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_147 bl[147] br[147] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_148 bl[148] br[148] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_149 bl[149] br[149] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_150 bl[150] br[150] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_151 bl[151] br[151] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_152 bl[152] br[152] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_153 bl[153] br[153] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_154 bl[154] br[154] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_155 bl[155] br[155] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_156 bl[156] br[156] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_157 bl[157] br[157] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_158 bl[158] br[158] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_159 bl[159] br[159] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_160 bl[160] br[160] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_161 bl[161] br[161] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_162 bl[162] br[162] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_163 bl[163] br[163] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_164 bl[164] br[164] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_165 bl[165] br[165] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_166 bl[166] br[166] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_167 bl[167] br[167] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_168 bl[168] br[168] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_169 bl[169] br[169] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_170 bl[170] br[170] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_171 bl[171] br[171] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_172 bl[172] br[172] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_173 bl[173] br[173] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_174 bl[174] br[174] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_175 bl[175] br[175] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_176 bl[176] br[176] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_177 bl[177] br[177] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_178 bl[178] br[178] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_179 bl[179] br[179] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_180 bl[180] br[180] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_181 bl[181] br[181] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_182 bl[182] br[182] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_183 bl[183] br[183] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_184 bl[184] br[184] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_185 bl[185] br[185] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_186 bl[186] br[186] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_187 bl[187] br[187] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_188 bl[188] br[188] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_189 bl[189] br[189] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_190 bl[190] br[190] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_191 bl[191] br[191] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_192 bl[192] br[192] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_193 bl[193] br[193] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_194 bl[194] br[194] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_195 bl[195] br[195] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_196 bl[196] br[196] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_197 bl[197] br[197] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_198 bl[198] br[198] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_199 bl[199] br[199] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_200 bl[200] br[200] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_201 bl[201] br[201] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_202 bl[202] br[202] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_203 bl[203] br[203] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_204 bl[204] br[204] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_205 bl[205] br[205] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_206 bl[206] br[206] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_207 bl[207] br[207] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_208 bl[208] br[208] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_209 bl[209] br[209] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_210 bl[210] br[210] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_211 bl[211] br[211] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_212 bl[212] br[212] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_213 bl[213] br[213] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_214 bl[214] br[214] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_215 bl[215] br[215] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_216 bl[216] br[216] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_217 bl[217] br[217] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_218 bl[218] br[218] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_219 bl[219] br[219] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_220 bl[220] br[220] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_221 bl[221] br[221] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_222 bl[222] br[222] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_223 bl[223] br[223] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_224 bl[224] br[224] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_225 bl[225] br[225] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_226 bl[226] br[226] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_227 bl[227] br[227] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_228 bl[228] br[228] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_229 bl[229] br[229] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_230 bl[230] br[230] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_231 bl[231] br[231] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_232 bl[232] br[232] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_233 bl[233] br[233] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_234 bl[234] br[234] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_235 bl[235] br[235] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_236 bl[236] br[236] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_237 bl[237] br[237] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_238 bl[238] br[238] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_239 bl[239] br[239] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_240 bl[240] br[240] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_241 bl[241] br[241] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_242 bl[242] br[242] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_243 bl[243] br[243] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_244 bl[244] br[244] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_245 bl[245] br[245] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_246 bl[246] br[246] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_247 bl[247] br[247] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_248 bl[248] br[248] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_249 bl[249] br[249] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_250 bl[250] br[250] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_251 bl[251] br[251] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_252 bl[252] br[252] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_253 bl[253] br[253] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_254 bl[254] br[254] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_255 bl[255] br[255] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_256 bl[256] br[256] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_257 bl[257] br[257] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_258 bl[258] br[258] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_259 bl[259] br[259] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_260 bl[260] br[260] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_261 bl[261] br[261] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_262 bl[262] br[262] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_263 bl[263] br[263] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_264 bl[264] br[264] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_265 bl[265] br[265] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_266 bl[266] br[266] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_267 bl[267] br[267] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_268 bl[268] br[268] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_269 bl[269] br[269] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_270 bl[270] br[270] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_271 bl[271] br[271] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_272 bl[272] br[272] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_273 bl[273] br[273] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_274 bl[274] br[274] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_275 bl[275] br[275] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_276 bl[276] br[276] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_277 bl[277] br[277] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_278 bl[278] br[278] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_279 bl[279] br[279] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_280 bl[280] br[280] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_281 bl[281] br[281] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_282 bl[282] br[282] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_283 bl[283] br[283] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_284 bl[284] br[284] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_285 bl[285] br[285] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_286 bl[286] br[286] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_287 bl[287] br[287] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_288 bl[288] br[288] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_289 bl[289] br[289] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_290 bl[290] br[290] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_291 bl[291] br[291] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_292 bl[292] br[292] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_293 bl[293] br[293] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_294 bl[294] br[294] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_295 bl[295] br[295] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_296 bl[296] br[296] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_297 bl[297] br[297] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_298 bl[298] br[298] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_299 bl[299] br[299] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_300 bl[300] br[300] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_301 bl[301] br[301] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_302 bl[302] br[302] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_303 bl[303] br[303] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_304 bl[304] br[304] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_305 bl[305] br[305] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_306 bl[306] br[306] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_307 bl[307] br[307] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_308 bl[308] br[308] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_309 bl[309] br[309] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_310 bl[310] br[310] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_311 bl[311] br[311] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_312 bl[312] br[312] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_313 bl[313] br[313] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_314 bl[314] br[314] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_315 bl[315] br[315] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_316 bl[316] br[316] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_317 bl[317] br[317] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_318 bl[318] br[318] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_319 bl[319] br[319] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_320 bl[320] br[320] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_321 bl[321] br[321] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_322 bl[322] br[322] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_323 bl[323] br[323] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_324 bl[324] br[324] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_325 bl[325] br[325] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_326 bl[326] br[326] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_327 bl[327] br[327] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_328 bl[328] br[328] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_329 bl[329] br[329] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_330 bl[330] br[330] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_331 bl[331] br[331] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_332 bl[332] br[332] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_333 bl[333] br[333] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_334 bl[334] br[334] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_335 bl[335] br[335] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_336 bl[336] br[336] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_337 bl[337] br[337] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_338 bl[338] br[338] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_339 bl[339] br[339] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_340 bl[340] br[340] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_341 bl[341] br[341] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_342 bl[342] br[342] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_343 bl[343] br[343] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_344 bl[344] br[344] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_345 bl[345] br[345] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_346 bl[346] br[346] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_347 bl[347] br[347] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_348 bl[348] br[348] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_349 bl[349] br[349] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_350 bl[350] br[350] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_351 bl[351] br[351] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_352 bl[352] br[352] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_353 bl[353] br[353] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_354 bl[354] br[354] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_355 bl[355] br[355] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_356 bl[356] br[356] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_357 bl[357] br[357] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_358 bl[358] br[358] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_359 bl[359] br[359] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_360 bl[360] br[360] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_361 bl[361] br[361] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_362 bl[362] br[362] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_363 bl[363] br[363] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_364 bl[364] br[364] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_365 bl[365] br[365] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_366 bl[366] br[366] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_367 bl[367] br[367] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_368 bl[368] br[368] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_369 bl[369] br[369] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_370 bl[370] br[370] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_371 bl[371] br[371] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_372 bl[372] br[372] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_373 bl[373] br[373] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_374 bl[374] br[374] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_375 bl[375] br[375] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_376 bl[376] br[376] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_377 bl[377] br[377] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_378 bl[378] br[378] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_379 bl[379] br[379] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_380 bl[380] br[380] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_381 bl[381] br[381] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_382 bl[382] br[382] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_383 bl[383] br[383] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_384 bl[384] br[384] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_385 bl[385] br[385] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_386 bl[386] br[386] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_387 bl[387] br[387] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_388 bl[388] br[388] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_389 bl[389] br[389] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_390 bl[390] br[390] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_391 bl[391] br[391] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_392 bl[392] br[392] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_393 bl[393] br[393] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_394 bl[394] br[394] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_395 bl[395] br[395] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_396 bl[396] br[396] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_397 bl[397] br[397] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_398 bl[398] br[398] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_399 bl[399] br[399] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_400 bl[400] br[400] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_401 bl[401] br[401] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_402 bl[402] br[402] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_403 bl[403] br[403] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_404 bl[404] br[404] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_405 bl[405] br[405] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_406 bl[406] br[406] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_407 bl[407] br[407] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_408 bl[408] br[408] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_409 bl[409] br[409] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_410 bl[410] br[410] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_411 bl[411] br[411] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_412 bl[412] br[412] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_413 bl[413] br[413] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_414 bl[414] br[414] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_415 bl[415] br[415] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_416 bl[416] br[416] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_417 bl[417] br[417] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_418 bl[418] br[418] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_419 bl[419] br[419] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_420 bl[420] br[420] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_421 bl[421] br[421] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_422 bl[422] br[422] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_423 bl[423] br[423] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_424 bl[424] br[424] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_425 bl[425] br[425] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_426 bl[426] br[426] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_427 bl[427] br[427] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_428 bl[428] br[428] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_429 bl[429] br[429] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_430 bl[430] br[430] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_431 bl[431] br[431] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_432 bl[432] br[432] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_433 bl[433] br[433] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_434 bl[434] br[434] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_435 bl[435] br[435] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_436 bl[436] br[436] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_437 bl[437] br[437] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_438 bl[438] br[438] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_439 bl[439] br[439] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_440 bl[440] br[440] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_441 bl[441] br[441] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_442 bl[442] br[442] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_443 bl[443] br[443] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_444 bl[444] br[444] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_445 bl[445] br[445] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_446 bl[446] br[446] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_447 bl[447] br[447] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_448 bl[448] br[448] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_449 bl[449] br[449] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_450 bl[450] br[450] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_451 bl[451] br[451] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_452 bl[452] br[452] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_453 bl[453] br[453] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_454 bl[454] br[454] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_455 bl[455] br[455] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_456 bl[456] br[456] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_457 bl[457] br[457] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_458 bl[458] br[458] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_459 bl[459] br[459] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_460 bl[460] br[460] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_461 bl[461] br[461] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_462 bl[462] br[462] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_463 bl[463] br[463] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_464 bl[464] br[464] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_465 bl[465] br[465] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_466 bl[466] br[466] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_467 bl[467] br[467] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_468 bl[468] br[468] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_469 bl[469] br[469] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_470 bl[470] br[470] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_471 bl[471] br[471] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_472 bl[472] br[472] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_473 bl[473] br[473] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_474 bl[474] br[474] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_475 bl[475] br[475] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_476 bl[476] br[476] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_477 bl[477] br[477] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_478 bl[478] br[478] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_479 bl[479] br[479] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_480 bl[480] br[480] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_481 bl[481] br[481] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_482 bl[482] br[482] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_483 bl[483] br[483] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_484 bl[484] br[484] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_485 bl[485] br[485] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_486 bl[486] br[486] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_487 bl[487] br[487] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_488 bl[488] br[488] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_489 bl[489] br[489] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_490 bl[490] br[490] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_491 bl[491] br[491] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_492 bl[492] br[492] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_493 bl[493] br[493] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_494 bl[494] br[494] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_495 bl[495] br[495] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_496 bl[496] br[496] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_497 bl[497] br[497] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_498 bl[498] br[498] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_499 bl[499] br[499] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_500 bl[500] br[500] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_501 bl[501] br[501] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_502 bl[502] br[502] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_503 bl[503] br[503] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_504 bl[504] br[504] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_505 bl[505] br[505] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_506 bl[506] br[506] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_507 bl[507] br[507] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_508 bl[508] br[508] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_509 bl[509] br[509] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_510 bl[510] br[510] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_7_511 bl[511] br[511] vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xcell_8_0 bl[0] br[0] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_1 bl[1] br[1] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_2 bl[2] br[2] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_3 bl[3] br[3] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_4 bl[4] br[4] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_5 bl[5] br[5] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_6 bl[6] br[6] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_7 bl[7] br[7] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_8 bl[8] br[8] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_9 bl[9] br[9] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_10 bl[10] br[10] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_11 bl[11] br[11] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_12 bl[12] br[12] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_13 bl[13] br[13] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_14 bl[14] br[14] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_15 bl[15] br[15] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_16 bl[16] br[16] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_17 bl[17] br[17] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_18 bl[18] br[18] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_19 bl[19] br[19] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_20 bl[20] br[20] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_21 bl[21] br[21] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_22 bl[22] br[22] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_23 bl[23] br[23] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_24 bl[24] br[24] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_25 bl[25] br[25] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_26 bl[26] br[26] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_27 bl[27] br[27] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_28 bl[28] br[28] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_29 bl[29] br[29] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_30 bl[30] br[30] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_31 bl[31] br[31] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_32 bl[32] br[32] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_33 bl[33] br[33] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_34 bl[34] br[34] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_35 bl[35] br[35] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_36 bl[36] br[36] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_37 bl[37] br[37] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_38 bl[38] br[38] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_39 bl[39] br[39] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_40 bl[40] br[40] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_41 bl[41] br[41] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_42 bl[42] br[42] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_43 bl[43] br[43] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_44 bl[44] br[44] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_45 bl[45] br[45] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_46 bl[46] br[46] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_47 bl[47] br[47] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_48 bl[48] br[48] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_49 bl[49] br[49] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_50 bl[50] br[50] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_51 bl[51] br[51] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_52 bl[52] br[52] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_53 bl[53] br[53] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_54 bl[54] br[54] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_55 bl[55] br[55] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_56 bl[56] br[56] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_57 bl[57] br[57] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_58 bl[58] br[58] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_59 bl[59] br[59] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_60 bl[60] br[60] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_61 bl[61] br[61] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_62 bl[62] br[62] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_63 bl[63] br[63] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_64 bl[64] br[64] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_65 bl[65] br[65] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_66 bl[66] br[66] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_67 bl[67] br[67] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_68 bl[68] br[68] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_69 bl[69] br[69] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_70 bl[70] br[70] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_71 bl[71] br[71] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_72 bl[72] br[72] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_73 bl[73] br[73] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_74 bl[74] br[74] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_75 bl[75] br[75] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_76 bl[76] br[76] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_77 bl[77] br[77] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_78 bl[78] br[78] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_79 bl[79] br[79] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_80 bl[80] br[80] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_81 bl[81] br[81] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_82 bl[82] br[82] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_83 bl[83] br[83] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_84 bl[84] br[84] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_85 bl[85] br[85] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_86 bl[86] br[86] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_87 bl[87] br[87] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_88 bl[88] br[88] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_89 bl[89] br[89] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_90 bl[90] br[90] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_91 bl[91] br[91] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_92 bl[92] br[92] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_93 bl[93] br[93] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_94 bl[94] br[94] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_95 bl[95] br[95] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_96 bl[96] br[96] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_97 bl[97] br[97] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_98 bl[98] br[98] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_99 bl[99] br[99] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_100 bl[100] br[100] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_101 bl[101] br[101] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_102 bl[102] br[102] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_103 bl[103] br[103] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_104 bl[104] br[104] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_105 bl[105] br[105] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_106 bl[106] br[106] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_107 bl[107] br[107] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_108 bl[108] br[108] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_109 bl[109] br[109] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_110 bl[110] br[110] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_111 bl[111] br[111] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_112 bl[112] br[112] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_113 bl[113] br[113] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_114 bl[114] br[114] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_115 bl[115] br[115] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_116 bl[116] br[116] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_117 bl[117] br[117] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_118 bl[118] br[118] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_119 bl[119] br[119] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_120 bl[120] br[120] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_121 bl[121] br[121] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_122 bl[122] br[122] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_123 bl[123] br[123] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_124 bl[124] br[124] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_125 bl[125] br[125] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_126 bl[126] br[126] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_127 bl[127] br[127] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_128 bl[128] br[128] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_129 bl[129] br[129] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_130 bl[130] br[130] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_131 bl[131] br[131] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_132 bl[132] br[132] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_133 bl[133] br[133] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_134 bl[134] br[134] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_135 bl[135] br[135] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_136 bl[136] br[136] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_137 bl[137] br[137] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_138 bl[138] br[138] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_139 bl[139] br[139] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_140 bl[140] br[140] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_141 bl[141] br[141] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_142 bl[142] br[142] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_143 bl[143] br[143] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_144 bl[144] br[144] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_145 bl[145] br[145] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_146 bl[146] br[146] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_147 bl[147] br[147] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_148 bl[148] br[148] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_149 bl[149] br[149] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_150 bl[150] br[150] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_151 bl[151] br[151] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_152 bl[152] br[152] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_153 bl[153] br[153] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_154 bl[154] br[154] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_155 bl[155] br[155] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_156 bl[156] br[156] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_157 bl[157] br[157] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_158 bl[158] br[158] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_159 bl[159] br[159] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_160 bl[160] br[160] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_161 bl[161] br[161] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_162 bl[162] br[162] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_163 bl[163] br[163] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_164 bl[164] br[164] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_165 bl[165] br[165] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_166 bl[166] br[166] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_167 bl[167] br[167] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_168 bl[168] br[168] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_169 bl[169] br[169] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_170 bl[170] br[170] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_171 bl[171] br[171] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_172 bl[172] br[172] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_173 bl[173] br[173] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_174 bl[174] br[174] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_175 bl[175] br[175] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_176 bl[176] br[176] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_177 bl[177] br[177] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_178 bl[178] br[178] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_179 bl[179] br[179] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_180 bl[180] br[180] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_181 bl[181] br[181] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_182 bl[182] br[182] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_183 bl[183] br[183] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_184 bl[184] br[184] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_185 bl[185] br[185] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_186 bl[186] br[186] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_187 bl[187] br[187] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_188 bl[188] br[188] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_189 bl[189] br[189] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_190 bl[190] br[190] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_191 bl[191] br[191] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_192 bl[192] br[192] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_193 bl[193] br[193] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_194 bl[194] br[194] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_195 bl[195] br[195] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_196 bl[196] br[196] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_197 bl[197] br[197] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_198 bl[198] br[198] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_199 bl[199] br[199] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_200 bl[200] br[200] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_201 bl[201] br[201] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_202 bl[202] br[202] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_203 bl[203] br[203] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_204 bl[204] br[204] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_205 bl[205] br[205] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_206 bl[206] br[206] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_207 bl[207] br[207] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_208 bl[208] br[208] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_209 bl[209] br[209] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_210 bl[210] br[210] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_211 bl[211] br[211] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_212 bl[212] br[212] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_213 bl[213] br[213] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_214 bl[214] br[214] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_215 bl[215] br[215] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_216 bl[216] br[216] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_217 bl[217] br[217] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_218 bl[218] br[218] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_219 bl[219] br[219] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_220 bl[220] br[220] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_221 bl[221] br[221] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_222 bl[222] br[222] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_223 bl[223] br[223] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_224 bl[224] br[224] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_225 bl[225] br[225] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_226 bl[226] br[226] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_227 bl[227] br[227] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_228 bl[228] br[228] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_229 bl[229] br[229] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_230 bl[230] br[230] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_231 bl[231] br[231] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_232 bl[232] br[232] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_233 bl[233] br[233] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_234 bl[234] br[234] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_235 bl[235] br[235] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_236 bl[236] br[236] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_237 bl[237] br[237] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_238 bl[238] br[238] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_239 bl[239] br[239] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_240 bl[240] br[240] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_241 bl[241] br[241] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_242 bl[242] br[242] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_243 bl[243] br[243] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_244 bl[244] br[244] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_245 bl[245] br[245] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_246 bl[246] br[246] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_247 bl[247] br[247] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_248 bl[248] br[248] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_249 bl[249] br[249] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_250 bl[250] br[250] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_251 bl[251] br[251] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_252 bl[252] br[252] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_253 bl[253] br[253] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_254 bl[254] br[254] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_255 bl[255] br[255] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_256 bl[256] br[256] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_257 bl[257] br[257] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_258 bl[258] br[258] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_259 bl[259] br[259] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_260 bl[260] br[260] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_261 bl[261] br[261] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_262 bl[262] br[262] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_263 bl[263] br[263] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_264 bl[264] br[264] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_265 bl[265] br[265] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_266 bl[266] br[266] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_267 bl[267] br[267] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_268 bl[268] br[268] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_269 bl[269] br[269] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_270 bl[270] br[270] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_271 bl[271] br[271] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_272 bl[272] br[272] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_273 bl[273] br[273] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_274 bl[274] br[274] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_275 bl[275] br[275] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_276 bl[276] br[276] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_277 bl[277] br[277] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_278 bl[278] br[278] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_279 bl[279] br[279] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_280 bl[280] br[280] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_281 bl[281] br[281] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_282 bl[282] br[282] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_283 bl[283] br[283] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_284 bl[284] br[284] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_285 bl[285] br[285] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_286 bl[286] br[286] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_287 bl[287] br[287] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_288 bl[288] br[288] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_289 bl[289] br[289] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_290 bl[290] br[290] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_291 bl[291] br[291] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_292 bl[292] br[292] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_293 bl[293] br[293] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_294 bl[294] br[294] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_295 bl[295] br[295] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_296 bl[296] br[296] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_297 bl[297] br[297] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_298 bl[298] br[298] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_299 bl[299] br[299] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_300 bl[300] br[300] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_301 bl[301] br[301] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_302 bl[302] br[302] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_303 bl[303] br[303] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_304 bl[304] br[304] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_305 bl[305] br[305] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_306 bl[306] br[306] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_307 bl[307] br[307] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_308 bl[308] br[308] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_309 bl[309] br[309] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_310 bl[310] br[310] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_311 bl[311] br[311] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_312 bl[312] br[312] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_313 bl[313] br[313] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_314 bl[314] br[314] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_315 bl[315] br[315] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_316 bl[316] br[316] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_317 bl[317] br[317] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_318 bl[318] br[318] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_319 bl[319] br[319] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_320 bl[320] br[320] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_321 bl[321] br[321] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_322 bl[322] br[322] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_323 bl[323] br[323] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_324 bl[324] br[324] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_325 bl[325] br[325] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_326 bl[326] br[326] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_327 bl[327] br[327] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_328 bl[328] br[328] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_329 bl[329] br[329] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_330 bl[330] br[330] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_331 bl[331] br[331] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_332 bl[332] br[332] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_333 bl[333] br[333] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_334 bl[334] br[334] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_335 bl[335] br[335] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_336 bl[336] br[336] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_337 bl[337] br[337] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_338 bl[338] br[338] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_339 bl[339] br[339] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_340 bl[340] br[340] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_341 bl[341] br[341] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_342 bl[342] br[342] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_343 bl[343] br[343] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_344 bl[344] br[344] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_345 bl[345] br[345] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_346 bl[346] br[346] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_347 bl[347] br[347] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_348 bl[348] br[348] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_349 bl[349] br[349] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_350 bl[350] br[350] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_351 bl[351] br[351] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_352 bl[352] br[352] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_353 bl[353] br[353] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_354 bl[354] br[354] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_355 bl[355] br[355] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_356 bl[356] br[356] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_357 bl[357] br[357] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_358 bl[358] br[358] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_359 bl[359] br[359] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_360 bl[360] br[360] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_361 bl[361] br[361] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_362 bl[362] br[362] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_363 bl[363] br[363] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_364 bl[364] br[364] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_365 bl[365] br[365] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_366 bl[366] br[366] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_367 bl[367] br[367] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_368 bl[368] br[368] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_369 bl[369] br[369] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_370 bl[370] br[370] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_371 bl[371] br[371] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_372 bl[372] br[372] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_373 bl[373] br[373] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_374 bl[374] br[374] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_375 bl[375] br[375] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_376 bl[376] br[376] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_377 bl[377] br[377] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_378 bl[378] br[378] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_379 bl[379] br[379] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_380 bl[380] br[380] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_381 bl[381] br[381] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_382 bl[382] br[382] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_383 bl[383] br[383] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_384 bl[384] br[384] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_385 bl[385] br[385] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_386 bl[386] br[386] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_387 bl[387] br[387] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_388 bl[388] br[388] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_389 bl[389] br[389] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_390 bl[390] br[390] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_391 bl[391] br[391] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_392 bl[392] br[392] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_393 bl[393] br[393] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_394 bl[394] br[394] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_395 bl[395] br[395] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_396 bl[396] br[396] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_397 bl[397] br[397] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_398 bl[398] br[398] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_399 bl[399] br[399] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_400 bl[400] br[400] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_401 bl[401] br[401] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_402 bl[402] br[402] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_403 bl[403] br[403] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_404 bl[404] br[404] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_405 bl[405] br[405] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_406 bl[406] br[406] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_407 bl[407] br[407] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_408 bl[408] br[408] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_409 bl[409] br[409] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_410 bl[410] br[410] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_411 bl[411] br[411] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_412 bl[412] br[412] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_413 bl[413] br[413] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_414 bl[414] br[414] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_415 bl[415] br[415] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_416 bl[416] br[416] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_417 bl[417] br[417] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_418 bl[418] br[418] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_419 bl[419] br[419] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_420 bl[420] br[420] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_421 bl[421] br[421] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_422 bl[422] br[422] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_423 bl[423] br[423] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_424 bl[424] br[424] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_425 bl[425] br[425] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_426 bl[426] br[426] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_427 bl[427] br[427] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_428 bl[428] br[428] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_429 bl[429] br[429] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_430 bl[430] br[430] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_431 bl[431] br[431] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_432 bl[432] br[432] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_433 bl[433] br[433] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_434 bl[434] br[434] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_435 bl[435] br[435] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_436 bl[436] br[436] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_437 bl[437] br[437] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_438 bl[438] br[438] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_439 bl[439] br[439] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_440 bl[440] br[440] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_441 bl[441] br[441] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_442 bl[442] br[442] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_443 bl[443] br[443] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_444 bl[444] br[444] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_445 bl[445] br[445] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_446 bl[446] br[446] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_447 bl[447] br[447] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_448 bl[448] br[448] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_449 bl[449] br[449] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_450 bl[450] br[450] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_451 bl[451] br[451] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_452 bl[452] br[452] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_453 bl[453] br[453] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_454 bl[454] br[454] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_455 bl[455] br[455] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_456 bl[456] br[456] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_457 bl[457] br[457] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_458 bl[458] br[458] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_459 bl[459] br[459] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_460 bl[460] br[460] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_461 bl[461] br[461] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_462 bl[462] br[462] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_463 bl[463] br[463] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_464 bl[464] br[464] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_465 bl[465] br[465] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_466 bl[466] br[466] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_467 bl[467] br[467] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_468 bl[468] br[468] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_469 bl[469] br[469] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_470 bl[470] br[470] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_471 bl[471] br[471] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_472 bl[472] br[472] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_473 bl[473] br[473] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_474 bl[474] br[474] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_475 bl[475] br[475] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_476 bl[476] br[476] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_477 bl[477] br[477] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_478 bl[478] br[478] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_479 bl[479] br[479] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_480 bl[480] br[480] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_481 bl[481] br[481] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_482 bl[482] br[482] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_483 bl[483] br[483] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_484 bl[484] br[484] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_485 bl[485] br[485] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_486 bl[486] br[486] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_487 bl[487] br[487] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_488 bl[488] br[488] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_489 bl[489] br[489] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_490 bl[490] br[490] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_491 bl[491] br[491] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_492 bl[492] br[492] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_493 bl[493] br[493] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_494 bl[494] br[494] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_495 bl[495] br[495] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_496 bl[496] br[496] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_497 bl[497] br[497] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_498 bl[498] br[498] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_499 bl[499] br[499] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_500 bl[500] br[500] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_501 bl[501] br[501] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_502 bl[502] br[502] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_503 bl[503] br[503] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_504 bl[504] br[504] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_505 bl[505] br[505] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_506 bl[506] br[506] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_507 bl[507] br[507] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_508 bl[508] br[508] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_509 bl[509] br[509] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_510 bl[510] br[510] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_8_511 bl[511] br[511] vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xcell_9_0 bl[0] br[0] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_1 bl[1] br[1] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_2 bl[2] br[2] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_3 bl[3] br[3] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_4 bl[4] br[4] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_5 bl[5] br[5] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_6 bl[6] br[6] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_7 bl[7] br[7] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_8 bl[8] br[8] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_9 bl[9] br[9] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_10 bl[10] br[10] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_11 bl[11] br[11] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_12 bl[12] br[12] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_13 bl[13] br[13] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_14 bl[14] br[14] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_15 bl[15] br[15] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_16 bl[16] br[16] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_17 bl[17] br[17] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_18 bl[18] br[18] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_19 bl[19] br[19] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_20 bl[20] br[20] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_21 bl[21] br[21] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_22 bl[22] br[22] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_23 bl[23] br[23] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_24 bl[24] br[24] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_25 bl[25] br[25] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_26 bl[26] br[26] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_27 bl[27] br[27] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_28 bl[28] br[28] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_29 bl[29] br[29] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_30 bl[30] br[30] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_31 bl[31] br[31] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_32 bl[32] br[32] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_33 bl[33] br[33] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_34 bl[34] br[34] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_35 bl[35] br[35] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_36 bl[36] br[36] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_37 bl[37] br[37] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_38 bl[38] br[38] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_39 bl[39] br[39] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_40 bl[40] br[40] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_41 bl[41] br[41] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_42 bl[42] br[42] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_43 bl[43] br[43] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_44 bl[44] br[44] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_45 bl[45] br[45] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_46 bl[46] br[46] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_47 bl[47] br[47] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_48 bl[48] br[48] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_49 bl[49] br[49] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_50 bl[50] br[50] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_51 bl[51] br[51] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_52 bl[52] br[52] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_53 bl[53] br[53] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_54 bl[54] br[54] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_55 bl[55] br[55] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_56 bl[56] br[56] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_57 bl[57] br[57] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_58 bl[58] br[58] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_59 bl[59] br[59] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_60 bl[60] br[60] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_61 bl[61] br[61] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_62 bl[62] br[62] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_63 bl[63] br[63] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_64 bl[64] br[64] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_65 bl[65] br[65] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_66 bl[66] br[66] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_67 bl[67] br[67] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_68 bl[68] br[68] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_69 bl[69] br[69] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_70 bl[70] br[70] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_71 bl[71] br[71] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_72 bl[72] br[72] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_73 bl[73] br[73] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_74 bl[74] br[74] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_75 bl[75] br[75] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_76 bl[76] br[76] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_77 bl[77] br[77] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_78 bl[78] br[78] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_79 bl[79] br[79] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_80 bl[80] br[80] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_81 bl[81] br[81] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_82 bl[82] br[82] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_83 bl[83] br[83] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_84 bl[84] br[84] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_85 bl[85] br[85] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_86 bl[86] br[86] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_87 bl[87] br[87] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_88 bl[88] br[88] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_89 bl[89] br[89] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_90 bl[90] br[90] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_91 bl[91] br[91] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_92 bl[92] br[92] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_93 bl[93] br[93] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_94 bl[94] br[94] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_95 bl[95] br[95] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_96 bl[96] br[96] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_97 bl[97] br[97] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_98 bl[98] br[98] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_99 bl[99] br[99] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_100 bl[100] br[100] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_101 bl[101] br[101] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_102 bl[102] br[102] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_103 bl[103] br[103] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_104 bl[104] br[104] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_105 bl[105] br[105] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_106 bl[106] br[106] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_107 bl[107] br[107] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_108 bl[108] br[108] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_109 bl[109] br[109] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_110 bl[110] br[110] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_111 bl[111] br[111] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_112 bl[112] br[112] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_113 bl[113] br[113] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_114 bl[114] br[114] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_115 bl[115] br[115] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_116 bl[116] br[116] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_117 bl[117] br[117] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_118 bl[118] br[118] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_119 bl[119] br[119] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_120 bl[120] br[120] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_121 bl[121] br[121] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_122 bl[122] br[122] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_123 bl[123] br[123] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_124 bl[124] br[124] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_125 bl[125] br[125] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_126 bl[126] br[126] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_127 bl[127] br[127] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_128 bl[128] br[128] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_129 bl[129] br[129] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_130 bl[130] br[130] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_131 bl[131] br[131] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_132 bl[132] br[132] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_133 bl[133] br[133] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_134 bl[134] br[134] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_135 bl[135] br[135] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_136 bl[136] br[136] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_137 bl[137] br[137] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_138 bl[138] br[138] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_139 bl[139] br[139] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_140 bl[140] br[140] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_141 bl[141] br[141] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_142 bl[142] br[142] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_143 bl[143] br[143] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_144 bl[144] br[144] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_145 bl[145] br[145] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_146 bl[146] br[146] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_147 bl[147] br[147] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_148 bl[148] br[148] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_149 bl[149] br[149] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_150 bl[150] br[150] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_151 bl[151] br[151] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_152 bl[152] br[152] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_153 bl[153] br[153] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_154 bl[154] br[154] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_155 bl[155] br[155] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_156 bl[156] br[156] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_157 bl[157] br[157] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_158 bl[158] br[158] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_159 bl[159] br[159] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_160 bl[160] br[160] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_161 bl[161] br[161] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_162 bl[162] br[162] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_163 bl[163] br[163] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_164 bl[164] br[164] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_165 bl[165] br[165] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_166 bl[166] br[166] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_167 bl[167] br[167] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_168 bl[168] br[168] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_169 bl[169] br[169] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_170 bl[170] br[170] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_171 bl[171] br[171] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_172 bl[172] br[172] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_173 bl[173] br[173] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_174 bl[174] br[174] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_175 bl[175] br[175] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_176 bl[176] br[176] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_177 bl[177] br[177] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_178 bl[178] br[178] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_179 bl[179] br[179] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_180 bl[180] br[180] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_181 bl[181] br[181] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_182 bl[182] br[182] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_183 bl[183] br[183] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_184 bl[184] br[184] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_185 bl[185] br[185] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_186 bl[186] br[186] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_187 bl[187] br[187] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_188 bl[188] br[188] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_189 bl[189] br[189] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_190 bl[190] br[190] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_191 bl[191] br[191] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_192 bl[192] br[192] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_193 bl[193] br[193] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_194 bl[194] br[194] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_195 bl[195] br[195] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_196 bl[196] br[196] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_197 bl[197] br[197] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_198 bl[198] br[198] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_199 bl[199] br[199] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_200 bl[200] br[200] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_201 bl[201] br[201] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_202 bl[202] br[202] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_203 bl[203] br[203] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_204 bl[204] br[204] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_205 bl[205] br[205] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_206 bl[206] br[206] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_207 bl[207] br[207] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_208 bl[208] br[208] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_209 bl[209] br[209] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_210 bl[210] br[210] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_211 bl[211] br[211] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_212 bl[212] br[212] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_213 bl[213] br[213] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_214 bl[214] br[214] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_215 bl[215] br[215] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_216 bl[216] br[216] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_217 bl[217] br[217] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_218 bl[218] br[218] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_219 bl[219] br[219] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_220 bl[220] br[220] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_221 bl[221] br[221] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_222 bl[222] br[222] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_223 bl[223] br[223] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_224 bl[224] br[224] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_225 bl[225] br[225] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_226 bl[226] br[226] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_227 bl[227] br[227] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_228 bl[228] br[228] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_229 bl[229] br[229] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_230 bl[230] br[230] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_231 bl[231] br[231] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_232 bl[232] br[232] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_233 bl[233] br[233] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_234 bl[234] br[234] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_235 bl[235] br[235] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_236 bl[236] br[236] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_237 bl[237] br[237] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_238 bl[238] br[238] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_239 bl[239] br[239] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_240 bl[240] br[240] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_241 bl[241] br[241] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_242 bl[242] br[242] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_243 bl[243] br[243] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_244 bl[244] br[244] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_245 bl[245] br[245] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_246 bl[246] br[246] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_247 bl[247] br[247] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_248 bl[248] br[248] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_249 bl[249] br[249] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_250 bl[250] br[250] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_251 bl[251] br[251] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_252 bl[252] br[252] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_253 bl[253] br[253] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_254 bl[254] br[254] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_255 bl[255] br[255] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_256 bl[256] br[256] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_257 bl[257] br[257] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_258 bl[258] br[258] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_259 bl[259] br[259] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_260 bl[260] br[260] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_261 bl[261] br[261] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_262 bl[262] br[262] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_263 bl[263] br[263] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_264 bl[264] br[264] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_265 bl[265] br[265] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_266 bl[266] br[266] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_267 bl[267] br[267] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_268 bl[268] br[268] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_269 bl[269] br[269] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_270 bl[270] br[270] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_271 bl[271] br[271] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_272 bl[272] br[272] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_273 bl[273] br[273] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_274 bl[274] br[274] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_275 bl[275] br[275] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_276 bl[276] br[276] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_277 bl[277] br[277] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_278 bl[278] br[278] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_279 bl[279] br[279] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_280 bl[280] br[280] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_281 bl[281] br[281] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_282 bl[282] br[282] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_283 bl[283] br[283] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_284 bl[284] br[284] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_285 bl[285] br[285] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_286 bl[286] br[286] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_287 bl[287] br[287] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_288 bl[288] br[288] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_289 bl[289] br[289] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_290 bl[290] br[290] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_291 bl[291] br[291] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_292 bl[292] br[292] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_293 bl[293] br[293] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_294 bl[294] br[294] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_295 bl[295] br[295] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_296 bl[296] br[296] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_297 bl[297] br[297] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_298 bl[298] br[298] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_299 bl[299] br[299] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_300 bl[300] br[300] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_301 bl[301] br[301] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_302 bl[302] br[302] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_303 bl[303] br[303] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_304 bl[304] br[304] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_305 bl[305] br[305] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_306 bl[306] br[306] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_307 bl[307] br[307] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_308 bl[308] br[308] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_309 bl[309] br[309] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_310 bl[310] br[310] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_311 bl[311] br[311] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_312 bl[312] br[312] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_313 bl[313] br[313] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_314 bl[314] br[314] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_315 bl[315] br[315] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_316 bl[316] br[316] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_317 bl[317] br[317] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_318 bl[318] br[318] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_319 bl[319] br[319] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_320 bl[320] br[320] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_321 bl[321] br[321] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_322 bl[322] br[322] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_323 bl[323] br[323] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_324 bl[324] br[324] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_325 bl[325] br[325] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_326 bl[326] br[326] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_327 bl[327] br[327] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_328 bl[328] br[328] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_329 bl[329] br[329] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_330 bl[330] br[330] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_331 bl[331] br[331] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_332 bl[332] br[332] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_333 bl[333] br[333] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_334 bl[334] br[334] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_335 bl[335] br[335] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_336 bl[336] br[336] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_337 bl[337] br[337] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_338 bl[338] br[338] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_339 bl[339] br[339] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_340 bl[340] br[340] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_341 bl[341] br[341] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_342 bl[342] br[342] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_343 bl[343] br[343] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_344 bl[344] br[344] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_345 bl[345] br[345] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_346 bl[346] br[346] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_347 bl[347] br[347] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_348 bl[348] br[348] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_349 bl[349] br[349] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_350 bl[350] br[350] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_351 bl[351] br[351] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_352 bl[352] br[352] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_353 bl[353] br[353] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_354 bl[354] br[354] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_355 bl[355] br[355] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_356 bl[356] br[356] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_357 bl[357] br[357] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_358 bl[358] br[358] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_359 bl[359] br[359] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_360 bl[360] br[360] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_361 bl[361] br[361] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_362 bl[362] br[362] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_363 bl[363] br[363] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_364 bl[364] br[364] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_365 bl[365] br[365] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_366 bl[366] br[366] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_367 bl[367] br[367] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_368 bl[368] br[368] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_369 bl[369] br[369] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_370 bl[370] br[370] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_371 bl[371] br[371] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_372 bl[372] br[372] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_373 bl[373] br[373] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_374 bl[374] br[374] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_375 bl[375] br[375] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_376 bl[376] br[376] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_377 bl[377] br[377] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_378 bl[378] br[378] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_379 bl[379] br[379] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_380 bl[380] br[380] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_381 bl[381] br[381] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_382 bl[382] br[382] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_383 bl[383] br[383] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_384 bl[384] br[384] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_385 bl[385] br[385] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_386 bl[386] br[386] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_387 bl[387] br[387] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_388 bl[388] br[388] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_389 bl[389] br[389] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_390 bl[390] br[390] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_391 bl[391] br[391] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_392 bl[392] br[392] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_393 bl[393] br[393] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_394 bl[394] br[394] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_395 bl[395] br[395] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_396 bl[396] br[396] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_397 bl[397] br[397] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_398 bl[398] br[398] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_399 bl[399] br[399] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_400 bl[400] br[400] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_401 bl[401] br[401] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_402 bl[402] br[402] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_403 bl[403] br[403] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_404 bl[404] br[404] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_405 bl[405] br[405] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_406 bl[406] br[406] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_407 bl[407] br[407] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_408 bl[408] br[408] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_409 bl[409] br[409] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_410 bl[410] br[410] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_411 bl[411] br[411] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_412 bl[412] br[412] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_413 bl[413] br[413] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_414 bl[414] br[414] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_415 bl[415] br[415] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_416 bl[416] br[416] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_417 bl[417] br[417] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_418 bl[418] br[418] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_419 bl[419] br[419] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_420 bl[420] br[420] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_421 bl[421] br[421] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_422 bl[422] br[422] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_423 bl[423] br[423] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_424 bl[424] br[424] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_425 bl[425] br[425] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_426 bl[426] br[426] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_427 bl[427] br[427] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_428 bl[428] br[428] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_429 bl[429] br[429] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_430 bl[430] br[430] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_431 bl[431] br[431] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_432 bl[432] br[432] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_433 bl[433] br[433] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_434 bl[434] br[434] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_435 bl[435] br[435] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_436 bl[436] br[436] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_437 bl[437] br[437] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_438 bl[438] br[438] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_439 bl[439] br[439] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_440 bl[440] br[440] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_441 bl[441] br[441] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_442 bl[442] br[442] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_443 bl[443] br[443] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_444 bl[444] br[444] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_445 bl[445] br[445] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_446 bl[446] br[446] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_447 bl[447] br[447] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_448 bl[448] br[448] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_449 bl[449] br[449] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_450 bl[450] br[450] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_451 bl[451] br[451] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_452 bl[452] br[452] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_453 bl[453] br[453] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_454 bl[454] br[454] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_455 bl[455] br[455] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_456 bl[456] br[456] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_457 bl[457] br[457] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_458 bl[458] br[458] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_459 bl[459] br[459] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_460 bl[460] br[460] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_461 bl[461] br[461] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_462 bl[462] br[462] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_463 bl[463] br[463] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_464 bl[464] br[464] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_465 bl[465] br[465] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_466 bl[466] br[466] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_467 bl[467] br[467] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_468 bl[468] br[468] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_469 bl[469] br[469] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_470 bl[470] br[470] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_471 bl[471] br[471] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_472 bl[472] br[472] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_473 bl[473] br[473] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_474 bl[474] br[474] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_475 bl[475] br[475] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_476 bl[476] br[476] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_477 bl[477] br[477] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_478 bl[478] br[478] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_479 bl[479] br[479] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_480 bl[480] br[480] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_481 bl[481] br[481] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_482 bl[482] br[482] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_483 bl[483] br[483] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_484 bl[484] br[484] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_485 bl[485] br[485] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_486 bl[486] br[486] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_487 bl[487] br[487] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_488 bl[488] br[488] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_489 bl[489] br[489] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_490 bl[490] br[490] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_491 bl[491] br[491] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_492 bl[492] br[492] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_493 bl[493] br[493] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_494 bl[494] br[494] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_495 bl[495] br[495] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_496 bl[496] br[496] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_497 bl[497] br[497] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_498 bl[498] br[498] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_499 bl[499] br[499] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_500 bl[500] br[500] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_501 bl[501] br[501] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_502 bl[502] br[502] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_503 bl[503] br[503] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_504 bl[504] br[504] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_505 bl[505] br[505] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_506 bl[506] br[506] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_507 bl[507] br[507] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_508 bl[508] br[508] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_509 bl[509] br[509] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_510 bl[510] br[510] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_9_511 bl[511] br[511] vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xcell_10_0 bl[0] br[0] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_1 bl[1] br[1] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_2 bl[2] br[2] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_3 bl[3] br[3] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_4 bl[4] br[4] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_5 bl[5] br[5] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_6 bl[6] br[6] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_7 bl[7] br[7] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_8 bl[8] br[8] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_9 bl[9] br[9] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_10 bl[10] br[10] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_11 bl[11] br[11] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_12 bl[12] br[12] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_13 bl[13] br[13] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_14 bl[14] br[14] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_15 bl[15] br[15] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_16 bl[16] br[16] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_17 bl[17] br[17] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_18 bl[18] br[18] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_19 bl[19] br[19] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_20 bl[20] br[20] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_21 bl[21] br[21] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_22 bl[22] br[22] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_23 bl[23] br[23] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_24 bl[24] br[24] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_25 bl[25] br[25] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_26 bl[26] br[26] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_27 bl[27] br[27] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_28 bl[28] br[28] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_29 bl[29] br[29] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_30 bl[30] br[30] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_31 bl[31] br[31] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_32 bl[32] br[32] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_33 bl[33] br[33] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_34 bl[34] br[34] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_35 bl[35] br[35] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_36 bl[36] br[36] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_37 bl[37] br[37] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_38 bl[38] br[38] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_39 bl[39] br[39] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_40 bl[40] br[40] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_41 bl[41] br[41] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_42 bl[42] br[42] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_43 bl[43] br[43] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_44 bl[44] br[44] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_45 bl[45] br[45] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_46 bl[46] br[46] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_47 bl[47] br[47] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_48 bl[48] br[48] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_49 bl[49] br[49] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_50 bl[50] br[50] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_51 bl[51] br[51] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_52 bl[52] br[52] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_53 bl[53] br[53] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_54 bl[54] br[54] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_55 bl[55] br[55] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_56 bl[56] br[56] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_57 bl[57] br[57] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_58 bl[58] br[58] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_59 bl[59] br[59] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_60 bl[60] br[60] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_61 bl[61] br[61] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_62 bl[62] br[62] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_63 bl[63] br[63] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_64 bl[64] br[64] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_65 bl[65] br[65] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_66 bl[66] br[66] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_67 bl[67] br[67] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_68 bl[68] br[68] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_69 bl[69] br[69] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_70 bl[70] br[70] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_71 bl[71] br[71] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_72 bl[72] br[72] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_73 bl[73] br[73] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_74 bl[74] br[74] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_75 bl[75] br[75] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_76 bl[76] br[76] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_77 bl[77] br[77] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_78 bl[78] br[78] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_79 bl[79] br[79] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_80 bl[80] br[80] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_81 bl[81] br[81] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_82 bl[82] br[82] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_83 bl[83] br[83] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_84 bl[84] br[84] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_85 bl[85] br[85] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_86 bl[86] br[86] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_87 bl[87] br[87] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_88 bl[88] br[88] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_89 bl[89] br[89] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_90 bl[90] br[90] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_91 bl[91] br[91] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_92 bl[92] br[92] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_93 bl[93] br[93] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_94 bl[94] br[94] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_95 bl[95] br[95] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_96 bl[96] br[96] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_97 bl[97] br[97] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_98 bl[98] br[98] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_99 bl[99] br[99] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_100 bl[100] br[100] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_101 bl[101] br[101] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_102 bl[102] br[102] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_103 bl[103] br[103] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_104 bl[104] br[104] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_105 bl[105] br[105] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_106 bl[106] br[106] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_107 bl[107] br[107] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_108 bl[108] br[108] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_109 bl[109] br[109] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_110 bl[110] br[110] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_111 bl[111] br[111] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_112 bl[112] br[112] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_113 bl[113] br[113] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_114 bl[114] br[114] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_115 bl[115] br[115] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_116 bl[116] br[116] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_117 bl[117] br[117] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_118 bl[118] br[118] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_119 bl[119] br[119] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_120 bl[120] br[120] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_121 bl[121] br[121] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_122 bl[122] br[122] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_123 bl[123] br[123] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_124 bl[124] br[124] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_125 bl[125] br[125] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_126 bl[126] br[126] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_127 bl[127] br[127] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_128 bl[128] br[128] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_129 bl[129] br[129] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_130 bl[130] br[130] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_131 bl[131] br[131] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_132 bl[132] br[132] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_133 bl[133] br[133] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_134 bl[134] br[134] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_135 bl[135] br[135] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_136 bl[136] br[136] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_137 bl[137] br[137] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_138 bl[138] br[138] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_139 bl[139] br[139] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_140 bl[140] br[140] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_141 bl[141] br[141] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_142 bl[142] br[142] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_143 bl[143] br[143] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_144 bl[144] br[144] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_145 bl[145] br[145] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_146 bl[146] br[146] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_147 bl[147] br[147] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_148 bl[148] br[148] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_149 bl[149] br[149] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_150 bl[150] br[150] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_151 bl[151] br[151] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_152 bl[152] br[152] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_153 bl[153] br[153] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_154 bl[154] br[154] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_155 bl[155] br[155] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_156 bl[156] br[156] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_157 bl[157] br[157] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_158 bl[158] br[158] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_159 bl[159] br[159] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_160 bl[160] br[160] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_161 bl[161] br[161] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_162 bl[162] br[162] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_163 bl[163] br[163] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_164 bl[164] br[164] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_165 bl[165] br[165] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_166 bl[166] br[166] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_167 bl[167] br[167] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_168 bl[168] br[168] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_169 bl[169] br[169] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_170 bl[170] br[170] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_171 bl[171] br[171] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_172 bl[172] br[172] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_173 bl[173] br[173] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_174 bl[174] br[174] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_175 bl[175] br[175] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_176 bl[176] br[176] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_177 bl[177] br[177] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_178 bl[178] br[178] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_179 bl[179] br[179] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_180 bl[180] br[180] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_181 bl[181] br[181] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_182 bl[182] br[182] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_183 bl[183] br[183] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_184 bl[184] br[184] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_185 bl[185] br[185] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_186 bl[186] br[186] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_187 bl[187] br[187] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_188 bl[188] br[188] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_189 bl[189] br[189] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_190 bl[190] br[190] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_191 bl[191] br[191] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_192 bl[192] br[192] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_193 bl[193] br[193] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_194 bl[194] br[194] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_195 bl[195] br[195] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_196 bl[196] br[196] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_197 bl[197] br[197] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_198 bl[198] br[198] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_199 bl[199] br[199] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_200 bl[200] br[200] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_201 bl[201] br[201] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_202 bl[202] br[202] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_203 bl[203] br[203] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_204 bl[204] br[204] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_205 bl[205] br[205] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_206 bl[206] br[206] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_207 bl[207] br[207] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_208 bl[208] br[208] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_209 bl[209] br[209] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_210 bl[210] br[210] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_211 bl[211] br[211] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_212 bl[212] br[212] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_213 bl[213] br[213] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_214 bl[214] br[214] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_215 bl[215] br[215] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_216 bl[216] br[216] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_217 bl[217] br[217] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_218 bl[218] br[218] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_219 bl[219] br[219] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_220 bl[220] br[220] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_221 bl[221] br[221] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_222 bl[222] br[222] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_223 bl[223] br[223] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_224 bl[224] br[224] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_225 bl[225] br[225] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_226 bl[226] br[226] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_227 bl[227] br[227] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_228 bl[228] br[228] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_229 bl[229] br[229] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_230 bl[230] br[230] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_231 bl[231] br[231] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_232 bl[232] br[232] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_233 bl[233] br[233] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_234 bl[234] br[234] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_235 bl[235] br[235] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_236 bl[236] br[236] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_237 bl[237] br[237] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_238 bl[238] br[238] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_239 bl[239] br[239] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_240 bl[240] br[240] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_241 bl[241] br[241] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_242 bl[242] br[242] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_243 bl[243] br[243] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_244 bl[244] br[244] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_245 bl[245] br[245] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_246 bl[246] br[246] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_247 bl[247] br[247] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_248 bl[248] br[248] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_249 bl[249] br[249] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_250 bl[250] br[250] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_251 bl[251] br[251] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_252 bl[252] br[252] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_253 bl[253] br[253] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_254 bl[254] br[254] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_255 bl[255] br[255] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_256 bl[256] br[256] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_257 bl[257] br[257] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_258 bl[258] br[258] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_259 bl[259] br[259] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_260 bl[260] br[260] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_261 bl[261] br[261] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_262 bl[262] br[262] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_263 bl[263] br[263] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_264 bl[264] br[264] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_265 bl[265] br[265] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_266 bl[266] br[266] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_267 bl[267] br[267] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_268 bl[268] br[268] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_269 bl[269] br[269] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_270 bl[270] br[270] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_271 bl[271] br[271] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_272 bl[272] br[272] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_273 bl[273] br[273] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_274 bl[274] br[274] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_275 bl[275] br[275] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_276 bl[276] br[276] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_277 bl[277] br[277] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_278 bl[278] br[278] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_279 bl[279] br[279] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_280 bl[280] br[280] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_281 bl[281] br[281] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_282 bl[282] br[282] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_283 bl[283] br[283] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_284 bl[284] br[284] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_285 bl[285] br[285] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_286 bl[286] br[286] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_287 bl[287] br[287] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_288 bl[288] br[288] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_289 bl[289] br[289] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_290 bl[290] br[290] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_291 bl[291] br[291] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_292 bl[292] br[292] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_293 bl[293] br[293] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_294 bl[294] br[294] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_295 bl[295] br[295] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_296 bl[296] br[296] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_297 bl[297] br[297] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_298 bl[298] br[298] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_299 bl[299] br[299] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_300 bl[300] br[300] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_301 bl[301] br[301] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_302 bl[302] br[302] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_303 bl[303] br[303] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_304 bl[304] br[304] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_305 bl[305] br[305] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_306 bl[306] br[306] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_307 bl[307] br[307] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_308 bl[308] br[308] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_309 bl[309] br[309] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_310 bl[310] br[310] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_311 bl[311] br[311] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_312 bl[312] br[312] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_313 bl[313] br[313] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_314 bl[314] br[314] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_315 bl[315] br[315] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_316 bl[316] br[316] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_317 bl[317] br[317] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_318 bl[318] br[318] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_319 bl[319] br[319] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_320 bl[320] br[320] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_321 bl[321] br[321] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_322 bl[322] br[322] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_323 bl[323] br[323] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_324 bl[324] br[324] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_325 bl[325] br[325] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_326 bl[326] br[326] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_327 bl[327] br[327] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_328 bl[328] br[328] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_329 bl[329] br[329] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_330 bl[330] br[330] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_331 bl[331] br[331] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_332 bl[332] br[332] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_333 bl[333] br[333] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_334 bl[334] br[334] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_335 bl[335] br[335] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_336 bl[336] br[336] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_337 bl[337] br[337] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_338 bl[338] br[338] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_339 bl[339] br[339] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_340 bl[340] br[340] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_341 bl[341] br[341] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_342 bl[342] br[342] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_343 bl[343] br[343] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_344 bl[344] br[344] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_345 bl[345] br[345] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_346 bl[346] br[346] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_347 bl[347] br[347] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_348 bl[348] br[348] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_349 bl[349] br[349] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_350 bl[350] br[350] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_351 bl[351] br[351] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_352 bl[352] br[352] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_353 bl[353] br[353] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_354 bl[354] br[354] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_355 bl[355] br[355] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_356 bl[356] br[356] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_357 bl[357] br[357] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_358 bl[358] br[358] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_359 bl[359] br[359] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_360 bl[360] br[360] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_361 bl[361] br[361] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_362 bl[362] br[362] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_363 bl[363] br[363] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_364 bl[364] br[364] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_365 bl[365] br[365] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_366 bl[366] br[366] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_367 bl[367] br[367] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_368 bl[368] br[368] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_369 bl[369] br[369] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_370 bl[370] br[370] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_371 bl[371] br[371] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_372 bl[372] br[372] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_373 bl[373] br[373] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_374 bl[374] br[374] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_375 bl[375] br[375] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_376 bl[376] br[376] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_377 bl[377] br[377] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_378 bl[378] br[378] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_379 bl[379] br[379] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_380 bl[380] br[380] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_381 bl[381] br[381] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_382 bl[382] br[382] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_383 bl[383] br[383] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_384 bl[384] br[384] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_385 bl[385] br[385] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_386 bl[386] br[386] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_387 bl[387] br[387] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_388 bl[388] br[388] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_389 bl[389] br[389] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_390 bl[390] br[390] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_391 bl[391] br[391] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_392 bl[392] br[392] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_393 bl[393] br[393] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_394 bl[394] br[394] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_395 bl[395] br[395] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_396 bl[396] br[396] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_397 bl[397] br[397] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_398 bl[398] br[398] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_399 bl[399] br[399] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_400 bl[400] br[400] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_401 bl[401] br[401] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_402 bl[402] br[402] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_403 bl[403] br[403] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_404 bl[404] br[404] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_405 bl[405] br[405] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_406 bl[406] br[406] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_407 bl[407] br[407] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_408 bl[408] br[408] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_409 bl[409] br[409] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_410 bl[410] br[410] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_411 bl[411] br[411] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_412 bl[412] br[412] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_413 bl[413] br[413] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_414 bl[414] br[414] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_415 bl[415] br[415] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_416 bl[416] br[416] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_417 bl[417] br[417] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_418 bl[418] br[418] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_419 bl[419] br[419] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_420 bl[420] br[420] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_421 bl[421] br[421] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_422 bl[422] br[422] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_423 bl[423] br[423] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_424 bl[424] br[424] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_425 bl[425] br[425] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_426 bl[426] br[426] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_427 bl[427] br[427] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_428 bl[428] br[428] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_429 bl[429] br[429] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_430 bl[430] br[430] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_431 bl[431] br[431] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_432 bl[432] br[432] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_433 bl[433] br[433] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_434 bl[434] br[434] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_435 bl[435] br[435] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_436 bl[436] br[436] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_437 bl[437] br[437] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_438 bl[438] br[438] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_439 bl[439] br[439] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_440 bl[440] br[440] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_441 bl[441] br[441] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_442 bl[442] br[442] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_443 bl[443] br[443] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_444 bl[444] br[444] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_445 bl[445] br[445] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_446 bl[446] br[446] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_447 bl[447] br[447] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_448 bl[448] br[448] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_449 bl[449] br[449] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_450 bl[450] br[450] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_451 bl[451] br[451] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_452 bl[452] br[452] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_453 bl[453] br[453] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_454 bl[454] br[454] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_455 bl[455] br[455] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_456 bl[456] br[456] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_457 bl[457] br[457] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_458 bl[458] br[458] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_459 bl[459] br[459] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_460 bl[460] br[460] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_461 bl[461] br[461] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_462 bl[462] br[462] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_463 bl[463] br[463] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_464 bl[464] br[464] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_465 bl[465] br[465] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_466 bl[466] br[466] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_467 bl[467] br[467] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_468 bl[468] br[468] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_469 bl[469] br[469] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_470 bl[470] br[470] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_471 bl[471] br[471] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_472 bl[472] br[472] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_473 bl[473] br[473] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_474 bl[474] br[474] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_475 bl[475] br[475] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_476 bl[476] br[476] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_477 bl[477] br[477] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_478 bl[478] br[478] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_479 bl[479] br[479] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_480 bl[480] br[480] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_481 bl[481] br[481] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_482 bl[482] br[482] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_483 bl[483] br[483] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_484 bl[484] br[484] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_485 bl[485] br[485] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_486 bl[486] br[486] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_487 bl[487] br[487] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_488 bl[488] br[488] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_489 bl[489] br[489] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_490 bl[490] br[490] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_491 bl[491] br[491] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_492 bl[492] br[492] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_493 bl[493] br[493] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_494 bl[494] br[494] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_495 bl[495] br[495] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_496 bl[496] br[496] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_497 bl[497] br[497] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_498 bl[498] br[498] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_499 bl[499] br[499] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_500 bl[500] br[500] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_501 bl[501] br[501] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_502 bl[502] br[502] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_503 bl[503] br[503] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_504 bl[504] br[504] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_505 bl[505] br[505] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_506 bl[506] br[506] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_507 bl[507] br[507] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_508 bl[508] br[508] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_509 bl[509] br[509] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_510 bl[510] br[510] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_10_511 bl[511] br[511] vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xcell_11_0 bl[0] br[0] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_1 bl[1] br[1] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_2 bl[2] br[2] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_3 bl[3] br[3] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_4 bl[4] br[4] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_5 bl[5] br[5] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_6 bl[6] br[6] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_7 bl[7] br[7] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_8 bl[8] br[8] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_9 bl[9] br[9] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_10 bl[10] br[10] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_11 bl[11] br[11] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_12 bl[12] br[12] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_13 bl[13] br[13] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_14 bl[14] br[14] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_15 bl[15] br[15] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_16 bl[16] br[16] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_17 bl[17] br[17] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_18 bl[18] br[18] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_19 bl[19] br[19] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_20 bl[20] br[20] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_21 bl[21] br[21] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_22 bl[22] br[22] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_23 bl[23] br[23] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_24 bl[24] br[24] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_25 bl[25] br[25] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_26 bl[26] br[26] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_27 bl[27] br[27] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_28 bl[28] br[28] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_29 bl[29] br[29] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_30 bl[30] br[30] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_31 bl[31] br[31] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_32 bl[32] br[32] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_33 bl[33] br[33] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_34 bl[34] br[34] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_35 bl[35] br[35] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_36 bl[36] br[36] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_37 bl[37] br[37] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_38 bl[38] br[38] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_39 bl[39] br[39] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_40 bl[40] br[40] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_41 bl[41] br[41] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_42 bl[42] br[42] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_43 bl[43] br[43] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_44 bl[44] br[44] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_45 bl[45] br[45] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_46 bl[46] br[46] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_47 bl[47] br[47] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_48 bl[48] br[48] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_49 bl[49] br[49] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_50 bl[50] br[50] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_51 bl[51] br[51] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_52 bl[52] br[52] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_53 bl[53] br[53] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_54 bl[54] br[54] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_55 bl[55] br[55] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_56 bl[56] br[56] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_57 bl[57] br[57] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_58 bl[58] br[58] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_59 bl[59] br[59] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_60 bl[60] br[60] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_61 bl[61] br[61] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_62 bl[62] br[62] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_63 bl[63] br[63] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_64 bl[64] br[64] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_65 bl[65] br[65] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_66 bl[66] br[66] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_67 bl[67] br[67] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_68 bl[68] br[68] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_69 bl[69] br[69] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_70 bl[70] br[70] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_71 bl[71] br[71] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_72 bl[72] br[72] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_73 bl[73] br[73] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_74 bl[74] br[74] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_75 bl[75] br[75] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_76 bl[76] br[76] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_77 bl[77] br[77] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_78 bl[78] br[78] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_79 bl[79] br[79] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_80 bl[80] br[80] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_81 bl[81] br[81] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_82 bl[82] br[82] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_83 bl[83] br[83] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_84 bl[84] br[84] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_85 bl[85] br[85] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_86 bl[86] br[86] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_87 bl[87] br[87] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_88 bl[88] br[88] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_89 bl[89] br[89] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_90 bl[90] br[90] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_91 bl[91] br[91] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_92 bl[92] br[92] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_93 bl[93] br[93] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_94 bl[94] br[94] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_95 bl[95] br[95] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_96 bl[96] br[96] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_97 bl[97] br[97] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_98 bl[98] br[98] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_99 bl[99] br[99] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_100 bl[100] br[100] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_101 bl[101] br[101] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_102 bl[102] br[102] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_103 bl[103] br[103] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_104 bl[104] br[104] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_105 bl[105] br[105] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_106 bl[106] br[106] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_107 bl[107] br[107] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_108 bl[108] br[108] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_109 bl[109] br[109] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_110 bl[110] br[110] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_111 bl[111] br[111] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_112 bl[112] br[112] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_113 bl[113] br[113] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_114 bl[114] br[114] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_115 bl[115] br[115] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_116 bl[116] br[116] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_117 bl[117] br[117] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_118 bl[118] br[118] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_119 bl[119] br[119] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_120 bl[120] br[120] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_121 bl[121] br[121] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_122 bl[122] br[122] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_123 bl[123] br[123] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_124 bl[124] br[124] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_125 bl[125] br[125] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_126 bl[126] br[126] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_127 bl[127] br[127] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_128 bl[128] br[128] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_129 bl[129] br[129] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_130 bl[130] br[130] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_131 bl[131] br[131] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_132 bl[132] br[132] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_133 bl[133] br[133] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_134 bl[134] br[134] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_135 bl[135] br[135] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_136 bl[136] br[136] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_137 bl[137] br[137] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_138 bl[138] br[138] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_139 bl[139] br[139] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_140 bl[140] br[140] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_141 bl[141] br[141] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_142 bl[142] br[142] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_143 bl[143] br[143] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_144 bl[144] br[144] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_145 bl[145] br[145] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_146 bl[146] br[146] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_147 bl[147] br[147] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_148 bl[148] br[148] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_149 bl[149] br[149] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_150 bl[150] br[150] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_151 bl[151] br[151] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_152 bl[152] br[152] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_153 bl[153] br[153] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_154 bl[154] br[154] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_155 bl[155] br[155] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_156 bl[156] br[156] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_157 bl[157] br[157] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_158 bl[158] br[158] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_159 bl[159] br[159] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_160 bl[160] br[160] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_161 bl[161] br[161] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_162 bl[162] br[162] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_163 bl[163] br[163] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_164 bl[164] br[164] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_165 bl[165] br[165] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_166 bl[166] br[166] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_167 bl[167] br[167] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_168 bl[168] br[168] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_169 bl[169] br[169] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_170 bl[170] br[170] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_171 bl[171] br[171] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_172 bl[172] br[172] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_173 bl[173] br[173] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_174 bl[174] br[174] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_175 bl[175] br[175] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_176 bl[176] br[176] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_177 bl[177] br[177] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_178 bl[178] br[178] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_179 bl[179] br[179] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_180 bl[180] br[180] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_181 bl[181] br[181] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_182 bl[182] br[182] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_183 bl[183] br[183] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_184 bl[184] br[184] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_185 bl[185] br[185] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_186 bl[186] br[186] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_187 bl[187] br[187] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_188 bl[188] br[188] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_189 bl[189] br[189] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_190 bl[190] br[190] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_191 bl[191] br[191] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_192 bl[192] br[192] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_193 bl[193] br[193] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_194 bl[194] br[194] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_195 bl[195] br[195] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_196 bl[196] br[196] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_197 bl[197] br[197] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_198 bl[198] br[198] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_199 bl[199] br[199] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_200 bl[200] br[200] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_201 bl[201] br[201] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_202 bl[202] br[202] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_203 bl[203] br[203] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_204 bl[204] br[204] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_205 bl[205] br[205] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_206 bl[206] br[206] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_207 bl[207] br[207] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_208 bl[208] br[208] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_209 bl[209] br[209] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_210 bl[210] br[210] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_211 bl[211] br[211] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_212 bl[212] br[212] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_213 bl[213] br[213] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_214 bl[214] br[214] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_215 bl[215] br[215] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_216 bl[216] br[216] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_217 bl[217] br[217] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_218 bl[218] br[218] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_219 bl[219] br[219] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_220 bl[220] br[220] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_221 bl[221] br[221] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_222 bl[222] br[222] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_223 bl[223] br[223] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_224 bl[224] br[224] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_225 bl[225] br[225] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_226 bl[226] br[226] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_227 bl[227] br[227] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_228 bl[228] br[228] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_229 bl[229] br[229] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_230 bl[230] br[230] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_231 bl[231] br[231] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_232 bl[232] br[232] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_233 bl[233] br[233] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_234 bl[234] br[234] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_235 bl[235] br[235] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_236 bl[236] br[236] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_237 bl[237] br[237] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_238 bl[238] br[238] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_239 bl[239] br[239] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_240 bl[240] br[240] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_241 bl[241] br[241] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_242 bl[242] br[242] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_243 bl[243] br[243] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_244 bl[244] br[244] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_245 bl[245] br[245] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_246 bl[246] br[246] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_247 bl[247] br[247] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_248 bl[248] br[248] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_249 bl[249] br[249] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_250 bl[250] br[250] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_251 bl[251] br[251] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_252 bl[252] br[252] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_253 bl[253] br[253] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_254 bl[254] br[254] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_255 bl[255] br[255] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_256 bl[256] br[256] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_257 bl[257] br[257] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_258 bl[258] br[258] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_259 bl[259] br[259] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_260 bl[260] br[260] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_261 bl[261] br[261] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_262 bl[262] br[262] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_263 bl[263] br[263] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_264 bl[264] br[264] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_265 bl[265] br[265] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_266 bl[266] br[266] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_267 bl[267] br[267] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_268 bl[268] br[268] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_269 bl[269] br[269] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_270 bl[270] br[270] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_271 bl[271] br[271] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_272 bl[272] br[272] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_273 bl[273] br[273] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_274 bl[274] br[274] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_275 bl[275] br[275] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_276 bl[276] br[276] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_277 bl[277] br[277] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_278 bl[278] br[278] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_279 bl[279] br[279] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_280 bl[280] br[280] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_281 bl[281] br[281] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_282 bl[282] br[282] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_283 bl[283] br[283] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_284 bl[284] br[284] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_285 bl[285] br[285] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_286 bl[286] br[286] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_287 bl[287] br[287] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_288 bl[288] br[288] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_289 bl[289] br[289] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_290 bl[290] br[290] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_291 bl[291] br[291] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_292 bl[292] br[292] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_293 bl[293] br[293] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_294 bl[294] br[294] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_295 bl[295] br[295] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_296 bl[296] br[296] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_297 bl[297] br[297] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_298 bl[298] br[298] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_299 bl[299] br[299] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_300 bl[300] br[300] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_301 bl[301] br[301] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_302 bl[302] br[302] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_303 bl[303] br[303] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_304 bl[304] br[304] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_305 bl[305] br[305] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_306 bl[306] br[306] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_307 bl[307] br[307] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_308 bl[308] br[308] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_309 bl[309] br[309] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_310 bl[310] br[310] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_311 bl[311] br[311] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_312 bl[312] br[312] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_313 bl[313] br[313] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_314 bl[314] br[314] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_315 bl[315] br[315] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_316 bl[316] br[316] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_317 bl[317] br[317] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_318 bl[318] br[318] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_319 bl[319] br[319] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_320 bl[320] br[320] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_321 bl[321] br[321] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_322 bl[322] br[322] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_323 bl[323] br[323] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_324 bl[324] br[324] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_325 bl[325] br[325] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_326 bl[326] br[326] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_327 bl[327] br[327] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_328 bl[328] br[328] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_329 bl[329] br[329] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_330 bl[330] br[330] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_331 bl[331] br[331] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_332 bl[332] br[332] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_333 bl[333] br[333] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_334 bl[334] br[334] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_335 bl[335] br[335] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_336 bl[336] br[336] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_337 bl[337] br[337] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_338 bl[338] br[338] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_339 bl[339] br[339] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_340 bl[340] br[340] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_341 bl[341] br[341] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_342 bl[342] br[342] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_343 bl[343] br[343] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_344 bl[344] br[344] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_345 bl[345] br[345] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_346 bl[346] br[346] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_347 bl[347] br[347] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_348 bl[348] br[348] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_349 bl[349] br[349] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_350 bl[350] br[350] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_351 bl[351] br[351] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_352 bl[352] br[352] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_353 bl[353] br[353] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_354 bl[354] br[354] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_355 bl[355] br[355] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_356 bl[356] br[356] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_357 bl[357] br[357] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_358 bl[358] br[358] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_359 bl[359] br[359] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_360 bl[360] br[360] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_361 bl[361] br[361] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_362 bl[362] br[362] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_363 bl[363] br[363] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_364 bl[364] br[364] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_365 bl[365] br[365] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_366 bl[366] br[366] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_367 bl[367] br[367] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_368 bl[368] br[368] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_369 bl[369] br[369] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_370 bl[370] br[370] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_371 bl[371] br[371] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_372 bl[372] br[372] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_373 bl[373] br[373] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_374 bl[374] br[374] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_375 bl[375] br[375] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_376 bl[376] br[376] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_377 bl[377] br[377] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_378 bl[378] br[378] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_379 bl[379] br[379] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_380 bl[380] br[380] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_381 bl[381] br[381] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_382 bl[382] br[382] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_383 bl[383] br[383] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_384 bl[384] br[384] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_385 bl[385] br[385] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_386 bl[386] br[386] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_387 bl[387] br[387] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_388 bl[388] br[388] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_389 bl[389] br[389] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_390 bl[390] br[390] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_391 bl[391] br[391] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_392 bl[392] br[392] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_393 bl[393] br[393] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_394 bl[394] br[394] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_395 bl[395] br[395] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_396 bl[396] br[396] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_397 bl[397] br[397] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_398 bl[398] br[398] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_399 bl[399] br[399] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_400 bl[400] br[400] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_401 bl[401] br[401] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_402 bl[402] br[402] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_403 bl[403] br[403] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_404 bl[404] br[404] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_405 bl[405] br[405] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_406 bl[406] br[406] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_407 bl[407] br[407] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_408 bl[408] br[408] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_409 bl[409] br[409] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_410 bl[410] br[410] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_411 bl[411] br[411] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_412 bl[412] br[412] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_413 bl[413] br[413] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_414 bl[414] br[414] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_415 bl[415] br[415] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_416 bl[416] br[416] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_417 bl[417] br[417] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_418 bl[418] br[418] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_419 bl[419] br[419] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_420 bl[420] br[420] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_421 bl[421] br[421] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_422 bl[422] br[422] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_423 bl[423] br[423] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_424 bl[424] br[424] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_425 bl[425] br[425] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_426 bl[426] br[426] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_427 bl[427] br[427] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_428 bl[428] br[428] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_429 bl[429] br[429] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_430 bl[430] br[430] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_431 bl[431] br[431] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_432 bl[432] br[432] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_433 bl[433] br[433] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_434 bl[434] br[434] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_435 bl[435] br[435] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_436 bl[436] br[436] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_437 bl[437] br[437] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_438 bl[438] br[438] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_439 bl[439] br[439] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_440 bl[440] br[440] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_441 bl[441] br[441] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_442 bl[442] br[442] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_443 bl[443] br[443] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_444 bl[444] br[444] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_445 bl[445] br[445] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_446 bl[446] br[446] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_447 bl[447] br[447] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_448 bl[448] br[448] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_449 bl[449] br[449] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_450 bl[450] br[450] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_451 bl[451] br[451] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_452 bl[452] br[452] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_453 bl[453] br[453] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_454 bl[454] br[454] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_455 bl[455] br[455] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_456 bl[456] br[456] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_457 bl[457] br[457] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_458 bl[458] br[458] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_459 bl[459] br[459] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_460 bl[460] br[460] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_461 bl[461] br[461] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_462 bl[462] br[462] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_463 bl[463] br[463] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_464 bl[464] br[464] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_465 bl[465] br[465] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_466 bl[466] br[466] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_467 bl[467] br[467] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_468 bl[468] br[468] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_469 bl[469] br[469] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_470 bl[470] br[470] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_471 bl[471] br[471] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_472 bl[472] br[472] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_473 bl[473] br[473] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_474 bl[474] br[474] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_475 bl[475] br[475] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_476 bl[476] br[476] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_477 bl[477] br[477] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_478 bl[478] br[478] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_479 bl[479] br[479] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_480 bl[480] br[480] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_481 bl[481] br[481] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_482 bl[482] br[482] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_483 bl[483] br[483] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_484 bl[484] br[484] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_485 bl[485] br[485] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_486 bl[486] br[486] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_487 bl[487] br[487] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_488 bl[488] br[488] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_489 bl[489] br[489] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_490 bl[490] br[490] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_491 bl[491] br[491] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_492 bl[492] br[492] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_493 bl[493] br[493] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_494 bl[494] br[494] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_495 bl[495] br[495] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_496 bl[496] br[496] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_497 bl[497] br[497] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_498 bl[498] br[498] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_499 bl[499] br[499] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_500 bl[500] br[500] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_501 bl[501] br[501] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_502 bl[502] br[502] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_503 bl[503] br[503] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_504 bl[504] br[504] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_505 bl[505] br[505] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_506 bl[506] br[506] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_507 bl[507] br[507] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_508 bl[508] br[508] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_509 bl[509] br[509] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_510 bl[510] br[510] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_11_511 bl[511] br[511] vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xcell_12_0 bl[0] br[0] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_1 bl[1] br[1] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_2 bl[2] br[2] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_3 bl[3] br[3] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_4 bl[4] br[4] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_5 bl[5] br[5] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_6 bl[6] br[6] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_7 bl[7] br[7] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_8 bl[8] br[8] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_9 bl[9] br[9] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_10 bl[10] br[10] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_11 bl[11] br[11] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_12 bl[12] br[12] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_13 bl[13] br[13] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_14 bl[14] br[14] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_15 bl[15] br[15] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_16 bl[16] br[16] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_17 bl[17] br[17] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_18 bl[18] br[18] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_19 bl[19] br[19] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_20 bl[20] br[20] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_21 bl[21] br[21] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_22 bl[22] br[22] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_23 bl[23] br[23] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_24 bl[24] br[24] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_25 bl[25] br[25] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_26 bl[26] br[26] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_27 bl[27] br[27] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_28 bl[28] br[28] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_29 bl[29] br[29] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_30 bl[30] br[30] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_31 bl[31] br[31] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_32 bl[32] br[32] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_33 bl[33] br[33] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_34 bl[34] br[34] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_35 bl[35] br[35] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_36 bl[36] br[36] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_37 bl[37] br[37] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_38 bl[38] br[38] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_39 bl[39] br[39] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_40 bl[40] br[40] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_41 bl[41] br[41] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_42 bl[42] br[42] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_43 bl[43] br[43] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_44 bl[44] br[44] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_45 bl[45] br[45] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_46 bl[46] br[46] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_47 bl[47] br[47] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_48 bl[48] br[48] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_49 bl[49] br[49] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_50 bl[50] br[50] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_51 bl[51] br[51] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_52 bl[52] br[52] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_53 bl[53] br[53] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_54 bl[54] br[54] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_55 bl[55] br[55] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_56 bl[56] br[56] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_57 bl[57] br[57] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_58 bl[58] br[58] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_59 bl[59] br[59] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_60 bl[60] br[60] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_61 bl[61] br[61] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_62 bl[62] br[62] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_63 bl[63] br[63] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_64 bl[64] br[64] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_65 bl[65] br[65] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_66 bl[66] br[66] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_67 bl[67] br[67] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_68 bl[68] br[68] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_69 bl[69] br[69] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_70 bl[70] br[70] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_71 bl[71] br[71] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_72 bl[72] br[72] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_73 bl[73] br[73] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_74 bl[74] br[74] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_75 bl[75] br[75] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_76 bl[76] br[76] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_77 bl[77] br[77] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_78 bl[78] br[78] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_79 bl[79] br[79] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_80 bl[80] br[80] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_81 bl[81] br[81] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_82 bl[82] br[82] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_83 bl[83] br[83] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_84 bl[84] br[84] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_85 bl[85] br[85] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_86 bl[86] br[86] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_87 bl[87] br[87] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_88 bl[88] br[88] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_89 bl[89] br[89] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_90 bl[90] br[90] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_91 bl[91] br[91] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_92 bl[92] br[92] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_93 bl[93] br[93] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_94 bl[94] br[94] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_95 bl[95] br[95] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_96 bl[96] br[96] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_97 bl[97] br[97] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_98 bl[98] br[98] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_99 bl[99] br[99] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_100 bl[100] br[100] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_101 bl[101] br[101] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_102 bl[102] br[102] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_103 bl[103] br[103] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_104 bl[104] br[104] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_105 bl[105] br[105] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_106 bl[106] br[106] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_107 bl[107] br[107] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_108 bl[108] br[108] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_109 bl[109] br[109] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_110 bl[110] br[110] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_111 bl[111] br[111] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_112 bl[112] br[112] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_113 bl[113] br[113] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_114 bl[114] br[114] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_115 bl[115] br[115] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_116 bl[116] br[116] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_117 bl[117] br[117] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_118 bl[118] br[118] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_119 bl[119] br[119] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_120 bl[120] br[120] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_121 bl[121] br[121] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_122 bl[122] br[122] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_123 bl[123] br[123] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_124 bl[124] br[124] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_125 bl[125] br[125] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_126 bl[126] br[126] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_127 bl[127] br[127] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_128 bl[128] br[128] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_129 bl[129] br[129] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_130 bl[130] br[130] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_131 bl[131] br[131] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_132 bl[132] br[132] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_133 bl[133] br[133] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_134 bl[134] br[134] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_135 bl[135] br[135] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_136 bl[136] br[136] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_137 bl[137] br[137] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_138 bl[138] br[138] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_139 bl[139] br[139] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_140 bl[140] br[140] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_141 bl[141] br[141] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_142 bl[142] br[142] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_143 bl[143] br[143] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_144 bl[144] br[144] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_145 bl[145] br[145] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_146 bl[146] br[146] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_147 bl[147] br[147] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_148 bl[148] br[148] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_149 bl[149] br[149] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_150 bl[150] br[150] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_151 bl[151] br[151] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_152 bl[152] br[152] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_153 bl[153] br[153] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_154 bl[154] br[154] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_155 bl[155] br[155] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_156 bl[156] br[156] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_157 bl[157] br[157] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_158 bl[158] br[158] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_159 bl[159] br[159] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_160 bl[160] br[160] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_161 bl[161] br[161] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_162 bl[162] br[162] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_163 bl[163] br[163] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_164 bl[164] br[164] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_165 bl[165] br[165] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_166 bl[166] br[166] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_167 bl[167] br[167] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_168 bl[168] br[168] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_169 bl[169] br[169] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_170 bl[170] br[170] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_171 bl[171] br[171] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_172 bl[172] br[172] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_173 bl[173] br[173] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_174 bl[174] br[174] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_175 bl[175] br[175] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_176 bl[176] br[176] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_177 bl[177] br[177] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_178 bl[178] br[178] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_179 bl[179] br[179] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_180 bl[180] br[180] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_181 bl[181] br[181] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_182 bl[182] br[182] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_183 bl[183] br[183] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_184 bl[184] br[184] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_185 bl[185] br[185] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_186 bl[186] br[186] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_187 bl[187] br[187] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_188 bl[188] br[188] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_189 bl[189] br[189] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_190 bl[190] br[190] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_191 bl[191] br[191] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_192 bl[192] br[192] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_193 bl[193] br[193] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_194 bl[194] br[194] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_195 bl[195] br[195] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_196 bl[196] br[196] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_197 bl[197] br[197] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_198 bl[198] br[198] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_199 bl[199] br[199] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_200 bl[200] br[200] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_201 bl[201] br[201] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_202 bl[202] br[202] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_203 bl[203] br[203] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_204 bl[204] br[204] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_205 bl[205] br[205] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_206 bl[206] br[206] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_207 bl[207] br[207] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_208 bl[208] br[208] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_209 bl[209] br[209] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_210 bl[210] br[210] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_211 bl[211] br[211] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_212 bl[212] br[212] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_213 bl[213] br[213] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_214 bl[214] br[214] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_215 bl[215] br[215] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_216 bl[216] br[216] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_217 bl[217] br[217] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_218 bl[218] br[218] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_219 bl[219] br[219] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_220 bl[220] br[220] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_221 bl[221] br[221] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_222 bl[222] br[222] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_223 bl[223] br[223] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_224 bl[224] br[224] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_225 bl[225] br[225] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_226 bl[226] br[226] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_227 bl[227] br[227] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_228 bl[228] br[228] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_229 bl[229] br[229] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_230 bl[230] br[230] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_231 bl[231] br[231] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_232 bl[232] br[232] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_233 bl[233] br[233] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_234 bl[234] br[234] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_235 bl[235] br[235] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_236 bl[236] br[236] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_237 bl[237] br[237] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_238 bl[238] br[238] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_239 bl[239] br[239] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_240 bl[240] br[240] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_241 bl[241] br[241] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_242 bl[242] br[242] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_243 bl[243] br[243] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_244 bl[244] br[244] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_245 bl[245] br[245] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_246 bl[246] br[246] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_247 bl[247] br[247] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_248 bl[248] br[248] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_249 bl[249] br[249] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_250 bl[250] br[250] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_251 bl[251] br[251] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_252 bl[252] br[252] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_253 bl[253] br[253] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_254 bl[254] br[254] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_255 bl[255] br[255] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_256 bl[256] br[256] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_257 bl[257] br[257] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_258 bl[258] br[258] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_259 bl[259] br[259] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_260 bl[260] br[260] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_261 bl[261] br[261] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_262 bl[262] br[262] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_263 bl[263] br[263] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_264 bl[264] br[264] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_265 bl[265] br[265] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_266 bl[266] br[266] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_267 bl[267] br[267] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_268 bl[268] br[268] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_269 bl[269] br[269] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_270 bl[270] br[270] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_271 bl[271] br[271] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_272 bl[272] br[272] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_273 bl[273] br[273] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_274 bl[274] br[274] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_275 bl[275] br[275] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_276 bl[276] br[276] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_277 bl[277] br[277] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_278 bl[278] br[278] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_279 bl[279] br[279] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_280 bl[280] br[280] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_281 bl[281] br[281] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_282 bl[282] br[282] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_283 bl[283] br[283] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_284 bl[284] br[284] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_285 bl[285] br[285] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_286 bl[286] br[286] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_287 bl[287] br[287] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_288 bl[288] br[288] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_289 bl[289] br[289] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_290 bl[290] br[290] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_291 bl[291] br[291] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_292 bl[292] br[292] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_293 bl[293] br[293] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_294 bl[294] br[294] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_295 bl[295] br[295] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_296 bl[296] br[296] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_297 bl[297] br[297] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_298 bl[298] br[298] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_299 bl[299] br[299] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_300 bl[300] br[300] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_301 bl[301] br[301] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_302 bl[302] br[302] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_303 bl[303] br[303] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_304 bl[304] br[304] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_305 bl[305] br[305] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_306 bl[306] br[306] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_307 bl[307] br[307] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_308 bl[308] br[308] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_309 bl[309] br[309] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_310 bl[310] br[310] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_311 bl[311] br[311] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_312 bl[312] br[312] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_313 bl[313] br[313] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_314 bl[314] br[314] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_315 bl[315] br[315] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_316 bl[316] br[316] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_317 bl[317] br[317] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_318 bl[318] br[318] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_319 bl[319] br[319] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_320 bl[320] br[320] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_321 bl[321] br[321] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_322 bl[322] br[322] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_323 bl[323] br[323] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_324 bl[324] br[324] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_325 bl[325] br[325] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_326 bl[326] br[326] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_327 bl[327] br[327] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_328 bl[328] br[328] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_329 bl[329] br[329] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_330 bl[330] br[330] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_331 bl[331] br[331] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_332 bl[332] br[332] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_333 bl[333] br[333] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_334 bl[334] br[334] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_335 bl[335] br[335] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_336 bl[336] br[336] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_337 bl[337] br[337] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_338 bl[338] br[338] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_339 bl[339] br[339] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_340 bl[340] br[340] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_341 bl[341] br[341] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_342 bl[342] br[342] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_343 bl[343] br[343] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_344 bl[344] br[344] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_345 bl[345] br[345] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_346 bl[346] br[346] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_347 bl[347] br[347] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_348 bl[348] br[348] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_349 bl[349] br[349] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_350 bl[350] br[350] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_351 bl[351] br[351] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_352 bl[352] br[352] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_353 bl[353] br[353] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_354 bl[354] br[354] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_355 bl[355] br[355] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_356 bl[356] br[356] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_357 bl[357] br[357] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_358 bl[358] br[358] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_359 bl[359] br[359] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_360 bl[360] br[360] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_361 bl[361] br[361] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_362 bl[362] br[362] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_363 bl[363] br[363] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_364 bl[364] br[364] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_365 bl[365] br[365] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_366 bl[366] br[366] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_367 bl[367] br[367] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_368 bl[368] br[368] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_369 bl[369] br[369] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_370 bl[370] br[370] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_371 bl[371] br[371] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_372 bl[372] br[372] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_373 bl[373] br[373] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_374 bl[374] br[374] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_375 bl[375] br[375] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_376 bl[376] br[376] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_377 bl[377] br[377] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_378 bl[378] br[378] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_379 bl[379] br[379] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_380 bl[380] br[380] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_381 bl[381] br[381] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_382 bl[382] br[382] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_383 bl[383] br[383] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_384 bl[384] br[384] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_385 bl[385] br[385] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_386 bl[386] br[386] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_387 bl[387] br[387] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_388 bl[388] br[388] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_389 bl[389] br[389] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_390 bl[390] br[390] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_391 bl[391] br[391] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_392 bl[392] br[392] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_393 bl[393] br[393] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_394 bl[394] br[394] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_395 bl[395] br[395] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_396 bl[396] br[396] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_397 bl[397] br[397] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_398 bl[398] br[398] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_399 bl[399] br[399] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_400 bl[400] br[400] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_401 bl[401] br[401] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_402 bl[402] br[402] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_403 bl[403] br[403] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_404 bl[404] br[404] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_405 bl[405] br[405] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_406 bl[406] br[406] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_407 bl[407] br[407] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_408 bl[408] br[408] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_409 bl[409] br[409] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_410 bl[410] br[410] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_411 bl[411] br[411] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_412 bl[412] br[412] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_413 bl[413] br[413] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_414 bl[414] br[414] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_415 bl[415] br[415] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_416 bl[416] br[416] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_417 bl[417] br[417] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_418 bl[418] br[418] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_419 bl[419] br[419] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_420 bl[420] br[420] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_421 bl[421] br[421] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_422 bl[422] br[422] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_423 bl[423] br[423] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_424 bl[424] br[424] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_425 bl[425] br[425] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_426 bl[426] br[426] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_427 bl[427] br[427] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_428 bl[428] br[428] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_429 bl[429] br[429] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_430 bl[430] br[430] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_431 bl[431] br[431] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_432 bl[432] br[432] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_433 bl[433] br[433] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_434 bl[434] br[434] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_435 bl[435] br[435] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_436 bl[436] br[436] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_437 bl[437] br[437] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_438 bl[438] br[438] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_439 bl[439] br[439] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_440 bl[440] br[440] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_441 bl[441] br[441] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_442 bl[442] br[442] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_443 bl[443] br[443] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_444 bl[444] br[444] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_445 bl[445] br[445] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_446 bl[446] br[446] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_447 bl[447] br[447] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_448 bl[448] br[448] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_449 bl[449] br[449] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_450 bl[450] br[450] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_451 bl[451] br[451] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_452 bl[452] br[452] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_453 bl[453] br[453] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_454 bl[454] br[454] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_455 bl[455] br[455] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_456 bl[456] br[456] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_457 bl[457] br[457] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_458 bl[458] br[458] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_459 bl[459] br[459] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_460 bl[460] br[460] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_461 bl[461] br[461] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_462 bl[462] br[462] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_463 bl[463] br[463] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_464 bl[464] br[464] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_465 bl[465] br[465] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_466 bl[466] br[466] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_467 bl[467] br[467] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_468 bl[468] br[468] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_469 bl[469] br[469] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_470 bl[470] br[470] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_471 bl[471] br[471] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_472 bl[472] br[472] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_473 bl[473] br[473] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_474 bl[474] br[474] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_475 bl[475] br[475] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_476 bl[476] br[476] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_477 bl[477] br[477] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_478 bl[478] br[478] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_479 bl[479] br[479] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_480 bl[480] br[480] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_481 bl[481] br[481] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_482 bl[482] br[482] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_483 bl[483] br[483] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_484 bl[484] br[484] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_485 bl[485] br[485] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_486 bl[486] br[486] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_487 bl[487] br[487] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_488 bl[488] br[488] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_489 bl[489] br[489] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_490 bl[490] br[490] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_491 bl[491] br[491] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_492 bl[492] br[492] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_493 bl[493] br[493] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_494 bl[494] br[494] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_495 bl[495] br[495] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_496 bl[496] br[496] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_497 bl[497] br[497] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_498 bl[498] br[498] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_499 bl[499] br[499] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_500 bl[500] br[500] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_501 bl[501] br[501] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_502 bl[502] br[502] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_503 bl[503] br[503] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_504 bl[504] br[504] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_505 bl[505] br[505] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_506 bl[506] br[506] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_507 bl[507] br[507] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_508 bl[508] br[508] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_509 bl[509] br[509] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_510 bl[510] br[510] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_12_511 bl[511] br[511] vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xcell_13_0 bl[0] br[0] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_1 bl[1] br[1] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_2 bl[2] br[2] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_3 bl[3] br[3] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_4 bl[4] br[4] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_5 bl[5] br[5] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_6 bl[6] br[6] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_7 bl[7] br[7] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_8 bl[8] br[8] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_9 bl[9] br[9] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_10 bl[10] br[10] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_11 bl[11] br[11] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_12 bl[12] br[12] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_13 bl[13] br[13] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_14 bl[14] br[14] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_15 bl[15] br[15] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_16 bl[16] br[16] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_17 bl[17] br[17] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_18 bl[18] br[18] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_19 bl[19] br[19] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_20 bl[20] br[20] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_21 bl[21] br[21] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_22 bl[22] br[22] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_23 bl[23] br[23] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_24 bl[24] br[24] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_25 bl[25] br[25] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_26 bl[26] br[26] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_27 bl[27] br[27] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_28 bl[28] br[28] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_29 bl[29] br[29] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_30 bl[30] br[30] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_31 bl[31] br[31] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_32 bl[32] br[32] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_33 bl[33] br[33] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_34 bl[34] br[34] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_35 bl[35] br[35] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_36 bl[36] br[36] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_37 bl[37] br[37] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_38 bl[38] br[38] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_39 bl[39] br[39] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_40 bl[40] br[40] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_41 bl[41] br[41] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_42 bl[42] br[42] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_43 bl[43] br[43] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_44 bl[44] br[44] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_45 bl[45] br[45] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_46 bl[46] br[46] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_47 bl[47] br[47] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_48 bl[48] br[48] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_49 bl[49] br[49] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_50 bl[50] br[50] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_51 bl[51] br[51] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_52 bl[52] br[52] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_53 bl[53] br[53] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_54 bl[54] br[54] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_55 bl[55] br[55] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_56 bl[56] br[56] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_57 bl[57] br[57] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_58 bl[58] br[58] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_59 bl[59] br[59] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_60 bl[60] br[60] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_61 bl[61] br[61] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_62 bl[62] br[62] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_63 bl[63] br[63] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_64 bl[64] br[64] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_65 bl[65] br[65] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_66 bl[66] br[66] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_67 bl[67] br[67] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_68 bl[68] br[68] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_69 bl[69] br[69] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_70 bl[70] br[70] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_71 bl[71] br[71] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_72 bl[72] br[72] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_73 bl[73] br[73] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_74 bl[74] br[74] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_75 bl[75] br[75] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_76 bl[76] br[76] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_77 bl[77] br[77] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_78 bl[78] br[78] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_79 bl[79] br[79] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_80 bl[80] br[80] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_81 bl[81] br[81] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_82 bl[82] br[82] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_83 bl[83] br[83] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_84 bl[84] br[84] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_85 bl[85] br[85] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_86 bl[86] br[86] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_87 bl[87] br[87] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_88 bl[88] br[88] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_89 bl[89] br[89] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_90 bl[90] br[90] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_91 bl[91] br[91] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_92 bl[92] br[92] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_93 bl[93] br[93] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_94 bl[94] br[94] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_95 bl[95] br[95] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_96 bl[96] br[96] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_97 bl[97] br[97] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_98 bl[98] br[98] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_99 bl[99] br[99] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_100 bl[100] br[100] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_101 bl[101] br[101] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_102 bl[102] br[102] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_103 bl[103] br[103] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_104 bl[104] br[104] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_105 bl[105] br[105] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_106 bl[106] br[106] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_107 bl[107] br[107] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_108 bl[108] br[108] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_109 bl[109] br[109] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_110 bl[110] br[110] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_111 bl[111] br[111] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_112 bl[112] br[112] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_113 bl[113] br[113] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_114 bl[114] br[114] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_115 bl[115] br[115] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_116 bl[116] br[116] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_117 bl[117] br[117] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_118 bl[118] br[118] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_119 bl[119] br[119] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_120 bl[120] br[120] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_121 bl[121] br[121] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_122 bl[122] br[122] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_123 bl[123] br[123] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_124 bl[124] br[124] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_125 bl[125] br[125] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_126 bl[126] br[126] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_127 bl[127] br[127] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_128 bl[128] br[128] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_129 bl[129] br[129] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_130 bl[130] br[130] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_131 bl[131] br[131] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_132 bl[132] br[132] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_133 bl[133] br[133] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_134 bl[134] br[134] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_135 bl[135] br[135] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_136 bl[136] br[136] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_137 bl[137] br[137] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_138 bl[138] br[138] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_139 bl[139] br[139] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_140 bl[140] br[140] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_141 bl[141] br[141] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_142 bl[142] br[142] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_143 bl[143] br[143] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_144 bl[144] br[144] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_145 bl[145] br[145] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_146 bl[146] br[146] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_147 bl[147] br[147] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_148 bl[148] br[148] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_149 bl[149] br[149] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_150 bl[150] br[150] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_151 bl[151] br[151] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_152 bl[152] br[152] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_153 bl[153] br[153] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_154 bl[154] br[154] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_155 bl[155] br[155] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_156 bl[156] br[156] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_157 bl[157] br[157] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_158 bl[158] br[158] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_159 bl[159] br[159] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_160 bl[160] br[160] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_161 bl[161] br[161] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_162 bl[162] br[162] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_163 bl[163] br[163] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_164 bl[164] br[164] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_165 bl[165] br[165] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_166 bl[166] br[166] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_167 bl[167] br[167] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_168 bl[168] br[168] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_169 bl[169] br[169] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_170 bl[170] br[170] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_171 bl[171] br[171] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_172 bl[172] br[172] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_173 bl[173] br[173] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_174 bl[174] br[174] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_175 bl[175] br[175] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_176 bl[176] br[176] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_177 bl[177] br[177] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_178 bl[178] br[178] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_179 bl[179] br[179] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_180 bl[180] br[180] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_181 bl[181] br[181] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_182 bl[182] br[182] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_183 bl[183] br[183] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_184 bl[184] br[184] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_185 bl[185] br[185] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_186 bl[186] br[186] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_187 bl[187] br[187] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_188 bl[188] br[188] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_189 bl[189] br[189] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_190 bl[190] br[190] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_191 bl[191] br[191] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_192 bl[192] br[192] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_193 bl[193] br[193] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_194 bl[194] br[194] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_195 bl[195] br[195] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_196 bl[196] br[196] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_197 bl[197] br[197] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_198 bl[198] br[198] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_199 bl[199] br[199] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_200 bl[200] br[200] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_201 bl[201] br[201] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_202 bl[202] br[202] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_203 bl[203] br[203] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_204 bl[204] br[204] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_205 bl[205] br[205] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_206 bl[206] br[206] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_207 bl[207] br[207] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_208 bl[208] br[208] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_209 bl[209] br[209] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_210 bl[210] br[210] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_211 bl[211] br[211] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_212 bl[212] br[212] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_213 bl[213] br[213] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_214 bl[214] br[214] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_215 bl[215] br[215] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_216 bl[216] br[216] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_217 bl[217] br[217] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_218 bl[218] br[218] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_219 bl[219] br[219] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_220 bl[220] br[220] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_221 bl[221] br[221] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_222 bl[222] br[222] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_223 bl[223] br[223] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_224 bl[224] br[224] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_225 bl[225] br[225] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_226 bl[226] br[226] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_227 bl[227] br[227] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_228 bl[228] br[228] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_229 bl[229] br[229] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_230 bl[230] br[230] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_231 bl[231] br[231] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_232 bl[232] br[232] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_233 bl[233] br[233] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_234 bl[234] br[234] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_235 bl[235] br[235] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_236 bl[236] br[236] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_237 bl[237] br[237] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_238 bl[238] br[238] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_239 bl[239] br[239] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_240 bl[240] br[240] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_241 bl[241] br[241] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_242 bl[242] br[242] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_243 bl[243] br[243] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_244 bl[244] br[244] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_245 bl[245] br[245] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_246 bl[246] br[246] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_247 bl[247] br[247] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_248 bl[248] br[248] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_249 bl[249] br[249] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_250 bl[250] br[250] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_251 bl[251] br[251] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_252 bl[252] br[252] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_253 bl[253] br[253] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_254 bl[254] br[254] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_255 bl[255] br[255] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_256 bl[256] br[256] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_257 bl[257] br[257] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_258 bl[258] br[258] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_259 bl[259] br[259] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_260 bl[260] br[260] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_261 bl[261] br[261] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_262 bl[262] br[262] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_263 bl[263] br[263] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_264 bl[264] br[264] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_265 bl[265] br[265] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_266 bl[266] br[266] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_267 bl[267] br[267] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_268 bl[268] br[268] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_269 bl[269] br[269] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_270 bl[270] br[270] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_271 bl[271] br[271] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_272 bl[272] br[272] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_273 bl[273] br[273] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_274 bl[274] br[274] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_275 bl[275] br[275] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_276 bl[276] br[276] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_277 bl[277] br[277] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_278 bl[278] br[278] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_279 bl[279] br[279] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_280 bl[280] br[280] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_281 bl[281] br[281] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_282 bl[282] br[282] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_283 bl[283] br[283] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_284 bl[284] br[284] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_285 bl[285] br[285] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_286 bl[286] br[286] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_287 bl[287] br[287] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_288 bl[288] br[288] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_289 bl[289] br[289] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_290 bl[290] br[290] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_291 bl[291] br[291] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_292 bl[292] br[292] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_293 bl[293] br[293] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_294 bl[294] br[294] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_295 bl[295] br[295] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_296 bl[296] br[296] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_297 bl[297] br[297] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_298 bl[298] br[298] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_299 bl[299] br[299] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_300 bl[300] br[300] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_301 bl[301] br[301] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_302 bl[302] br[302] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_303 bl[303] br[303] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_304 bl[304] br[304] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_305 bl[305] br[305] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_306 bl[306] br[306] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_307 bl[307] br[307] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_308 bl[308] br[308] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_309 bl[309] br[309] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_310 bl[310] br[310] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_311 bl[311] br[311] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_312 bl[312] br[312] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_313 bl[313] br[313] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_314 bl[314] br[314] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_315 bl[315] br[315] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_316 bl[316] br[316] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_317 bl[317] br[317] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_318 bl[318] br[318] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_319 bl[319] br[319] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_320 bl[320] br[320] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_321 bl[321] br[321] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_322 bl[322] br[322] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_323 bl[323] br[323] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_324 bl[324] br[324] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_325 bl[325] br[325] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_326 bl[326] br[326] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_327 bl[327] br[327] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_328 bl[328] br[328] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_329 bl[329] br[329] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_330 bl[330] br[330] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_331 bl[331] br[331] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_332 bl[332] br[332] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_333 bl[333] br[333] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_334 bl[334] br[334] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_335 bl[335] br[335] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_336 bl[336] br[336] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_337 bl[337] br[337] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_338 bl[338] br[338] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_339 bl[339] br[339] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_340 bl[340] br[340] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_341 bl[341] br[341] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_342 bl[342] br[342] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_343 bl[343] br[343] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_344 bl[344] br[344] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_345 bl[345] br[345] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_346 bl[346] br[346] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_347 bl[347] br[347] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_348 bl[348] br[348] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_349 bl[349] br[349] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_350 bl[350] br[350] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_351 bl[351] br[351] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_352 bl[352] br[352] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_353 bl[353] br[353] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_354 bl[354] br[354] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_355 bl[355] br[355] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_356 bl[356] br[356] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_357 bl[357] br[357] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_358 bl[358] br[358] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_359 bl[359] br[359] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_360 bl[360] br[360] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_361 bl[361] br[361] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_362 bl[362] br[362] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_363 bl[363] br[363] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_364 bl[364] br[364] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_365 bl[365] br[365] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_366 bl[366] br[366] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_367 bl[367] br[367] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_368 bl[368] br[368] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_369 bl[369] br[369] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_370 bl[370] br[370] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_371 bl[371] br[371] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_372 bl[372] br[372] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_373 bl[373] br[373] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_374 bl[374] br[374] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_375 bl[375] br[375] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_376 bl[376] br[376] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_377 bl[377] br[377] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_378 bl[378] br[378] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_379 bl[379] br[379] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_380 bl[380] br[380] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_381 bl[381] br[381] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_382 bl[382] br[382] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_383 bl[383] br[383] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_384 bl[384] br[384] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_385 bl[385] br[385] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_386 bl[386] br[386] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_387 bl[387] br[387] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_388 bl[388] br[388] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_389 bl[389] br[389] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_390 bl[390] br[390] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_391 bl[391] br[391] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_392 bl[392] br[392] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_393 bl[393] br[393] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_394 bl[394] br[394] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_395 bl[395] br[395] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_396 bl[396] br[396] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_397 bl[397] br[397] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_398 bl[398] br[398] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_399 bl[399] br[399] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_400 bl[400] br[400] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_401 bl[401] br[401] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_402 bl[402] br[402] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_403 bl[403] br[403] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_404 bl[404] br[404] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_405 bl[405] br[405] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_406 bl[406] br[406] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_407 bl[407] br[407] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_408 bl[408] br[408] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_409 bl[409] br[409] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_410 bl[410] br[410] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_411 bl[411] br[411] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_412 bl[412] br[412] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_413 bl[413] br[413] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_414 bl[414] br[414] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_415 bl[415] br[415] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_416 bl[416] br[416] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_417 bl[417] br[417] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_418 bl[418] br[418] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_419 bl[419] br[419] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_420 bl[420] br[420] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_421 bl[421] br[421] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_422 bl[422] br[422] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_423 bl[423] br[423] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_424 bl[424] br[424] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_425 bl[425] br[425] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_426 bl[426] br[426] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_427 bl[427] br[427] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_428 bl[428] br[428] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_429 bl[429] br[429] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_430 bl[430] br[430] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_431 bl[431] br[431] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_432 bl[432] br[432] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_433 bl[433] br[433] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_434 bl[434] br[434] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_435 bl[435] br[435] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_436 bl[436] br[436] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_437 bl[437] br[437] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_438 bl[438] br[438] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_439 bl[439] br[439] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_440 bl[440] br[440] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_441 bl[441] br[441] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_442 bl[442] br[442] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_443 bl[443] br[443] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_444 bl[444] br[444] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_445 bl[445] br[445] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_446 bl[446] br[446] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_447 bl[447] br[447] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_448 bl[448] br[448] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_449 bl[449] br[449] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_450 bl[450] br[450] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_451 bl[451] br[451] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_452 bl[452] br[452] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_453 bl[453] br[453] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_454 bl[454] br[454] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_455 bl[455] br[455] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_456 bl[456] br[456] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_457 bl[457] br[457] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_458 bl[458] br[458] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_459 bl[459] br[459] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_460 bl[460] br[460] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_461 bl[461] br[461] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_462 bl[462] br[462] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_463 bl[463] br[463] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_464 bl[464] br[464] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_465 bl[465] br[465] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_466 bl[466] br[466] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_467 bl[467] br[467] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_468 bl[468] br[468] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_469 bl[469] br[469] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_470 bl[470] br[470] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_471 bl[471] br[471] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_472 bl[472] br[472] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_473 bl[473] br[473] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_474 bl[474] br[474] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_475 bl[475] br[475] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_476 bl[476] br[476] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_477 bl[477] br[477] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_478 bl[478] br[478] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_479 bl[479] br[479] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_480 bl[480] br[480] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_481 bl[481] br[481] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_482 bl[482] br[482] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_483 bl[483] br[483] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_484 bl[484] br[484] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_485 bl[485] br[485] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_486 bl[486] br[486] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_487 bl[487] br[487] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_488 bl[488] br[488] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_489 bl[489] br[489] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_490 bl[490] br[490] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_491 bl[491] br[491] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_492 bl[492] br[492] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_493 bl[493] br[493] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_494 bl[494] br[494] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_495 bl[495] br[495] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_496 bl[496] br[496] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_497 bl[497] br[497] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_498 bl[498] br[498] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_499 bl[499] br[499] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_500 bl[500] br[500] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_501 bl[501] br[501] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_502 bl[502] br[502] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_503 bl[503] br[503] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_504 bl[504] br[504] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_505 bl[505] br[505] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_506 bl[506] br[506] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_507 bl[507] br[507] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_508 bl[508] br[508] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_509 bl[509] br[509] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_510 bl[510] br[510] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_13_511 bl[511] br[511] vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xcell_14_0 bl[0] br[0] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_1 bl[1] br[1] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_2 bl[2] br[2] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_3 bl[3] br[3] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_4 bl[4] br[4] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_5 bl[5] br[5] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_6 bl[6] br[6] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_7 bl[7] br[7] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_8 bl[8] br[8] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_9 bl[9] br[9] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_10 bl[10] br[10] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_11 bl[11] br[11] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_12 bl[12] br[12] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_13 bl[13] br[13] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_14 bl[14] br[14] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_15 bl[15] br[15] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_16 bl[16] br[16] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_17 bl[17] br[17] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_18 bl[18] br[18] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_19 bl[19] br[19] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_20 bl[20] br[20] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_21 bl[21] br[21] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_22 bl[22] br[22] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_23 bl[23] br[23] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_24 bl[24] br[24] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_25 bl[25] br[25] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_26 bl[26] br[26] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_27 bl[27] br[27] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_28 bl[28] br[28] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_29 bl[29] br[29] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_30 bl[30] br[30] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_31 bl[31] br[31] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_32 bl[32] br[32] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_33 bl[33] br[33] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_34 bl[34] br[34] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_35 bl[35] br[35] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_36 bl[36] br[36] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_37 bl[37] br[37] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_38 bl[38] br[38] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_39 bl[39] br[39] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_40 bl[40] br[40] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_41 bl[41] br[41] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_42 bl[42] br[42] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_43 bl[43] br[43] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_44 bl[44] br[44] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_45 bl[45] br[45] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_46 bl[46] br[46] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_47 bl[47] br[47] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_48 bl[48] br[48] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_49 bl[49] br[49] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_50 bl[50] br[50] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_51 bl[51] br[51] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_52 bl[52] br[52] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_53 bl[53] br[53] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_54 bl[54] br[54] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_55 bl[55] br[55] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_56 bl[56] br[56] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_57 bl[57] br[57] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_58 bl[58] br[58] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_59 bl[59] br[59] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_60 bl[60] br[60] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_61 bl[61] br[61] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_62 bl[62] br[62] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_63 bl[63] br[63] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_64 bl[64] br[64] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_65 bl[65] br[65] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_66 bl[66] br[66] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_67 bl[67] br[67] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_68 bl[68] br[68] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_69 bl[69] br[69] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_70 bl[70] br[70] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_71 bl[71] br[71] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_72 bl[72] br[72] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_73 bl[73] br[73] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_74 bl[74] br[74] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_75 bl[75] br[75] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_76 bl[76] br[76] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_77 bl[77] br[77] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_78 bl[78] br[78] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_79 bl[79] br[79] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_80 bl[80] br[80] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_81 bl[81] br[81] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_82 bl[82] br[82] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_83 bl[83] br[83] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_84 bl[84] br[84] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_85 bl[85] br[85] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_86 bl[86] br[86] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_87 bl[87] br[87] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_88 bl[88] br[88] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_89 bl[89] br[89] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_90 bl[90] br[90] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_91 bl[91] br[91] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_92 bl[92] br[92] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_93 bl[93] br[93] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_94 bl[94] br[94] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_95 bl[95] br[95] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_96 bl[96] br[96] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_97 bl[97] br[97] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_98 bl[98] br[98] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_99 bl[99] br[99] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_100 bl[100] br[100] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_101 bl[101] br[101] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_102 bl[102] br[102] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_103 bl[103] br[103] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_104 bl[104] br[104] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_105 bl[105] br[105] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_106 bl[106] br[106] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_107 bl[107] br[107] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_108 bl[108] br[108] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_109 bl[109] br[109] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_110 bl[110] br[110] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_111 bl[111] br[111] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_112 bl[112] br[112] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_113 bl[113] br[113] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_114 bl[114] br[114] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_115 bl[115] br[115] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_116 bl[116] br[116] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_117 bl[117] br[117] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_118 bl[118] br[118] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_119 bl[119] br[119] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_120 bl[120] br[120] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_121 bl[121] br[121] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_122 bl[122] br[122] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_123 bl[123] br[123] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_124 bl[124] br[124] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_125 bl[125] br[125] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_126 bl[126] br[126] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_127 bl[127] br[127] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_128 bl[128] br[128] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_129 bl[129] br[129] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_130 bl[130] br[130] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_131 bl[131] br[131] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_132 bl[132] br[132] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_133 bl[133] br[133] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_134 bl[134] br[134] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_135 bl[135] br[135] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_136 bl[136] br[136] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_137 bl[137] br[137] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_138 bl[138] br[138] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_139 bl[139] br[139] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_140 bl[140] br[140] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_141 bl[141] br[141] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_142 bl[142] br[142] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_143 bl[143] br[143] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_144 bl[144] br[144] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_145 bl[145] br[145] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_146 bl[146] br[146] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_147 bl[147] br[147] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_148 bl[148] br[148] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_149 bl[149] br[149] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_150 bl[150] br[150] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_151 bl[151] br[151] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_152 bl[152] br[152] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_153 bl[153] br[153] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_154 bl[154] br[154] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_155 bl[155] br[155] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_156 bl[156] br[156] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_157 bl[157] br[157] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_158 bl[158] br[158] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_159 bl[159] br[159] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_160 bl[160] br[160] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_161 bl[161] br[161] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_162 bl[162] br[162] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_163 bl[163] br[163] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_164 bl[164] br[164] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_165 bl[165] br[165] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_166 bl[166] br[166] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_167 bl[167] br[167] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_168 bl[168] br[168] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_169 bl[169] br[169] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_170 bl[170] br[170] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_171 bl[171] br[171] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_172 bl[172] br[172] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_173 bl[173] br[173] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_174 bl[174] br[174] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_175 bl[175] br[175] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_176 bl[176] br[176] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_177 bl[177] br[177] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_178 bl[178] br[178] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_179 bl[179] br[179] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_180 bl[180] br[180] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_181 bl[181] br[181] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_182 bl[182] br[182] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_183 bl[183] br[183] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_184 bl[184] br[184] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_185 bl[185] br[185] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_186 bl[186] br[186] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_187 bl[187] br[187] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_188 bl[188] br[188] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_189 bl[189] br[189] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_190 bl[190] br[190] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_191 bl[191] br[191] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_192 bl[192] br[192] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_193 bl[193] br[193] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_194 bl[194] br[194] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_195 bl[195] br[195] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_196 bl[196] br[196] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_197 bl[197] br[197] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_198 bl[198] br[198] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_199 bl[199] br[199] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_200 bl[200] br[200] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_201 bl[201] br[201] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_202 bl[202] br[202] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_203 bl[203] br[203] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_204 bl[204] br[204] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_205 bl[205] br[205] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_206 bl[206] br[206] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_207 bl[207] br[207] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_208 bl[208] br[208] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_209 bl[209] br[209] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_210 bl[210] br[210] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_211 bl[211] br[211] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_212 bl[212] br[212] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_213 bl[213] br[213] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_214 bl[214] br[214] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_215 bl[215] br[215] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_216 bl[216] br[216] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_217 bl[217] br[217] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_218 bl[218] br[218] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_219 bl[219] br[219] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_220 bl[220] br[220] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_221 bl[221] br[221] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_222 bl[222] br[222] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_223 bl[223] br[223] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_224 bl[224] br[224] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_225 bl[225] br[225] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_226 bl[226] br[226] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_227 bl[227] br[227] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_228 bl[228] br[228] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_229 bl[229] br[229] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_230 bl[230] br[230] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_231 bl[231] br[231] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_232 bl[232] br[232] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_233 bl[233] br[233] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_234 bl[234] br[234] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_235 bl[235] br[235] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_236 bl[236] br[236] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_237 bl[237] br[237] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_238 bl[238] br[238] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_239 bl[239] br[239] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_240 bl[240] br[240] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_241 bl[241] br[241] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_242 bl[242] br[242] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_243 bl[243] br[243] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_244 bl[244] br[244] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_245 bl[245] br[245] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_246 bl[246] br[246] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_247 bl[247] br[247] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_248 bl[248] br[248] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_249 bl[249] br[249] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_250 bl[250] br[250] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_251 bl[251] br[251] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_252 bl[252] br[252] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_253 bl[253] br[253] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_254 bl[254] br[254] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_255 bl[255] br[255] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_256 bl[256] br[256] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_257 bl[257] br[257] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_258 bl[258] br[258] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_259 bl[259] br[259] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_260 bl[260] br[260] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_261 bl[261] br[261] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_262 bl[262] br[262] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_263 bl[263] br[263] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_264 bl[264] br[264] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_265 bl[265] br[265] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_266 bl[266] br[266] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_267 bl[267] br[267] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_268 bl[268] br[268] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_269 bl[269] br[269] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_270 bl[270] br[270] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_271 bl[271] br[271] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_272 bl[272] br[272] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_273 bl[273] br[273] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_274 bl[274] br[274] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_275 bl[275] br[275] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_276 bl[276] br[276] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_277 bl[277] br[277] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_278 bl[278] br[278] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_279 bl[279] br[279] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_280 bl[280] br[280] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_281 bl[281] br[281] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_282 bl[282] br[282] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_283 bl[283] br[283] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_284 bl[284] br[284] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_285 bl[285] br[285] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_286 bl[286] br[286] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_287 bl[287] br[287] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_288 bl[288] br[288] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_289 bl[289] br[289] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_290 bl[290] br[290] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_291 bl[291] br[291] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_292 bl[292] br[292] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_293 bl[293] br[293] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_294 bl[294] br[294] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_295 bl[295] br[295] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_296 bl[296] br[296] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_297 bl[297] br[297] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_298 bl[298] br[298] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_299 bl[299] br[299] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_300 bl[300] br[300] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_301 bl[301] br[301] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_302 bl[302] br[302] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_303 bl[303] br[303] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_304 bl[304] br[304] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_305 bl[305] br[305] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_306 bl[306] br[306] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_307 bl[307] br[307] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_308 bl[308] br[308] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_309 bl[309] br[309] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_310 bl[310] br[310] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_311 bl[311] br[311] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_312 bl[312] br[312] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_313 bl[313] br[313] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_314 bl[314] br[314] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_315 bl[315] br[315] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_316 bl[316] br[316] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_317 bl[317] br[317] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_318 bl[318] br[318] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_319 bl[319] br[319] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_320 bl[320] br[320] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_321 bl[321] br[321] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_322 bl[322] br[322] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_323 bl[323] br[323] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_324 bl[324] br[324] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_325 bl[325] br[325] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_326 bl[326] br[326] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_327 bl[327] br[327] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_328 bl[328] br[328] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_329 bl[329] br[329] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_330 bl[330] br[330] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_331 bl[331] br[331] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_332 bl[332] br[332] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_333 bl[333] br[333] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_334 bl[334] br[334] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_335 bl[335] br[335] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_336 bl[336] br[336] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_337 bl[337] br[337] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_338 bl[338] br[338] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_339 bl[339] br[339] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_340 bl[340] br[340] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_341 bl[341] br[341] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_342 bl[342] br[342] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_343 bl[343] br[343] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_344 bl[344] br[344] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_345 bl[345] br[345] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_346 bl[346] br[346] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_347 bl[347] br[347] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_348 bl[348] br[348] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_349 bl[349] br[349] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_350 bl[350] br[350] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_351 bl[351] br[351] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_352 bl[352] br[352] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_353 bl[353] br[353] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_354 bl[354] br[354] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_355 bl[355] br[355] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_356 bl[356] br[356] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_357 bl[357] br[357] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_358 bl[358] br[358] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_359 bl[359] br[359] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_360 bl[360] br[360] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_361 bl[361] br[361] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_362 bl[362] br[362] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_363 bl[363] br[363] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_364 bl[364] br[364] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_365 bl[365] br[365] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_366 bl[366] br[366] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_367 bl[367] br[367] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_368 bl[368] br[368] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_369 bl[369] br[369] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_370 bl[370] br[370] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_371 bl[371] br[371] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_372 bl[372] br[372] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_373 bl[373] br[373] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_374 bl[374] br[374] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_375 bl[375] br[375] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_376 bl[376] br[376] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_377 bl[377] br[377] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_378 bl[378] br[378] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_379 bl[379] br[379] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_380 bl[380] br[380] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_381 bl[381] br[381] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_382 bl[382] br[382] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_383 bl[383] br[383] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_384 bl[384] br[384] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_385 bl[385] br[385] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_386 bl[386] br[386] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_387 bl[387] br[387] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_388 bl[388] br[388] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_389 bl[389] br[389] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_390 bl[390] br[390] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_391 bl[391] br[391] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_392 bl[392] br[392] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_393 bl[393] br[393] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_394 bl[394] br[394] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_395 bl[395] br[395] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_396 bl[396] br[396] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_397 bl[397] br[397] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_398 bl[398] br[398] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_399 bl[399] br[399] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_400 bl[400] br[400] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_401 bl[401] br[401] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_402 bl[402] br[402] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_403 bl[403] br[403] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_404 bl[404] br[404] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_405 bl[405] br[405] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_406 bl[406] br[406] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_407 bl[407] br[407] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_408 bl[408] br[408] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_409 bl[409] br[409] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_410 bl[410] br[410] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_411 bl[411] br[411] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_412 bl[412] br[412] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_413 bl[413] br[413] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_414 bl[414] br[414] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_415 bl[415] br[415] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_416 bl[416] br[416] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_417 bl[417] br[417] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_418 bl[418] br[418] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_419 bl[419] br[419] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_420 bl[420] br[420] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_421 bl[421] br[421] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_422 bl[422] br[422] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_423 bl[423] br[423] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_424 bl[424] br[424] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_425 bl[425] br[425] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_426 bl[426] br[426] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_427 bl[427] br[427] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_428 bl[428] br[428] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_429 bl[429] br[429] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_430 bl[430] br[430] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_431 bl[431] br[431] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_432 bl[432] br[432] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_433 bl[433] br[433] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_434 bl[434] br[434] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_435 bl[435] br[435] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_436 bl[436] br[436] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_437 bl[437] br[437] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_438 bl[438] br[438] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_439 bl[439] br[439] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_440 bl[440] br[440] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_441 bl[441] br[441] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_442 bl[442] br[442] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_443 bl[443] br[443] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_444 bl[444] br[444] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_445 bl[445] br[445] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_446 bl[446] br[446] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_447 bl[447] br[447] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_448 bl[448] br[448] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_449 bl[449] br[449] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_450 bl[450] br[450] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_451 bl[451] br[451] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_452 bl[452] br[452] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_453 bl[453] br[453] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_454 bl[454] br[454] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_455 bl[455] br[455] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_456 bl[456] br[456] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_457 bl[457] br[457] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_458 bl[458] br[458] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_459 bl[459] br[459] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_460 bl[460] br[460] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_461 bl[461] br[461] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_462 bl[462] br[462] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_463 bl[463] br[463] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_464 bl[464] br[464] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_465 bl[465] br[465] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_466 bl[466] br[466] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_467 bl[467] br[467] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_468 bl[468] br[468] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_469 bl[469] br[469] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_470 bl[470] br[470] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_471 bl[471] br[471] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_472 bl[472] br[472] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_473 bl[473] br[473] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_474 bl[474] br[474] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_475 bl[475] br[475] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_476 bl[476] br[476] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_477 bl[477] br[477] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_478 bl[478] br[478] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_479 bl[479] br[479] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_480 bl[480] br[480] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_481 bl[481] br[481] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_482 bl[482] br[482] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_483 bl[483] br[483] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_484 bl[484] br[484] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_485 bl[485] br[485] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_486 bl[486] br[486] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_487 bl[487] br[487] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_488 bl[488] br[488] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_489 bl[489] br[489] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_490 bl[490] br[490] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_491 bl[491] br[491] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_492 bl[492] br[492] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_493 bl[493] br[493] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_494 bl[494] br[494] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_495 bl[495] br[495] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_496 bl[496] br[496] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_497 bl[497] br[497] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_498 bl[498] br[498] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_499 bl[499] br[499] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_500 bl[500] br[500] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_501 bl[501] br[501] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_502 bl[502] br[502] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_503 bl[503] br[503] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_504 bl[504] br[504] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_505 bl[505] br[505] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_506 bl[506] br[506] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_507 bl[507] br[507] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_508 bl[508] br[508] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_509 bl[509] br[509] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_510 bl[510] br[510] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_14_511 bl[511] br[511] vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xcell_15_0 bl[0] br[0] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_1 bl[1] br[1] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_2 bl[2] br[2] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_3 bl[3] br[3] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_4 bl[4] br[4] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_5 bl[5] br[5] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_6 bl[6] br[6] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_7 bl[7] br[7] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_8 bl[8] br[8] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_9 bl[9] br[9] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_10 bl[10] br[10] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_11 bl[11] br[11] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_12 bl[12] br[12] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_13 bl[13] br[13] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_14 bl[14] br[14] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_15 bl[15] br[15] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_16 bl[16] br[16] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_17 bl[17] br[17] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_18 bl[18] br[18] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_19 bl[19] br[19] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_20 bl[20] br[20] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_21 bl[21] br[21] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_22 bl[22] br[22] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_23 bl[23] br[23] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_24 bl[24] br[24] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_25 bl[25] br[25] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_26 bl[26] br[26] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_27 bl[27] br[27] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_28 bl[28] br[28] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_29 bl[29] br[29] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_30 bl[30] br[30] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_31 bl[31] br[31] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_32 bl[32] br[32] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_33 bl[33] br[33] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_34 bl[34] br[34] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_35 bl[35] br[35] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_36 bl[36] br[36] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_37 bl[37] br[37] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_38 bl[38] br[38] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_39 bl[39] br[39] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_40 bl[40] br[40] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_41 bl[41] br[41] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_42 bl[42] br[42] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_43 bl[43] br[43] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_44 bl[44] br[44] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_45 bl[45] br[45] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_46 bl[46] br[46] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_47 bl[47] br[47] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_48 bl[48] br[48] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_49 bl[49] br[49] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_50 bl[50] br[50] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_51 bl[51] br[51] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_52 bl[52] br[52] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_53 bl[53] br[53] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_54 bl[54] br[54] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_55 bl[55] br[55] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_56 bl[56] br[56] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_57 bl[57] br[57] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_58 bl[58] br[58] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_59 bl[59] br[59] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_60 bl[60] br[60] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_61 bl[61] br[61] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_62 bl[62] br[62] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_63 bl[63] br[63] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_64 bl[64] br[64] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_65 bl[65] br[65] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_66 bl[66] br[66] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_67 bl[67] br[67] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_68 bl[68] br[68] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_69 bl[69] br[69] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_70 bl[70] br[70] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_71 bl[71] br[71] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_72 bl[72] br[72] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_73 bl[73] br[73] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_74 bl[74] br[74] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_75 bl[75] br[75] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_76 bl[76] br[76] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_77 bl[77] br[77] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_78 bl[78] br[78] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_79 bl[79] br[79] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_80 bl[80] br[80] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_81 bl[81] br[81] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_82 bl[82] br[82] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_83 bl[83] br[83] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_84 bl[84] br[84] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_85 bl[85] br[85] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_86 bl[86] br[86] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_87 bl[87] br[87] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_88 bl[88] br[88] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_89 bl[89] br[89] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_90 bl[90] br[90] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_91 bl[91] br[91] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_92 bl[92] br[92] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_93 bl[93] br[93] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_94 bl[94] br[94] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_95 bl[95] br[95] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_96 bl[96] br[96] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_97 bl[97] br[97] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_98 bl[98] br[98] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_99 bl[99] br[99] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_100 bl[100] br[100] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_101 bl[101] br[101] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_102 bl[102] br[102] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_103 bl[103] br[103] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_104 bl[104] br[104] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_105 bl[105] br[105] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_106 bl[106] br[106] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_107 bl[107] br[107] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_108 bl[108] br[108] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_109 bl[109] br[109] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_110 bl[110] br[110] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_111 bl[111] br[111] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_112 bl[112] br[112] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_113 bl[113] br[113] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_114 bl[114] br[114] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_115 bl[115] br[115] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_116 bl[116] br[116] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_117 bl[117] br[117] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_118 bl[118] br[118] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_119 bl[119] br[119] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_120 bl[120] br[120] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_121 bl[121] br[121] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_122 bl[122] br[122] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_123 bl[123] br[123] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_124 bl[124] br[124] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_125 bl[125] br[125] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_126 bl[126] br[126] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_127 bl[127] br[127] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_128 bl[128] br[128] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_129 bl[129] br[129] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_130 bl[130] br[130] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_131 bl[131] br[131] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_132 bl[132] br[132] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_133 bl[133] br[133] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_134 bl[134] br[134] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_135 bl[135] br[135] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_136 bl[136] br[136] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_137 bl[137] br[137] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_138 bl[138] br[138] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_139 bl[139] br[139] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_140 bl[140] br[140] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_141 bl[141] br[141] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_142 bl[142] br[142] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_143 bl[143] br[143] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_144 bl[144] br[144] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_145 bl[145] br[145] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_146 bl[146] br[146] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_147 bl[147] br[147] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_148 bl[148] br[148] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_149 bl[149] br[149] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_150 bl[150] br[150] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_151 bl[151] br[151] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_152 bl[152] br[152] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_153 bl[153] br[153] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_154 bl[154] br[154] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_155 bl[155] br[155] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_156 bl[156] br[156] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_157 bl[157] br[157] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_158 bl[158] br[158] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_159 bl[159] br[159] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_160 bl[160] br[160] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_161 bl[161] br[161] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_162 bl[162] br[162] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_163 bl[163] br[163] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_164 bl[164] br[164] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_165 bl[165] br[165] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_166 bl[166] br[166] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_167 bl[167] br[167] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_168 bl[168] br[168] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_169 bl[169] br[169] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_170 bl[170] br[170] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_171 bl[171] br[171] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_172 bl[172] br[172] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_173 bl[173] br[173] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_174 bl[174] br[174] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_175 bl[175] br[175] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_176 bl[176] br[176] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_177 bl[177] br[177] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_178 bl[178] br[178] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_179 bl[179] br[179] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_180 bl[180] br[180] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_181 bl[181] br[181] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_182 bl[182] br[182] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_183 bl[183] br[183] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_184 bl[184] br[184] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_185 bl[185] br[185] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_186 bl[186] br[186] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_187 bl[187] br[187] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_188 bl[188] br[188] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_189 bl[189] br[189] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_190 bl[190] br[190] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_191 bl[191] br[191] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_192 bl[192] br[192] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_193 bl[193] br[193] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_194 bl[194] br[194] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_195 bl[195] br[195] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_196 bl[196] br[196] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_197 bl[197] br[197] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_198 bl[198] br[198] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_199 bl[199] br[199] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_200 bl[200] br[200] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_201 bl[201] br[201] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_202 bl[202] br[202] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_203 bl[203] br[203] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_204 bl[204] br[204] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_205 bl[205] br[205] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_206 bl[206] br[206] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_207 bl[207] br[207] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_208 bl[208] br[208] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_209 bl[209] br[209] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_210 bl[210] br[210] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_211 bl[211] br[211] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_212 bl[212] br[212] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_213 bl[213] br[213] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_214 bl[214] br[214] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_215 bl[215] br[215] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_216 bl[216] br[216] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_217 bl[217] br[217] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_218 bl[218] br[218] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_219 bl[219] br[219] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_220 bl[220] br[220] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_221 bl[221] br[221] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_222 bl[222] br[222] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_223 bl[223] br[223] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_224 bl[224] br[224] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_225 bl[225] br[225] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_226 bl[226] br[226] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_227 bl[227] br[227] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_228 bl[228] br[228] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_229 bl[229] br[229] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_230 bl[230] br[230] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_231 bl[231] br[231] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_232 bl[232] br[232] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_233 bl[233] br[233] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_234 bl[234] br[234] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_235 bl[235] br[235] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_236 bl[236] br[236] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_237 bl[237] br[237] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_238 bl[238] br[238] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_239 bl[239] br[239] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_240 bl[240] br[240] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_241 bl[241] br[241] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_242 bl[242] br[242] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_243 bl[243] br[243] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_244 bl[244] br[244] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_245 bl[245] br[245] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_246 bl[246] br[246] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_247 bl[247] br[247] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_248 bl[248] br[248] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_249 bl[249] br[249] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_250 bl[250] br[250] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_251 bl[251] br[251] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_252 bl[252] br[252] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_253 bl[253] br[253] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_254 bl[254] br[254] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_255 bl[255] br[255] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_256 bl[256] br[256] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_257 bl[257] br[257] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_258 bl[258] br[258] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_259 bl[259] br[259] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_260 bl[260] br[260] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_261 bl[261] br[261] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_262 bl[262] br[262] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_263 bl[263] br[263] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_264 bl[264] br[264] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_265 bl[265] br[265] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_266 bl[266] br[266] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_267 bl[267] br[267] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_268 bl[268] br[268] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_269 bl[269] br[269] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_270 bl[270] br[270] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_271 bl[271] br[271] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_272 bl[272] br[272] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_273 bl[273] br[273] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_274 bl[274] br[274] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_275 bl[275] br[275] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_276 bl[276] br[276] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_277 bl[277] br[277] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_278 bl[278] br[278] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_279 bl[279] br[279] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_280 bl[280] br[280] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_281 bl[281] br[281] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_282 bl[282] br[282] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_283 bl[283] br[283] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_284 bl[284] br[284] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_285 bl[285] br[285] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_286 bl[286] br[286] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_287 bl[287] br[287] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_288 bl[288] br[288] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_289 bl[289] br[289] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_290 bl[290] br[290] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_291 bl[291] br[291] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_292 bl[292] br[292] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_293 bl[293] br[293] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_294 bl[294] br[294] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_295 bl[295] br[295] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_296 bl[296] br[296] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_297 bl[297] br[297] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_298 bl[298] br[298] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_299 bl[299] br[299] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_300 bl[300] br[300] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_301 bl[301] br[301] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_302 bl[302] br[302] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_303 bl[303] br[303] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_304 bl[304] br[304] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_305 bl[305] br[305] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_306 bl[306] br[306] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_307 bl[307] br[307] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_308 bl[308] br[308] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_309 bl[309] br[309] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_310 bl[310] br[310] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_311 bl[311] br[311] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_312 bl[312] br[312] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_313 bl[313] br[313] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_314 bl[314] br[314] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_315 bl[315] br[315] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_316 bl[316] br[316] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_317 bl[317] br[317] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_318 bl[318] br[318] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_319 bl[319] br[319] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_320 bl[320] br[320] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_321 bl[321] br[321] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_322 bl[322] br[322] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_323 bl[323] br[323] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_324 bl[324] br[324] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_325 bl[325] br[325] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_326 bl[326] br[326] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_327 bl[327] br[327] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_328 bl[328] br[328] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_329 bl[329] br[329] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_330 bl[330] br[330] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_331 bl[331] br[331] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_332 bl[332] br[332] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_333 bl[333] br[333] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_334 bl[334] br[334] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_335 bl[335] br[335] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_336 bl[336] br[336] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_337 bl[337] br[337] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_338 bl[338] br[338] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_339 bl[339] br[339] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_340 bl[340] br[340] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_341 bl[341] br[341] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_342 bl[342] br[342] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_343 bl[343] br[343] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_344 bl[344] br[344] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_345 bl[345] br[345] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_346 bl[346] br[346] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_347 bl[347] br[347] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_348 bl[348] br[348] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_349 bl[349] br[349] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_350 bl[350] br[350] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_351 bl[351] br[351] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_352 bl[352] br[352] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_353 bl[353] br[353] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_354 bl[354] br[354] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_355 bl[355] br[355] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_356 bl[356] br[356] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_357 bl[357] br[357] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_358 bl[358] br[358] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_359 bl[359] br[359] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_360 bl[360] br[360] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_361 bl[361] br[361] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_362 bl[362] br[362] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_363 bl[363] br[363] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_364 bl[364] br[364] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_365 bl[365] br[365] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_366 bl[366] br[366] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_367 bl[367] br[367] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_368 bl[368] br[368] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_369 bl[369] br[369] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_370 bl[370] br[370] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_371 bl[371] br[371] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_372 bl[372] br[372] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_373 bl[373] br[373] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_374 bl[374] br[374] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_375 bl[375] br[375] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_376 bl[376] br[376] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_377 bl[377] br[377] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_378 bl[378] br[378] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_379 bl[379] br[379] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_380 bl[380] br[380] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_381 bl[381] br[381] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_382 bl[382] br[382] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_383 bl[383] br[383] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_384 bl[384] br[384] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_385 bl[385] br[385] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_386 bl[386] br[386] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_387 bl[387] br[387] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_388 bl[388] br[388] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_389 bl[389] br[389] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_390 bl[390] br[390] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_391 bl[391] br[391] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_392 bl[392] br[392] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_393 bl[393] br[393] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_394 bl[394] br[394] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_395 bl[395] br[395] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_396 bl[396] br[396] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_397 bl[397] br[397] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_398 bl[398] br[398] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_399 bl[399] br[399] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_400 bl[400] br[400] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_401 bl[401] br[401] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_402 bl[402] br[402] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_403 bl[403] br[403] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_404 bl[404] br[404] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_405 bl[405] br[405] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_406 bl[406] br[406] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_407 bl[407] br[407] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_408 bl[408] br[408] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_409 bl[409] br[409] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_410 bl[410] br[410] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_411 bl[411] br[411] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_412 bl[412] br[412] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_413 bl[413] br[413] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_414 bl[414] br[414] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_415 bl[415] br[415] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_416 bl[416] br[416] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_417 bl[417] br[417] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_418 bl[418] br[418] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_419 bl[419] br[419] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_420 bl[420] br[420] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_421 bl[421] br[421] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_422 bl[422] br[422] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_423 bl[423] br[423] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_424 bl[424] br[424] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_425 bl[425] br[425] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_426 bl[426] br[426] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_427 bl[427] br[427] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_428 bl[428] br[428] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_429 bl[429] br[429] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_430 bl[430] br[430] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_431 bl[431] br[431] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_432 bl[432] br[432] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_433 bl[433] br[433] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_434 bl[434] br[434] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_435 bl[435] br[435] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_436 bl[436] br[436] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_437 bl[437] br[437] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_438 bl[438] br[438] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_439 bl[439] br[439] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_440 bl[440] br[440] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_441 bl[441] br[441] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_442 bl[442] br[442] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_443 bl[443] br[443] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_444 bl[444] br[444] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_445 bl[445] br[445] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_446 bl[446] br[446] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_447 bl[447] br[447] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_448 bl[448] br[448] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_449 bl[449] br[449] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_450 bl[450] br[450] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_451 bl[451] br[451] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_452 bl[452] br[452] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_453 bl[453] br[453] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_454 bl[454] br[454] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_455 bl[455] br[455] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_456 bl[456] br[456] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_457 bl[457] br[457] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_458 bl[458] br[458] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_459 bl[459] br[459] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_460 bl[460] br[460] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_461 bl[461] br[461] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_462 bl[462] br[462] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_463 bl[463] br[463] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_464 bl[464] br[464] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_465 bl[465] br[465] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_466 bl[466] br[466] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_467 bl[467] br[467] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_468 bl[468] br[468] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_469 bl[469] br[469] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_470 bl[470] br[470] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_471 bl[471] br[471] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_472 bl[472] br[472] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_473 bl[473] br[473] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_474 bl[474] br[474] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_475 bl[475] br[475] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_476 bl[476] br[476] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_477 bl[477] br[477] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_478 bl[478] br[478] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_479 bl[479] br[479] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_480 bl[480] br[480] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_481 bl[481] br[481] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_482 bl[482] br[482] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_483 bl[483] br[483] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_484 bl[484] br[484] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_485 bl[485] br[485] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_486 bl[486] br[486] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_487 bl[487] br[487] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_488 bl[488] br[488] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_489 bl[489] br[489] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_490 bl[490] br[490] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_491 bl[491] br[491] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_492 bl[492] br[492] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_493 bl[493] br[493] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_494 bl[494] br[494] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_495 bl[495] br[495] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_496 bl[496] br[496] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_497 bl[497] br[497] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_498 bl[498] br[498] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_499 bl[499] br[499] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_500 bl[500] br[500] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_501 bl[501] br[501] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_502 bl[502] br[502] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_503 bl[503] br[503] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_504 bl[504] br[504] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_505 bl[505] br[505] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_506 bl[506] br[506] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_507 bl[507] br[507] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_508 bl[508] br[508] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_509 bl[509] br[509] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_510 bl[510] br[510] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_15_511 bl[511] br[511] vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xcell_16_0 bl[0] br[0] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_1 bl[1] br[1] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_2 bl[2] br[2] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_3 bl[3] br[3] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_4 bl[4] br[4] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_5 bl[5] br[5] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_6 bl[6] br[6] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_7 bl[7] br[7] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_8 bl[8] br[8] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_9 bl[9] br[9] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_10 bl[10] br[10] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_11 bl[11] br[11] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_12 bl[12] br[12] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_13 bl[13] br[13] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_14 bl[14] br[14] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_15 bl[15] br[15] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_16 bl[16] br[16] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_17 bl[17] br[17] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_18 bl[18] br[18] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_19 bl[19] br[19] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_20 bl[20] br[20] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_21 bl[21] br[21] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_22 bl[22] br[22] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_23 bl[23] br[23] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_24 bl[24] br[24] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_25 bl[25] br[25] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_26 bl[26] br[26] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_27 bl[27] br[27] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_28 bl[28] br[28] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_29 bl[29] br[29] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_30 bl[30] br[30] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_31 bl[31] br[31] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_32 bl[32] br[32] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_33 bl[33] br[33] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_34 bl[34] br[34] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_35 bl[35] br[35] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_36 bl[36] br[36] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_37 bl[37] br[37] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_38 bl[38] br[38] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_39 bl[39] br[39] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_40 bl[40] br[40] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_41 bl[41] br[41] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_42 bl[42] br[42] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_43 bl[43] br[43] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_44 bl[44] br[44] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_45 bl[45] br[45] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_46 bl[46] br[46] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_47 bl[47] br[47] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_48 bl[48] br[48] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_49 bl[49] br[49] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_50 bl[50] br[50] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_51 bl[51] br[51] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_52 bl[52] br[52] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_53 bl[53] br[53] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_54 bl[54] br[54] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_55 bl[55] br[55] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_56 bl[56] br[56] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_57 bl[57] br[57] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_58 bl[58] br[58] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_59 bl[59] br[59] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_60 bl[60] br[60] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_61 bl[61] br[61] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_62 bl[62] br[62] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_63 bl[63] br[63] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_64 bl[64] br[64] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_65 bl[65] br[65] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_66 bl[66] br[66] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_67 bl[67] br[67] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_68 bl[68] br[68] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_69 bl[69] br[69] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_70 bl[70] br[70] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_71 bl[71] br[71] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_72 bl[72] br[72] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_73 bl[73] br[73] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_74 bl[74] br[74] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_75 bl[75] br[75] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_76 bl[76] br[76] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_77 bl[77] br[77] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_78 bl[78] br[78] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_79 bl[79] br[79] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_80 bl[80] br[80] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_81 bl[81] br[81] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_82 bl[82] br[82] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_83 bl[83] br[83] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_84 bl[84] br[84] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_85 bl[85] br[85] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_86 bl[86] br[86] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_87 bl[87] br[87] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_88 bl[88] br[88] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_89 bl[89] br[89] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_90 bl[90] br[90] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_91 bl[91] br[91] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_92 bl[92] br[92] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_93 bl[93] br[93] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_94 bl[94] br[94] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_95 bl[95] br[95] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_96 bl[96] br[96] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_97 bl[97] br[97] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_98 bl[98] br[98] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_99 bl[99] br[99] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_100 bl[100] br[100] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_101 bl[101] br[101] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_102 bl[102] br[102] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_103 bl[103] br[103] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_104 bl[104] br[104] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_105 bl[105] br[105] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_106 bl[106] br[106] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_107 bl[107] br[107] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_108 bl[108] br[108] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_109 bl[109] br[109] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_110 bl[110] br[110] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_111 bl[111] br[111] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_112 bl[112] br[112] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_113 bl[113] br[113] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_114 bl[114] br[114] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_115 bl[115] br[115] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_116 bl[116] br[116] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_117 bl[117] br[117] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_118 bl[118] br[118] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_119 bl[119] br[119] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_120 bl[120] br[120] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_121 bl[121] br[121] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_122 bl[122] br[122] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_123 bl[123] br[123] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_124 bl[124] br[124] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_125 bl[125] br[125] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_126 bl[126] br[126] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_127 bl[127] br[127] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_128 bl[128] br[128] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_129 bl[129] br[129] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_130 bl[130] br[130] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_131 bl[131] br[131] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_132 bl[132] br[132] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_133 bl[133] br[133] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_134 bl[134] br[134] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_135 bl[135] br[135] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_136 bl[136] br[136] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_137 bl[137] br[137] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_138 bl[138] br[138] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_139 bl[139] br[139] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_140 bl[140] br[140] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_141 bl[141] br[141] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_142 bl[142] br[142] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_143 bl[143] br[143] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_144 bl[144] br[144] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_145 bl[145] br[145] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_146 bl[146] br[146] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_147 bl[147] br[147] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_148 bl[148] br[148] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_149 bl[149] br[149] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_150 bl[150] br[150] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_151 bl[151] br[151] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_152 bl[152] br[152] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_153 bl[153] br[153] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_154 bl[154] br[154] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_155 bl[155] br[155] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_156 bl[156] br[156] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_157 bl[157] br[157] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_158 bl[158] br[158] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_159 bl[159] br[159] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_160 bl[160] br[160] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_161 bl[161] br[161] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_162 bl[162] br[162] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_163 bl[163] br[163] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_164 bl[164] br[164] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_165 bl[165] br[165] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_166 bl[166] br[166] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_167 bl[167] br[167] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_168 bl[168] br[168] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_169 bl[169] br[169] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_170 bl[170] br[170] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_171 bl[171] br[171] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_172 bl[172] br[172] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_173 bl[173] br[173] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_174 bl[174] br[174] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_175 bl[175] br[175] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_176 bl[176] br[176] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_177 bl[177] br[177] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_178 bl[178] br[178] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_179 bl[179] br[179] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_180 bl[180] br[180] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_181 bl[181] br[181] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_182 bl[182] br[182] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_183 bl[183] br[183] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_184 bl[184] br[184] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_185 bl[185] br[185] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_186 bl[186] br[186] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_187 bl[187] br[187] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_188 bl[188] br[188] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_189 bl[189] br[189] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_190 bl[190] br[190] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_191 bl[191] br[191] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_192 bl[192] br[192] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_193 bl[193] br[193] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_194 bl[194] br[194] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_195 bl[195] br[195] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_196 bl[196] br[196] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_197 bl[197] br[197] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_198 bl[198] br[198] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_199 bl[199] br[199] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_200 bl[200] br[200] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_201 bl[201] br[201] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_202 bl[202] br[202] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_203 bl[203] br[203] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_204 bl[204] br[204] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_205 bl[205] br[205] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_206 bl[206] br[206] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_207 bl[207] br[207] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_208 bl[208] br[208] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_209 bl[209] br[209] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_210 bl[210] br[210] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_211 bl[211] br[211] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_212 bl[212] br[212] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_213 bl[213] br[213] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_214 bl[214] br[214] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_215 bl[215] br[215] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_216 bl[216] br[216] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_217 bl[217] br[217] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_218 bl[218] br[218] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_219 bl[219] br[219] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_220 bl[220] br[220] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_221 bl[221] br[221] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_222 bl[222] br[222] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_223 bl[223] br[223] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_224 bl[224] br[224] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_225 bl[225] br[225] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_226 bl[226] br[226] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_227 bl[227] br[227] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_228 bl[228] br[228] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_229 bl[229] br[229] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_230 bl[230] br[230] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_231 bl[231] br[231] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_232 bl[232] br[232] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_233 bl[233] br[233] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_234 bl[234] br[234] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_235 bl[235] br[235] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_236 bl[236] br[236] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_237 bl[237] br[237] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_238 bl[238] br[238] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_239 bl[239] br[239] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_240 bl[240] br[240] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_241 bl[241] br[241] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_242 bl[242] br[242] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_243 bl[243] br[243] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_244 bl[244] br[244] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_245 bl[245] br[245] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_246 bl[246] br[246] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_247 bl[247] br[247] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_248 bl[248] br[248] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_249 bl[249] br[249] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_250 bl[250] br[250] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_251 bl[251] br[251] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_252 bl[252] br[252] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_253 bl[253] br[253] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_254 bl[254] br[254] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_255 bl[255] br[255] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_256 bl[256] br[256] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_257 bl[257] br[257] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_258 bl[258] br[258] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_259 bl[259] br[259] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_260 bl[260] br[260] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_261 bl[261] br[261] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_262 bl[262] br[262] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_263 bl[263] br[263] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_264 bl[264] br[264] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_265 bl[265] br[265] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_266 bl[266] br[266] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_267 bl[267] br[267] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_268 bl[268] br[268] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_269 bl[269] br[269] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_270 bl[270] br[270] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_271 bl[271] br[271] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_272 bl[272] br[272] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_273 bl[273] br[273] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_274 bl[274] br[274] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_275 bl[275] br[275] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_276 bl[276] br[276] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_277 bl[277] br[277] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_278 bl[278] br[278] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_279 bl[279] br[279] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_280 bl[280] br[280] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_281 bl[281] br[281] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_282 bl[282] br[282] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_283 bl[283] br[283] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_284 bl[284] br[284] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_285 bl[285] br[285] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_286 bl[286] br[286] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_287 bl[287] br[287] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_288 bl[288] br[288] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_289 bl[289] br[289] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_290 bl[290] br[290] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_291 bl[291] br[291] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_292 bl[292] br[292] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_293 bl[293] br[293] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_294 bl[294] br[294] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_295 bl[295] br[295] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_296 bl[296] br[296] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_297 bl[297] br[297] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_298 bl[298] br[298] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_299 bl[299] br[299] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_300 bl[300] br[300] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_301 bl[301] br[301] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_302 bl[302] br[302] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_303 bl[303] br[303] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_304 bl[304] br[304] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_305 bl[305] br[305] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_306 bl[306] br[306] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_307 bl[307] br[307] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_308 bl[308] br[308] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_309 bl[309] br[309] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_310 bl[310] br[310] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_311 bl[311] br[311] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_312 bl[312] br[312] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_313 bl[313] br[313] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_314 bl[314] br[314] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_315 bl[315] br[315] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_316 bl[316] br[316] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_317 bl[317] br[317] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_318 bl[318] br[318] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_319 bl[319] br[319] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_320 bl[320] br[320] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_321 bl[321] br[321] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_322 bl[322] br[322] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_323 bl[323] br[323] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_324 bl[324] br[324] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_325 bl[325] br[325] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_326 bl[326] br[326] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_327 bl[327] br[327] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_328 bl[328] br[328] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_329 bl[329] br[329] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_330 bl[330] br[330] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_331 bl[331] br[331] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_332 bl[332] br[332] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_333 bl[333] br[333] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_334 bl[334] br[334] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_335 bl[335] br[335] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_336 bl[336] br[336] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_337 bl[337] br[337] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_338 bl[338] br[338] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_339 bl[339] br[339] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_340 bl[340] br[340] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_341 bl[341] br[341] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_342 bl[342] br[342] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_343 bl[343] br[343] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_344 bl[344] br[344] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_345 bl[345] br[345] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_346 bl[346] br[346] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_347 bl[347] br[347] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_348 bl[348] br[348] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_349 bl[349] br[349] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_350 bl[350] br[350] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_351 bl[351] br[351] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_352 bl[352] br[352] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_353 bl[353] br[353] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_354 bl[354] br[354] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_355 bl[355] br[355] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_356 bl[356] br[356] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_357 bl[357] br[357] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_358 bl[358] br[358] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_359 bl[359] br[359] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_360 bl[360] br[360] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_361 bl[361] br[361] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_362 bl[362] br[362] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_363 bl[363] br[363] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_364 bl[364] br[364] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_365 bl[365] br[365] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_366 bl[366] br[366] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_367 bl[367] br[367] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_368 bl[368] br[368] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_369 bl[369] br[369] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_370 bl[370] br[370] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_371 bl[371] br[371] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_372 bl[372] br[372] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_373 bl[373] br[373] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_374 bl[374] br[374] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_375 bl[375] br[375] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_376 bl[376] br[376] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_377 bl[377] br[377] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_378 bl[378] br[378] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_379 bl[379] br[379] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_380 bl[380] br[380] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_381 bl[381] br[381] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_382 bl[382] br[382] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_383 bl[383] br[383] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_384 bl[384] br[384] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_385 bl[385] br[385] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_386 bl[386] br[386] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_387 bl[387] br[387] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_388 bl[388] br[388] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_389 bl[389] br[389] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_390 bl[390] br[390] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_391 bl[391] br[391] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_392 bl[392] br[392] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_393 bl[393] br[393] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_394 bl[394] br[394] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_395 bl[395] br[395] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_396 bl[396] br[396] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_397 bl[397] br[397] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_398 bl[398] br[398] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_399 bl[399] br[399] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_400 bl[400] br[400] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_401 bl[401] br[401] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_402 bl[402] br[402] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_403 bl[403] br[403] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_404 bl[404] br[404] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_405 bl[405] br[405] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_406 bl[406] br[406] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_407 bl[407] br[407] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_408 bl[408] br[408] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_409 bl[409] br[409] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_410 bl[410] br[410] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_411 bl[411] br[411] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_412 bl[412] br[412] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_413 bl[413] br[413] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_414 bl[414] br[414] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_415 bl[415] br[415] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_416 bl[416] br[416] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_417 bl[417] br[417] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_418 bl[418] br[418] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_419 bl[419] br[419] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_420 bl[420] br[420] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_421 bl[421] br[421] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_422 bl[422] br[422] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_423 bl[423] br[423] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_424 bl[424] br[424] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_425 bl[425] br[425] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_426 bl[426] br[426] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_427 bl[427] br[427] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_428 bl[428] br[428] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_429 bl[429] br[429] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_430 bl[430] br[430] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_431 bl[431] br[431] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_432 bl[432] br[432] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_433 bl[433] br[433] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_434 bl[434] br[434] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_435 bl[435] br[435] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_436 bl[436] br[436] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_437 bl[437] br[437] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_438 bl[438] br[438] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_439 bl[439] br[439] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_440 bl[440] br[440] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_441 bl[441] br[441] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_442 bl[442] br[442] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_443 bl[443] br[443] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_444 bl[444] br[444] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_445 bl[445] br[445] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_446 bl[446] br[446] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_447 bl[447] br[447] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_448 bl[448] br[448] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_449 bl[449] br[449] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_450 bl[450] br[450] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_451 bl[451] br[451] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_452 bl[452] br[452] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_453 bl[453] br[453] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_454 bl[454] br[454] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_455 bl[455] br[455] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_456 bl[456] br[456] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_457 bl[457] br[457] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_458 bl[458] br[458] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_459 bl[459] br[459] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_460 bl[460] br[460] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_461 bl[461] br[461] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_462 bl[462] br[462] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_463 bl[463] br[463] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_464 bl[464] br[464] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_465 bl[465] br[465] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_466 bl[466] br[466] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_467 bl[467] br[467] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_468 bl[468] br[468] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_469 bl[469] br[469] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_470 bl[470] br[470] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_471 bl[471] br[471] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_472 bl[472] br[472] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_473 bl[473] br[473] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_474 bl[474] br[474] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_475 bl[475] br[475] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_476 bl[476] br[476] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_477 bl[477] br[477] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_478 bl[478] br[478] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_479 bl[479] br[479] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_480 bl[480] br[480] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_481 bl[481] br[481] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_482 bl[482] br[482] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_483 bl[483] br[483] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_484 bl[484] br[484] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_485 bl[485] br[485] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_486 bl[486] br[486] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_487 bl[487] br[487] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_488 bl[488] br[488] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_489 bl[489] br[489] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_490 bl[490] br[490] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_491 bl[491] br[491] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_492 bl[492] br[492] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_493 bl[493] br[493] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_494 bl[494] br[494] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_495 bl[495] br[495] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_496 bl[496] br[496] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_497 bl[497] br[497] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_498 bl[498] br[498] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_499 bl[499] br[499] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_500 bl[500] br[500] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_501 bl[501] br[501] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_502 bl[502] br[502] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_503 bl[503] br[503] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_504 bl[504] br[504] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_505 bl[505] br[505] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_506 bl[506] br[506] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_507 bl[507] br[507] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_508 bl[508] br[508] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_509 bl[509] br[509] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_510 bl[510] br[510] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_16_511 bl[511] br[511] vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xcell_17_0 bl[0] br[0] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_1 bl[1] br[1] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_2 bl[2] br[2] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_3 bl[3] br[3] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_4 bl[4] br[4] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_5 bl[5] br[5] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_6 bl[6] br[6] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_7 bl[7] br[7] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_8 bl[8] br[8] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_9 bl[9] br[9] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_10 bl[10] br[10] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_11 bl[11] br[11] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_12 bl[12] br[12] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_13 bl[13] br[13] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_14 bl[14] br[14] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_15 bl[15] br[15] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_16 bl[16] br[16] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_17 bl[17] br[17] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_18 bl[18] br[18] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_19 bl[19] br[19] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_20 bl[20] br[20] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_21 bl[21] br[21] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_22 bl[22] br[22] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_23 bl[23] br[23] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_24 bl[24] br[24] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_25 bl[25] br[25] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_26 bl[26] br[26] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_27 bl[27] br[27] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_28 bl[28] br[28] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_29 bl[29] br[29] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_30 bl[30] br[30] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_31 bl[31] br[31] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_32 bl[32] br[32] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_33 bl[33] br[33] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_34 bl[34] br[34] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_35 bl[35] br[35] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_36 bl[36] br[36] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_37 bl[37] br[37] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_38 bl[38] br[38] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_39 bl[39] br[39] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_40 bl[40] br[40] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_41 bl[41] br[41] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_42 bl[42] br[42] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_43 bl[43] br[43] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_44 bl[44] br[44] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_45 bl[45] br[45] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_46 bl[46] br[46] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_47 bl[47] br[47] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_48 bl[48] br[48] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_49 bl[49] br[49] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_50 bl[50] br[50] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_51 bl[51] br[51] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_52 bl[52] br[52] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_53 bl[53] br[53] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_54 bl[54] br[54] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_55 bl[55] br[55] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_56 bl[56] br[56] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_57 bl[57] br[57] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_58 bl[58] br[58] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_59 bl[59] br[59] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_60 bl[60] br[60] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_61 bl[61] br[61] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_62 bl[62] br[62] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_63 bl[63] br[63] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_64 bl[64] br[64] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_65 bl[65] br[65] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_66 bl[66] br[66] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_67 bl[67] br[67] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_68 bl[68] br[68] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_69 bl[69] br[69] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_70 bl[70] br[70] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_71 bl[71] br[71] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_72 bl[72] br[72] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_73 bl[73] br[73] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_74 bl[74] br[74] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_75 bl[75] br[75] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_76 bl[76] br[76] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_77 bl[77] br[77] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_78 bl[78] br[78] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_79 bl[79] br[79] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_80 bl[80] br[80] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_81 bl[81] br[81] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_82 bl[82] br[82] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_83 bl[83] br[83] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_84 bl[84] br[84] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_85 bl[85] br[85] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_86 bl[86] br[86] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_87 bl[87] br[87] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_88 bl[88] br[88] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_89 bl[89] br[89] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_90 bl[90] br[90] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_91 bl[91] br[91] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_92 bl[92] br[92] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_93 bl[93] br[93] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_94 bl[94] br[94] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_95 bl[95] br[95] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_96 bl[96] br[96] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_97 bl[97] br[97] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_98 bl[98] br[98] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_99 bl[99] br[99] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_100 bl[100] br[100] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_101 bl[101] br[101] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_102 bl[102] br[102] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_103 bl[103] br[103] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_104 bl[104] br[104] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_105 bl[105] br[105] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_106 bl[106] br[106] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_107 bl[107] br[107] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_108 bl[108] br[108] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_109 bl[109] br[109] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_110 bl[110] br[110] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_111 bl[111] br[111] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_112 bl[112] br[112] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_113 bl[113] br[113] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_114 bl[114] br[114] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_115 bl[115] br[115] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_116 bl[116] br[116] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_117 bl[117] br[117] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_118 bl[118] br[118] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_119 bl[119] br[119] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_120 bl[120] br[120] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_121 bl[121] br[121] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_122 bl[122] br[122] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_123 bl[123] br[123] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_124 bl[124] br[124] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_125 bl[125] br[125] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_126 bl[126] br[126] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_127 bl[127] br[127] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_128 bl[128] br[128] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_129 bl[129] br[129] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_130 bl[130] br[130] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_131 bl[131] br[131] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_132 bl[132] br[132] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_133 bl[133] br[133] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_134 bl[134] br[134] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_135 bl[135] br[135] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_136 bl[136] br[136] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_137 bl[137] br[137] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_138 bl[138] br[138] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_139 bl[139] br[139] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_140 bl[140] br[140] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_141 bl[141] br[141] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_142 bl[142] br[142] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_143 bl[143] br[143] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_144 bl[144] br[144] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_145 bl[145] br[145] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_146 bl[146] br[146] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_147 bl[147] br[147] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_148 bl[148] br[148] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_149 bl[149] br[149] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_150 bl[150] br[150] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_151 bl[151] br[151] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_152 bl[152] br[152] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_153 bl[153] br[153] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_154 bl[154] br[154] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_155 bl[155] br[155] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_156 bl[156] br[156] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_157 bl[157] br[157] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_158 bl[158] br[158] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_159 bl[159] br[159] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_160 bl[160] br[160] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_161 bl[161] br[161] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_162 bl[162] br[162] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_163 bl[163] br[163] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_164 bl[164] br[164] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_165 bl[165] br[165] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_166 bl[166] br[166] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_167 bl[167] br[167] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_168 bl[168] br[168] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_169 bl[169] br[169] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_170 bl[170] br[170] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_171 bl[171] br[171] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_172 bl[172] br[172] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_173 bl[173] br[173] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_174 bl[174] br[174] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_175 bl[175] br[175] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_176 bl[176] br[176] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_177 bl[177] br[177] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_178 bl[178] br[178] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_179 bl[179] br[179] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_180 bl[180] br[180] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_181 bl[181] br[181] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_182 bl[182] br[182] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_183 bl[183] br[183] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_184 bl[184] br[184] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_185 bl[185] br[185] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_186 bl[186] br[186] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_187 bl[187] br[187] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_188 bl[188] br[188] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_189 bl[189] br[189] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_190 bl[190] br[190] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_191 bl[191] br[191] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_192 bl[192] br[192] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_193 bl[193] br[193] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_194 bl[194] br[194] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_195 bl[195] br[195] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_196 bl[196] br[196] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_197 bl[197] br[197] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_198 bl[198] br[198] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_199 bl[199] br[199] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_200 bl[200] br[200] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_201 bl[201] br[201] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_202 bl[202] br[202] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_203 bl[203] br[203] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_204 bl[204] br[204] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_205 bl[205] br[205] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_206 bl[206] br[206] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_207 bl[207] br[207] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_208 bl[208] br[208] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_209 bl[209] br[209] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_210 bl[210] br[210] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_211 bl[211] br[211] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_212 bl[212] br[212] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_213 bl[213] br[213] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_214 bl[214] br[214] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_215 bl[215] br[215] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_216 bl[216] br[216] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_217 bl[217] br[217] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_218 bl[218] br[218] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_219 bl[219] br[219] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_220 bl[220] br[220] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_221 bl[221] br[221] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_222 bl[222] br[222] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_223 bl[223] br[223] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_224 bl[224] br[224] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_225 bl[225] br[225] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_226 bl[226] br[226] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_227 bl[227] br[227] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_228 bl[228] br[228] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_229 bl[229] br[229] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_230 bl[230] br[230] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_231 bl[231] br[231] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_232 bl[232] br[232] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_233 bl[233] br[233] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_234 bl[234] br[234] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_235 bl[235] br[235] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_236 bl[236] br[236] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_237 bl[237] br[237] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_238 bl[238] br[238] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_239 bl[239] br[239] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_240 bl[240] br[240] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_241 bl[241] br[241] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_242 bl[242] br[242] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_243 bl[243] br[243] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_244 bl[244] br[244] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_245 bl[245] br[245] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_246 bl[246] br[246] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_247 bl[247] br[247] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_248 bl[248] br[248] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_249 bl[249] br[249] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_250 bl[250] br[250] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_251 bl[251] br[251] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_252 bl[252] br[252] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_253 bl[253] br[253] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_254 bl[254] br[254] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_255 bl[255] br[255] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_256 bl[256] br[256] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_257 bl[257] br[257] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_258 bl[258] br[258] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_259 bl[259] br[259] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_260 bl[260] br[260] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_261 bl[261] br[261] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_262 bl[262] br[262] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_263 bl[263] br[263] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_264 bl[264] br[264] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_265 bl[265] br[265] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_266 bl[266] br[266] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_267 bl[267] br[267] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_268 bl[268] br[268] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_269 bl[269] br[269] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_270 bl[270] br[270] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_271 bl[271] br[271] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_272 bl[272] br[272] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_273 bl[273] br[273] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_274 bl[274] br[274] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_275 bl[275] br[275] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_276 bl[276] br[276] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_277 bl[277] br[277] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_278 bl[278] br[278] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_279 bl[279] br[279] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_280 bl[280] br[280] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_281 bl[281] br[281] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_282 bl[282] br[282] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_283 bl[283] br[283] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_284 bl[284] br[284] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_285 bl[285] br[285] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_286 bl[286] br[286] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_287 bl[287] br[287] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_288 bl[288] br[288] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_289 bl[289] br[289] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_290 bl[290] br[290] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_291 bl[291] br[291] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_292 bl[292] br[292] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_293 bl[293] br[293] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_294 bl[294] br[294] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_295 bl[295] br[295] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_296 bl[296] br[296] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_297 bl[297] br[297] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_298 bl[298] br[298] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_299 bl[299] br[299] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_300 bl[300] br[300] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_301 bl[301] br[301] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_302 bl[302] br[302] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_303 bl[303] br[303] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_304 bl[304] br[304] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_305 bl[305] br[305] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_306 bl[306] br[306] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_307 bl[307] br[307] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_308 bl[308] br[308] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_309 bl[309] br[309] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_310 bl[310] br[310] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_311 bl[311] br[311] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_312 bl[312] br[312] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_313 bl[313] br[313] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_314 bl[314] br[314] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_315 bl[315] br[315] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_316 bl[316] br[316] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_317 bl[317] br[317] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_318 bl[318] br[318] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_319 bl[319] br[319] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_320 bl[320] br[320] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_321 bl[321] br[321] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_322 bl[322] br[322] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_323 bl[323] br[323] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_324 bl[324] br[324] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_325 bl[325] br[325] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_326 bl[326] br[326] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_327 bl[327] br[327] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_328 bl[328] br[328] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_329 bl[329] br[329] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_330 bl[330] br[330] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_331 bl[331] br[331] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_332 bl[332] br[332] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_333 bl[333] br[333] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_334 bl[334] br[334] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_335 bl[335] br[335] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_336 bl[336] br[336] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_337 bl[337] br[337] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_338 bl[338] br[338] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_339 bl[339] br[339] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_340 bl[340] br[340] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_341 bl[341] br[341] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_342 bl[342] br[342] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_343 bl[343] br[343] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_344 bl[344] br[344] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_345 bl[345] br[345] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_346 bl[346] br[346] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_347 bl[347] br[347] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_348 bl[348] br[348] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_349 bl[349] br[349] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_350 bl[350] br[350] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_351 bl[351] br[351] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_352 bl[352] br[352] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_353 bl[353] br[353] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_354 bl[354] br[354] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_355 bl[355] br[355] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_356 bl[356] br[356] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_357 bl[357] br[357] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_358 bl[358] br[358] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_359 bl[359] br[359] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_360 bl[360] br[360] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_361 bl[361] br[361] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_362 bl[362] br[362] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_363 bl[363] br[363] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_364 bl[364] br[364] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_365 bl[365] br[365] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_366 bl[366] br[366] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_367 bl[367] br[367] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_368 bl[368] br[368] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_369 bl[369] br[369] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_370 bl[370] br[370] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_371 bl[371] br[371] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_372 bl[372] br[372] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_373 bl[373] br[373] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_374 bl[374] br[374] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_375 bl[375] br[375] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_376 bl[376] br[376] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_377 bl[377] br[377] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_378 bl[378] br[378] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_379 bl[379] br[379] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_380 bl[380] br[380] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_381 bl[381] br[381] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_382 bl[382] br[382] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_383 bl[383] br[383] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_384 bl[384] br[384] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_385 bl[385] br[385] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_386 bl[386] br[386] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_387 bl[387] br[387] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_388 bl[388] br[388] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_389 bl[389] br[389] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_390 bl[390] br[390] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_391 bl[391] br[391] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_392 bl[392] br[392] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_393 bl[393] br[393] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_394 bl[394] br[394] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_395 bl[395] br[395] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_396 bl[396] br[396] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_397 bl[397] br[397] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_398 bl[398] br[398] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_399 bl[399] br[399] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_400 bl[400] br[400] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_401 bl[401] br[401] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_402 bl[402] br[402] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_403 bl[403] br[403] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_404 bl[404] br[404] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_405 bl[405] br[405] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_406 bl[406] br[406] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_407 bl[407] br[407] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_408 bl[408] br[408] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_409 bl[409] br[409] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_410 bl[410] br[410] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_411 bl[411] br[411] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_412 bl[412] br[412] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_413 bl[413] br[413] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_414 bl[414] br[414] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_415 bl[415] br[415] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_416 bl[416] br[416] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_417 bl[417] br[417] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_418 bl[418] br[418] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_419 bl[419] br[419] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_420 bl[420] br[420] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_421 bl[421] br[421] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_422 bl[422] br[422] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_423 bl[423] br[423] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_424 bl[424] br[424] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_425 bl[425] br[425] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_426 bl[426] br[426] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_427 bl[427] br[427] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_428 bl[428] br[428] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_429 bl[429] br[429] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_430 bl[430] br[430] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_431 bl[431] br[431] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_432 bl[432] br[432] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_433 bl[433] br[433] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_434 bl[434] br[434] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_435 bl[435] br[435] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_436 bl[436] br[436] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_437 bl[437] br[437] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_438 bl[438] br[438] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_439 bl[439] br[439] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_440 bl[440] br[440] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_441 bl[441] br[441] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_442 bl[442] br[442] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_443 bl[443] br[443] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_444 bl[444] br[444] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_445 bl[445] br[445] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_446 bl[446] br[446] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_447 bl[447] br[447] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_448 bl[448] br[448] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_449 bl[449] br[449] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_450 bl[450] br[450] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_451 bl[451] br[451] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_452 bl[452] br[452] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_453 bl[453] br[453] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_454 bl[454] br[454] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_455 bl[455] br[455] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_456 bl[456] br[456] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_457 bl[457] br[457] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_458 bl[458] br[458] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_459 bl[459] br[459] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_460 bl[460] br[460] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_461 bl[461] br[461] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_462 bl[462] br[462] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_463 bl[463] br[463] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_464 bl[464] br[464] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_465 bl[465] br[465] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_466 bl[466] br[466] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_467 bl[467] br[467] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_468 bl[468] br[468] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_469 bl[469] br[469] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_470 bl[470] br[470] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_471 bl[471] br[471] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_472 bl[472] br[472] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_473 bl[473] br[473] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_474 bl[474] br[474] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_475 bl[475] br[475] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_476 bl[476] br[476] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_477 bl[477] br[477] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_478 bl[478] br[478] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_479 bl[479] br[479] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_480 bl[480] br[480] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_481 bl[481] br[481] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_482 bl[482] br[482] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_483 bl[483] br[483] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_484 bl[484] br[484] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_485 bl[485] br[485] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_486 bl[486] br[486] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_487 bl[487] br[487] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_488 bl[488] br[488] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_489 bl[489] br[489] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_490 bl[490] br[490] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_491 bl[491] br[491] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_492 bl[492] br[492] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_493 bl[493] br[493] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_494 bl[494] br[494] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_495 bl[495] br[495] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_496 bl[496] br[496] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_497 bl[497] br[497] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_498 bl[498] br[498] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_499 bl[499] br[499] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_500 bl[500] br[500] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_501 bl[501] br[501] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_502 bl[502] br[502] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_503 bl[503] br[503] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_504 bl[504] br[504] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_505 bl[505] br[505] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_506 bl[506] br[506] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_507 bl[507] br[507] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_508 bl[508] br[508] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_509 bl[509] br[509] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_510 bl[510] br[510] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_17_511 bl[511] br[511] vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xcell_18_0 bl[0] br[0] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_1 bl[1] br[1] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_2 bl[2] br[2] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_3 bl[3] br[3] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_4 bl[4] br[4] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_5 bl[5] br[5] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_6 bl[6] br[6] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_7 bl[7] br[7] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_8 bl[8] br[8] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_9 bl[9] br[9] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_10 bl[10] br[10] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_11 bl[11] br[11] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_12 bl[12] br[12] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_13 bl[13] br[13] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_14 bl[14] br[14] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_15 bl[15] br[15] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_16 bl[16] br[16] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_17 bl[17] br[17] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_18 bl[18] br[18] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_19 bl[19] br[19] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_20 bl[20] br[20] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_21 bl[21] br[21] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_22 bl[22] br[22] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_23 bl[23] br[23] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_24 bl[24] br[24] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_25 bl[25] br[25] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_26 bl[26] br[26] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_27 bl[27] br[27] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_28 bl[28] br[28] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_29 bl[29] br[29] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_30 bl[30] br[30] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_31 bl[31] br[31] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_32 bl[32] br[32] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_33 bl[33] br[33] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_34 bl[34] br[34] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_35 bl[35] br[35] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_36 bl[36] br[36] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_37 bl[37] br[37] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_38 bl[38] br[38] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_39 bl[39] br[39] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_40 bl[40] br[40] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_41 bl[41] br[41] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_42 bl[42] br[42] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_43 bl[43] br[43] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_44 bl[44] br[44] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_45 bl[45] br[45] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_46 bl[46] br[46] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_47 bl[47] br[47] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_48 bl[48] br[48] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_49 bl[49] br[49] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_50 bl[50] br[50] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_51 bl[51] br[51] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_52 bl[52] br[52] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_53 bl[53] br[53] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_54 bl[54] br[54] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_55 bl[55] br[55] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_56 bl[56] br[56] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_57 bl[57] br[57] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_58 bl[58] br[58] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_59 bl[59] br[59] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_60 bl[60] br[60] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_61 bl[61] br[61] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_62 bl[62] br[62] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_63 bl[63] br[63] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_64 bl[64] br[64] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_65 bl[65] br[65] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_66 bl[66] br[66] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_67 bl[67] br[67] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_68 bl[68] br[68] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_69 bl[69] br[69] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_70 bl[70] br[70] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_71 bl[71] br[71] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_72 bl[72] br[72] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_73 bl[73] br[73] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_74 bl[74] br[74] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_75 bl[75] br[75] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_76 bl[76] br[76] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_77 bl[77] br[77] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_78 bl[78] br[78] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_79 bl[79] br[79] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_80 bl[80] br[80] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_81 bl[81] br[81] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_82 bl[82] br[82] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_83 bl[83] br[83] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_84 bl[84] br[84] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_85 bl[85] br[85] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_86 bl[86] br[86] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_87 bl[87] br[87] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_88 bl[88] br[88] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_89 bl[89] br[89] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_90 bl[90] br[90] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_91 bl[91] br[91] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_92 bl[92] br[92] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_93 bl[93] br[93] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_94 bl[94] br[94] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_95 bl[95] br[95] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_96 bl[96] br[96] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_97 bl[97] br[97] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_98 bl[98] br[98] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_99 bl[99] br[99] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_100 bl[100] br[100] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_101 bl[101] br[101] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_102 bl[102] br[102] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_103 bl[103] br[103] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_104 bl[104] br[104] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_105 bl[105] br[105] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_106 bl[106] br[106] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_107 bl[107] br[107] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_108 bl[108] br[108] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_109 bl[109] br[109] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_110 bl[110] br[110] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_111 bl[111] br[111] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_112 bl[112] br[112] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_113 bl[113] br[113] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_114 bl[114] br[114] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_115 bl[115] br[115] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_116 bl[116] br[116] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_117 bl[117] br[117] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_118 bl[118] br[118] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_119 bl[119] br[119] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_120 bl[120] br[120] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_121 bl[121] br[121] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_122 bl[122] br[122] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_123 bl[123] br[123] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_124 bl[124] br[124] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_125 bl[125] br[125] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_126 bl[126] br[126] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_127 bl[127] br[127] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_128 bl[128] br[128] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_129 bl[129] br[129] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_130 bl[130] br[130] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_131 bl[131] br[131] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_132 bl[132] br[132] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_133 bl[133] br[133] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_134 bl[134] br[134] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_135 bl[135] br[135] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_136 bl[136] br[136] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_137 bl[137] br[137] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_138 bl[138] br[138] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_139 bl[139] br[139] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_140 bl[140] br[140] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_141 bl[141] br[141] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_142 bl[142] br[142] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_143 bl[143] br[143] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_144 bl[144] br[144] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_145 bl[145] br[145] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_146 bl[146] br[146] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_147 bl[147] br[147] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_148 bl[148] br[148] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_149 bl[149] br[149] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_150 bl[150] br[150] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_151 bl[151] br[151] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_152 bl[152] br[152] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_153 bl[153] br[153] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_154 bl[154] br[154] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_155 bl[155] br[155] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_156 bl[156] br[156] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_157 bl[157] br[157] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_158 bl[158] br[158] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_159 bl[159] br[159] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_160 bl[160] br[160] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_161 bl[161] br[161] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_162 bl[162] br[162] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_163 bl[163] br[163] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_164 bl[164] br[164] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_165 bl[165] br[165] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_166 bl[166] br[166] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_167 bl[167] br[167] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_168 bl[168] br[168] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_169 bl[169] br[169] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_170 bl[170] br[170] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_171 bl[171] br[171] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_172 bl[172] br[172] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_173 bl[173] br[173] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_174 bl[174] br[174] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_175 bl[175] br[175] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_176 bl[176] br[176] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_177 bl[177] br[177] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_178 bl[178] br[178] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_179 bl[179] br[179] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_180 bl[180] br[180] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_181 bl[181] br[181] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_182 bl[182] br[182] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_183 bl[183] br[183] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_184 bl[184] br[184] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_185 bl[185] br[185] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_186 bl[186] br[186] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_187 bl[187] br[187] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_188 bl[188] br[188] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_189 bl[189] br[189] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_190 bl[190] br[190] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_191 bl[191] br[191] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_192 bl[192] br[192] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_193 bl[193] br[193] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_194 bl[194] br[194] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_195 bl[195] br[195] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_196 bl[196] br[196] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_197 bl[197] br[197] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_198 bl[198] br[198] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_199 bl[199] br[199] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_200 bl[200] br[200] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_201 bl[201] br[201] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_202 bl[202] br[202] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_203 bl[203] br[203] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_204 bl[204] br[204] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_205 bl[205] br[205] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_206 bl[206] br[206] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_207 bl[207] br[207] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_208 bl[208] br[208] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_209 bl[209] br[209] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_210 bl[210] br[210] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_211 bl[211] br[211] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_212 bl[212] br[212] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_213 bl[213] br[213] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_214 bl[214] br[214] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_215 bl[215] br[215] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_216 bl[216] br[216] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_217 bl[217] br[217] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_218 bl[218] br[218] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_219 bl[219] br[219] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_220 bl[220] br[220] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_221 bl[221] br[221] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_222 bl[222] br[222] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_223 bl[223] br[223] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_224 bl[224] br[224] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_225 bl[225] br[225] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_226 bl[226] br[226] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_227 bl[227] br[227] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_228 bl[228] br[228] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_229 bl[229] br[229] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_230 bl[230] br[230] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_231 bl[231] br[231] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_232 bl[232] br[232] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_233 bl[233] br[233] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_234 bl[234] br[234] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_235 bl[235] br[235] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_236 bl[236] br[236] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_237 bl[237] br[237] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_238 bl[238] br[238] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_239 bl[239] br[239] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_240 bl[240] br[240] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_241 bl[241] br[241] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_242 bl[242] br[242] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_243 bl[243] br[243] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_244 bl[244] br[244] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_245 bl[245] br[245] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_246 bl[246] br[246] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_247 bl[247] br[247] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_248 bl[248] br[248] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_249 bl[249] br[249] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_250 bl[250] br[250] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_251 bl[251] br[251] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_252 bl[252] br[252] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_253 bl[253] br[253] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_254 bl[254] br[254] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_255 bl[255] br[255] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_256 bl[256] br[256] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_257 bl[257] br[257] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_258 bl[258] br[258] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_259 bl[259] br[259] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_260 bl[260] br[260] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_261 bl[261] br[261] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_262 bl[262] br[262] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_263 bl[263] br[263] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_264 bl[264] br[264] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_265 bl[265] br[265] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_266 bl[266] br[266] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_267 bl[267] br[267] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_268 bl[268] br[268] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_269 bl[269] br[269] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_270 bl[270] br[270] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_271 bl[271] br[271] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_272 bl[272] br[272] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_273 bl[273] br[273] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_274 bl[274] br[274] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_275 bl[275] br[275] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_276 bl[276] br[276] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_277 bl[277] br[277] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_278 bl[278] br[278] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_279 bl[279] br[279] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_280 bl[280] br[280] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_281 bl[281] br[281] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_282 bl[282] br[282] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_283 bl[283] br[283] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_284 bl[284] br[284] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_285 bl[285] br[285] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_286 bl[286] br[286] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_287 bl[287] br[287] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_288 bl[288] br[288] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_289 bl[289] br[289] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_290 bl[290] br[290] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_291 bl[291] br[291] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_292 bl[292] br[292] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_293 bl[293] br[293] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_294 bl[294] br[294] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_295 bl[295] br[295] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_296 bl[296] br[296] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_297 bl[297] br[297] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_298 bl[298] br[298] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_299 bl[299] br[299] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_300 bl[300] br[300] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_301 bl[301] br[301] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_302 bl[302] br[302] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_303 bl[303] br[303] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_304 bl[304] br[304] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_305 bl[305] br[305] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_306 bl[306] br[306] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_307 bl[307] br[307] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_308 bl[308] br[308] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_309 bl[309] br[309] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_310 bl[310] br[310] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_311 bl[311] br[311] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_312 bl[312] br[312] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_313 bl[313] br[313] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_314 bl[314] br[314] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_315 bl[315] br[315] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_316 bl[316] br[316] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_317 bl[317] br[317] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_318 bl[318] br[318] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_319 bl[319] br[319] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_320 bl[320] br[320] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_321 bl[321] br[321] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_322 bl[322] br[322] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_323 bl[323] br[323] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_324 bl[324] br[324] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_325 bl[325] br[325] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_326 bl[326] br[326] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_327 bl[327] br[327] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_328 bl[328] br[328] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_329 bl[329] br[329] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_330 bl[330] br[330] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_331 bl[331] br[331] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_332 bl[332] br[332] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_333 bl[333] br[333] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_334 bl[334] br[334] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_335 bl[335] br[335] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_336 bl[336] br[336] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_337 bl[337] br[337] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_338 bl[338] br[338] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_339 bl[339] br[339] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_340 bl[340] br[340] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_341 bl[341] br[341] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_342 bl[342] br[342] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_343 bl[343] br[343] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_344 bl[344] br[344] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_345 bl[345] br[345] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_346 bl[346] br[346] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_347 bl[347] br[347] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_348 bl[348] br[348] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_349 bl[349] br[349] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_350 bl[350] br[350] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_351 bl[351] br[351] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_352 bl[352] br[352] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_353 bl[353] br[353] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_354 bl[354] br[354] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_355 bl[355] br[355] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_356 bl[356] br[356] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_357 bl[357] br[357] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_358 bl[358] br[358] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_359 bl[359] br[359] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_360 bl[360] br[360] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_361 bl[361] br[361] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_362 bl[362] br[362] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_363 bl[363] br[363] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_364 bl[364] br[364] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_365 bl[365] br[365] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_366 bl[366] br[366] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_367 bl[367] br[367] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_368 bl[368] br[368] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_369 bl[369] br[369] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_370 bl[370] br[370] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_371 bl[371] br[371] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_372 bl[372] br[372] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_373 bl[373] br[373] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_374 bl[374] br[374] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_375 bl[375] br[375] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_376 bl[376] br[376] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_377 bl[377] br[377] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_378 bl[378] br[378] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_379 bl[379] br[379] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_380 bl[380] br[380] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_381 bl[381] br[381] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_382 bl[382] br[382] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_383 bl[383] br[383] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_384 bl[384] br[384] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_385 bl[385] br[385] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_386 bl[386] br[386] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_387 bl[387] br[387] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_388 bl[388] br[388] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_389 bl[389] br[389] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_390 bl[390] br[390] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_391 bl[391] br[391] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_392 bl[392] br[392] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_393 bl[393] br[393] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_394 bl[394] br[394] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_395 bl[395] br[395] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_396 bl[396] br[396] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_397 bl[397] br[397] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_398 bl[398] br[398] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_399 bl[399] br[399] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_400 bl[400] br[400] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_401 bl[401] br[401] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_402 bl[402] br[402] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_403 bl[403] br[403] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_404 bl[404] br[404] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_405 bl[405] br[405] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_406 bl[406] br[406] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_407 bl[407] br[407] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_408 bl[408] br[408] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_409 bl[409] br[409] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_410 bl[410] br[410] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_411 bl[411] br[411] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_412 bl[412] br[412] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_413 bl[413] br[413] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_414 bl[414] br[414] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_415 bl[415] br[415] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_416 bl[416] br[416] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_417 bl[417] br[417] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_418 bl[418] br[418] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_419 bl[419] br[419] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_420 bl[420] br[420] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_421 bl[421] br[421] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_422 bl[422] br[422] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_423 bl[423] br[423] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_424 bl[424] br[424] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_425 bl[425] br[425] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_426 bl[426] br[426] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_427 bl[427] br[427] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_428 bl[428] br[428] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_429 bl[429] br[429] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_430 bl[430] br[430] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_431 bl[431] br[431] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_432 bl[432] br[432] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_433 bl[433] br[433] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_434 bl[434] br[434] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_435 bl[435] br[435] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_436 bl[436] br[436] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_437 bl[437] br[437] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_438 bl[438] br[438] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_439 bl[439] br[439] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_440 bl[440] br[440] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_441 bl[441] br[441] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_442 bl[442] br[442] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_443 bl[443] br[443] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_444 bl[444] br[444] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_445 bl[445] br[445] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_446 bl[446] br[446] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_447 bl[447] br[447] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_448 bl[448] br[448] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_449 bl[449] br[449] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_450 bl[450] br[450] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_451 bl[451] br[451] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_452 bl[452] br[452] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_453 bl[453] br[453] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_454 bl[454] br[454] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_455 bl[455] br[455] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_456 bl[456] br[456] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_457 bl[457] br[457] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_458 bl[458] br[458] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_459 bl[459] br[459] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_460 bl[460] br[460] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_461 bl[461] br[461] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_462 bl[462] br[462] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_463 bl[463] br[463] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_464 bl[464] br[464] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_465 bl[465] br[465] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_466 bl[466] br[466] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_467 bl[467] br[467] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_468 bl[468] br[468] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_469 bl[469] br[469] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_470 bl[470] br[470] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_471 bl[471] br[471] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_472 bl[472] br[472] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_473 bl[473] br[473] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_474 bl[474] br[474] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_475 bl[475] br[475] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_476 bl[476] br[476] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_477 bl[477] br[477] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_478 bl[478] br[478] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_479 bl[479] br[479] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_480 bl[480] br[480] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_481 bl[481] br[481] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_482 bl[482] br[482] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_483 bl[483] br[483] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_484 bl[484] br[484] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_485 bl[485] br[485] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_486 bl[486] br[486] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_487 bl[487] br[487] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_488 bl[488] br[488] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_489 bl[489] br[489] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_490 bl[490] br[490] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_491 bl[491] br[491] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_492 bl[492] br[492] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_493 bl[493] br[493] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_494 bl[494] br[494] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_495 bl[495] br[495] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_496 bl[496] br[496] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_497 bl[497] br[497] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_498 bl[498] br[498] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_499 bl[499] br[499] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_500 bl[500] br[500] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_501 bl[501] br[501] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_502 bl[502] br[502] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_503 bl[503] br[503] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_504 bl[504] br[504] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_505 bl[505] br[505] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_506 bl[506] br[506] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_507 bl[507] br[507] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_508 bl[508] br[508] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_509 bl[509] br[509] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_510 bl[510] br[510] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_18_511 bl[511] br[511] vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xcell_19_0 bl[0] br[0] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_1 bl[1] br[1] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_2 bl[2] br[2] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_3 bl[3] br[3] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_4 bl[4] br[4] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_5 bl[5] br[5] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_6 bl[6] br[6] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_7 bl[7] br[7] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_8 bl[8] br[8] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_9 bl[9] br[9] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_10 bl[10] br[10] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_11 bl[11] br[11] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_12 bl[12] br[12] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_13 bl[13] br[13] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_14 bl[14] br[14] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_15 bl[15] br[15] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_16 bl[16] br[16] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_17 bl[17] br[17] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_18 bl[18] br[18] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_19 bl[19] br[19] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_20 bl[20] br[20] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_21 bl[21] br[21] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_22 bl[22] br[22] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_23 bl[23] br[23] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_24 bl[24] br[24] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_25 bl[25] br[25] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_26 bl[26] br[26] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_27 bl[27] br[27] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_28 bl[28] br[28] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_29 bl[29] br[29] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_30 bl[30] br[30] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_31 bl[31] br[31] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_32 bl[32] br[32] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_33 bl[33] br[33] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_34 bl[34] br[34] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_35 bl[35] br[35] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_36 bl[36] br[36] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_37 bl[37] br[37] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_38 bl[38] br[38] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_39 bl[39] br[39] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_40 bl[40] br[40] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_41 bl[41] br[41] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_42 bl[42] br[42] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_43 bl[43] br[43] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_44 bl[44] br[44] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_45 bl[45] br[45] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_46 bl[46] br[46] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_47 bl[47] br[47] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_48 bl[48] br[48] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_49 bl[49] br[49] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_50 bl[50] br[50] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_51 bl[51] br[51] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_52 bl[52] br[52] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_53 bl[53] br[53] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_54 bl[54] br[54] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_55 bl[55] br[55] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_56 bl[56] br[56] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_57 bl[57] br[57] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_58 bl[58] br[58] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_59 bl[59] br[59] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_60 bl[60] br[60] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_61 bl[61] br[61] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_62 bl[62] br[62] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_63 bl[63] br[63] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_64 bl[64] br[64] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_65 bl[65] br[65] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_66 bl[66] br[66] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_67 bl[67] br[67] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_68 bl[68] br[68] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_69 bl[69] br[69] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_70 bl[70] br[70] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_71 bl[71] br[71] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_72 bl[72] br[72] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_73 bl[73] br[73] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_74 bl[74] br[74] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_75 bl[75] br[75] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_76 bl[76] br[76] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_77 bl[77] br[77] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_78 bl[78] br[78] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_79 bl[79] br[79] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_80 bl[80] br[80] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_81 bl[81] br[81] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_82 bl[82] br[82] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_83 bl[83] br[83] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_84 bl[84] br[84] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_85 bl[85] br[85] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_86 bl[86] br[86] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_87 bl[87] br[87] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_88 bl[88] br[88] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_89 bl[89] br[89] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_90 bl[90] br[90] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_91 bl[91] br[91] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_92 bl[92] br[92] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_93 bl[93] br[93] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_94 bl[94] br[94] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_95 bl[95] br[95] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_96 bl[96] br[96] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_97 bl[97] br[97] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_98 bl[98] br[98] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_99 bl[99] br[99] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_100 bl[100] br[100] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_101 bl[101] br[101] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_102 bl[102] br[102] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_103 bl[103] br[103] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_104 bl[104] br[104] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_105 bl[105] br[105] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_106 bl[106] br[106] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_107 bl[107] br[107] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_108 bl[108] br[108] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_109 bl[109] br[109] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_110 bl[110] br[110] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_111 bl[111] br[111] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_112 bl[112] br[112] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_113 bl[113] br[113] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_114 bl[114] br[114] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_115 bl[115] br[115] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_116 bl[116] br[116] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_117 bl[117] br[117] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_118 bl[118] br[118] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_119 bl[119] br[119] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_120 bl[120] br[120] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_121 bl[121] br[121] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_122 bl[122] br[122] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_123 bl[123] br[123] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_124 bl[124] br[124] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_125 bl[125] br[125] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_126 bl[126] br[126] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_127 bl[127] br[127] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_128 bl[128] br[128] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_129 bl[129] br[129] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_130 bl[130] br[130] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_131 bl[131] br[131] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_132 bl[132] br[132] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_133 bl[133] br[133] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_134 bl[134] br[134] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_135 bl[135] br[135] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_136 bl[136] br[136] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_137 bl[137] br[137] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_138 bl[138] br[138] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_139 bl[139] br[139] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_140 bl[140] br[140] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_141 bl[141] br[141] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_142 bl[142] br[142] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_143 bl[143] br[143] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_144 bl[144] br[144] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_145 bl[145] br[145] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_146 bl[146] br[146] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_147 bl[147] br[147] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_148 bl[148] br[148] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_149 bl[149] br[149] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_150 bl[150] br[150] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_151 bl[151] br[151] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_152 bl[152] br[152] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_153 bl[153] br[153] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_154 bl[154] br[154] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_155 bl[155] br[155] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_156 bl[156] br[156] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_157 bl[157] br[157] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_158 bl[158] br[158] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_159 bl[159] br[159] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_160 bl[160] br[160] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_161 bl[161] br[161] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_162 bl[162] br[162] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_163 bl[163] br[163] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_164 bl[164] br[164] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_165 bl[165] br[165] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_166 bl[166] br[166] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_167 bl[167] br[167] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_168 bl[168] br[168] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_169 bl[169] br[169] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_170 bl[170] br[170] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_171 bl[171] br[171] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_172 bl[172] br[172] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_173 bl[173] br[173] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_174 bl[174] br[174] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_175 bl[175] br[175] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_176 bl[176] br[176] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_177 bl[177] br[177] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_178 bl[178] br[178] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_179 bl[179] br[179] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_180 bl[180] br[180] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_181 bl[181] br[181] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_182 bl[182] br[182] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_183 bl[183] br[183] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_184 bl[184] br[184] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_185 bl[185] br[185] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_186 bl[186] br[186] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_187 bl[187] br[187] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_188 bl[188] br[188] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_189 bl[189] br[189] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_190 bl[190] br[190] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_191 bl[191] br[191] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_192 bl[192] br[192] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_193 bl[193] br[193] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_194 bl[194] br[194] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_195 bl[195] br[195] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_196 bl[196] br[196] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_197 bl[197] br[197] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_198 bl[198] br[198] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_199 bl[199] br[199] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_200 bl[200] br[200] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_201 bl[201] br[201] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_202 bl[202] br[202] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_203 bl[203] br[203] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_204 bl[204] br[204] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_205 bl[205] br[205] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_206 bl[206] br[206] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_207 bl[207] br[207] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_208 bl[208] br[208] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_209 bl[209] br[209] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_210 bl[210] br[210] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_211 bl[211] br[211] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_212 bl[212] br[212] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_213 bl[213] br[213] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_214 bl[214] br[214] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_215 bl[215] br[215] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_216 bl[216] br[216] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_217 bl[217] br[217] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_218 bl[218] br[218] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_219 bl[219] br[219] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_220 bl[220] br[220] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_221 bl[221] br[221] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_222 bl[222] br[222] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_223 bl[223] br[223] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_224 bl[224] br[224] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_225 bl[225] br[225] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_226 bl[226] br[226] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_227 bl[227] br[227] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_228 bl[228] br[228] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_229 bl[229] br[229] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_230 bl[230] br[230] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_231 bl[231] br[231] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_232 bl[232] br[232] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_233 bl[233] br[233] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_234 bl[234] br[234] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_235 bl[235] br[235] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_236 bl[236] br[236] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_237 bl[237] br[237] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_238 bl[238] br[238] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_239 bl[239] br[239] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_240 bl[240] br[240] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_241 bl[241] br[241] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_242 bl[242] br[242] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_243 bl[243] br[243] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_244 bl[244] br[244] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_245 bl[245] br[245] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_246 bl[246] br[246] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_247 bl[247] br[247] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_248 bl[248] br[248] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_249 bl[249] br[249] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_250 bl[250] br[250] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_251 bl[251] br[251] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_252 bl[252] br[252] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_253 bl[253] br[253] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_254 bl[254] br[254] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_255 bl[255] br[255] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_256 bl[256] br[256] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_257 bl[257] br[257] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_258 bl[258] br[258] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_259 bl[259] br[259] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_260 bl[260] br[260] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_261 bl[261] br[261] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_262 bl[262] br[262] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_263 bl[263] br[263] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_264 bl[264] br[264] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_265 bl[265] br[265] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_266 bl[266] br[266] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_267 bl[267] br[267] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_268 bl[268] br[268] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_269 bl[269] br[269] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_270 bl[270] br[270] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_271 bl[271] br[271] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_272 bl[272] br[272] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_273 bl[273] br[273] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_274 bl[274] br[274] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_275 bl[275] br[275] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_276 bl[276] br[276] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_277 bl[277] br[277] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_278 bl[278] br[278] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_279 bl[279] br[279] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_280 bl[280] br[280] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_281 bl[281] br[281] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_282 bl[282] br[282] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_283 bl[283] br[283] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_284 bl[284] br[284] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_285 bl[285] br[285] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_286 bl[286] br[286] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_287 bl[287] br[287] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_288 bl[288] br[288] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_289 bl[289] br[289] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_290 bl[290] br[290] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_291 bl[291] br[291] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_292 bl[292] br[292] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_293 bl[293] br[293] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_294 bl[294] br[294] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_295 bl[295] br[295] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_296 bl[296] br[296] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_297 bl[297] br[297] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_298 bl[298] br[298] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_299 bl[299] br[299] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_300 bl[300] br[300] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_301 bl[301] br[301] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_302 bl[302] br[302] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_303 bl[303] br[303] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_304 bl[304] br[304] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_305 bl[305] br[305] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_306 bl[306] br[306] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_307 bl[307] br[307] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_308 bl[308] br[308] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_309 bl[309] br[309] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_310 bl[310] br[310] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_311 bl[311] br[311] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_312 bl[312] br[312] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_313 bl[313] br[313] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_314 bl[314] br[314] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_315 bl[315] br[315] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_316 bl[316] br[316] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_317 bl[317] br[317] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_318 bl[318] br[318] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_319 bl[319] br[319] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_320 bl[320] br[320] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_321 bl[321] br[321] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_322 bl[322] br[322] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_323 bl[323] br[323] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_324 bl[324] br[324] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_325 bl[325] br[325] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_326 bl[326] br[326] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_327 bl[327] br[327] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_328 bl[328] br[328] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_329 bl[329] br[329] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_330 bl[330] br[330] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_331 bl[331] br[331] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_332 bl[332] br[332] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_333 bl[333] br[333] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_334 bl[334] br[334] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_335 bl[335] br[335] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_336 bl[336] br[336] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_337 bl[337] br[337] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_338 bl[338] br[338] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_339 bl[339] br[339] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_340 bl[340] br[340] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_341 bl[341] br[341] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_342 bl[342] br[342] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_343 bl[343] br[343] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_344 bl[344] br[344] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_345 bl[345] br[345] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_346 bl[346] br[346] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_347 bl[347] br[347] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_348 bl[348] br[348] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_349 bl[349] br[349] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_350 bl[350] br[350] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_351 bl[351] br[351] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_352 bl[352] br[352] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_353 bl[353] br[353] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_354 bl[354] br[354] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_355 bl[355] br[355] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_356 bl[356] br[356] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_357 bl[357] br[357] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_358 bl[358] br[358] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_359 bl[359] br[359] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_360 bl[360] br[360] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_361 bl[361] br[361] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_362 bl[362] br[362] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_363 bl[363] br[363] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_364 bl[364] br[364] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_365 bl[365] br[365] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_366 bl[366] br[366] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_367 bl[367] br[367] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_368 bl[368] br[368] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_369 bl[369] br[369] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_370 bl[370] br[370] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_371 bl[371] br[371] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_372 bl[372] br[372] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_373 bl[373] br[373] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_374 bl[374] br[374] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_375 bl[375] br[375] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_376 bl[376] br[376] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_377 bl[377] br[377] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_378 bl[378] br[378] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_379 bl[379] br[379] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_380 bl[380] br[380] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_381 bl[381] br[381] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_382 bl[382] br[382] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_383 bl[383] br[383] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_384 bl[384] br[384] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_385 bl[385] br[385] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_386 bl[386] br[386] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_387 bl[387] br[387] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_388 bl[388] br[388] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_389 bl[389] br[389] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_390 bl[390] br[390] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_391 bl[391] br[391] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_392 bl[392] br[392] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_393 bl[393] br[393] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_394 bl[394] br[394] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_395 bl[395] br[395] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_396 bl[396] br[396] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_397 bl[397] br[397] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_398 bl[398] br[398] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_399 bl[399] br[399] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_400 bl[400] br[400] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_401 bl[401] br[401] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_402 bl[402] br[402] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_403 bl[403] br[403] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_404 bl[404] br[404] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_405 bl[405] br[405] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_406 bl[406] br[406] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_407 bl[407] br[407] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_408 bl[408] br[408] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_409 bl[409] br[409] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_410 bl[410] br[410] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_411 bl[411] br[411] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_412 bl[412] br[412] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_413 bl[413] br[413] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_414 bl[414] br[414] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_415 bl[415] br[415] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_416 bl[416] br[416] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_417 bl[417] br[417] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_418 bl[418] br[418] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_419 bl[419] br[419] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_420 bl[420] br[420] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_421 bl[421] br[421] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_422 bl[422] br[422] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_423 bl[423] br[423] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_424 bl[424] br[424] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_425 bl[425] br[425] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_426 bl[426] br[426] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_427 bl[427] br[427] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_428 bl[428] br[428] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_429 bl[429] br[429] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_430 bl[430] br[430] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_431 bl[431] br[431] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_432 bl[432] br[432] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_433 bl[433] br[433] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_434 bl[434] br[434] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_435 bl[435] br[435] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_436 bl[436] br[436] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_437 bl[437] br[437] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_438 bl[438] br[438] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_439 bl[439] br[439] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_440 bl[440] br[440] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_441 bl[441] br[441] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_442 bl[442] br[442] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_443 bl[443] br[443] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_444 bl[444] br[444] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_445 bl[445] br[445] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_446 bl[446] br[446] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_447 bl[447] br[447] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_448 bl[448] br[448] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_449 bl[449] br[449] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_450 bl[450] br[450] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_451 bl[451] br[451] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_452 bl[452] br[452] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_453 bl[453] br[453] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_454 bl[454] br[454] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_455 bl[455] br[455] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_456 bl[456] br[456] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_457 bl[457] br[457] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_458 bl[458] br[458] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_459 bl[459] br[459] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_460 bl[460] br[460] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_461 bl[461] br[461] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_462 bl[462] br[462] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_463 bl[463] br[463] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_464 bl[464] br[464] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_465 bl[465] br[465] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_466 bl[466] br[466] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_467 bl[467] br[467] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_468 bl[468] br[468] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_469 bl[469] br[469] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_470 bl[470] br[470] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_471 bl[471] br[471] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_472 bl[472] br[472] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_473 bl[473] br[473] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_474 bl[474] br[474] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_475 bl[475] br[475] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_476 bl[476] br[476] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_477 bl[477] br[477] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_478 bl[478] br[478] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_479 bl[479] br[479] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_480 bl[480] br[480] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_481 bl[481] br[481] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_482 bl[482] br[482] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_483 bl[483] br[483] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_484 bl[484] br[484] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_485 bl[485] br[485] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_486 bl[486] br[486] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_487 bl[487] br[487] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_488 bl[488] br[488] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_489 bl[489] br[489] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_490 bl[490] br[490] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_491 bl[491] br[491] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_492 bl[492] br[492] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_493 bl[493] br[493] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_494 bl[494] br[494] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_495 bl[495] br[495] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_496 bl[496] br[496] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_497 bl[497] br[497] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_498 bl[498] br[498] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_499 bl[499] br[499] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_500 bl[500] br[500] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_501 bl[501] br[501] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_502 bl[502] br[502] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_503 bl[503] br[503] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_504 bl[504] br[504] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_505 bl[505] br[505] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_506 bl[506] br[506] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_507 bl[507] br[507] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_508 bl[508] br[508] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_509 bl[509] br[509] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_510 bl[510] br[510] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_19_511 bl[511] br[511] vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xcell_20_0 bl[0] br[0] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_1 bl[1] br[1] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_2 bl[2] br[2] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_3 bl[3] br[3] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_4 bl[4] br[4] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_5 bl[5] br[5] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_6 bl[6] br[6] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_7 bl[7] br[7] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_8 bl[8] br[8] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_9 bl[9] br[9] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_10 bl[10] br[10] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_11 bl[11] br[11] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_12 bl[12] br[12] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_13 bl[13] br[13] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_14 bl[14] br[14] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_15 bl[15] br[15] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_16 bl[16] br[16] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_17 bl[17] br[17] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_18 bl[18] br[18] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_19 bl[19] br[19] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_20 bl[20] br[20] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_21 bl[21] br[21] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_22 bl[22] br[22] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_23 bl[23] br[23] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_24 bl[24] br[24] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_25 bl[25] br[25] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_26 bl[26] br[26] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_27 bl[27] br[27] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_28 bl[28] br[28] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_29 bl[29] br[29] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_30 bl[30] br[30] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_31 bl[31] br[31] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_32 bl[32] br[32] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_33 bl[33] br[33] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_34 bl[34] br[34] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_35 bl[35] br[35] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_36 bl[36] br[36] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_37 bl[37] br[37] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_38 bl[38] br[38] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_39 bl[39] br[39] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_40 bl[40] br[40] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_41 bl[41] br[41] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_42 bl[42] br[42] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_43 bl[43] br[43] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_44 bl[44] br[44] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_45 bl[45] br[45] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_46 bl[46] br[46] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_47 bl[47] br[47] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_48 bl[48] br[48] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_49 bl[49] br[49] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_50 bl[50] br[50] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_51 bl[51] br[51] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_52 bl[52] br[52] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_53 bl[53] br[53] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_54 bl[54] br[54] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_55 bl[55] br[55] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_56 bl[56] br[56] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_57 bl[57] br[57] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_58 bl[58] br[58] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_59 bl[59] br[59] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_60 bl[60] br[60] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_61 bl[61] br[61] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_62 bl[62] br[62] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_63 bl[63] br[63] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_64 bl[64] br[64] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_65 bl[65] br[65] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_66 bl[66] br[66] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_67 bl[67] br[67] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_68 bl[68] br[68] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_69 bl[69] br[69] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_70 bl[70] br[70] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_71 bl[71] br[71] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_72 bl[72] br[72] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_73 bl[73] br[73] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_74 bl[74] br[74] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_75 bl[75] br[75] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_76 bl[76] br[76] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_77 bl[77] br[77] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_78 bl[78] br[78] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_79 bl[79] br[79] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_80 bl[80] br[80] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_81 bl[81] br[81] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_82 bl[82] br[82] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_83 bl[83] br[83] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_84 bl[84] br[84] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_85 bl[85] br[85] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_86 bl[86] br[86] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_87 bl[87] br[87] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_88 bl[88] br[88] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_89 bl[89] br[89] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_90 bl[90] br[90] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_91 bl[91] br[91] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_92 bl[92] br[92] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_93 bl[93] br[93] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_94 bl[94] br[94] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_95 bl[95] br[95] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_96 bl[96] br[96] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_97 bl[97] br[97] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_98 bl[98] br[98] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_99 bl[99] br[99] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_100 bl[100] br[100] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_101 bl[101] br[101] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_102 bl[102] br[102] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_103 bl[103] br[103] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_104 bl[104] br[104] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_105 bl[105] br[105] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_106 bl[106] br[106] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_107 bl[107] br[107] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_108 bl[108] br[108] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_109 bl[109] br[109] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_110 bl[110] br[110] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_111 bl[111] br[111] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_112 bl[112] br[112] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_113 bl[113] br[113] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_114 bl[114] br[114] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_115 bl[115] br[115] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_116 bl[116] br[116] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_117 bl[117] br[117] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_118 bl[118] br[118] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_119 bl[119] br[119] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_120 bl[120] br[120] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_121 bl[121] br[121] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_122 bl[122] br[122] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_123 bl[123] br[123] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_124 bl[124] br[124] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_125 bl[125] br[125] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_126 bl[126] br[126] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_127 bl[127] br[127] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_128 bl[128] br[128] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_129 bl[129] br[129] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_130 bl[130] br[130] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_131 bl[131] br[131] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_132 bl[132] br[132] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_133 bl[133] br[133] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_134 bl[134] br[134] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_135 bl[135] br[135] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_136 bl[136] br[136] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_137 bl[137] br[137] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_138 bl[138] br[138] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_139 bl[139] br[139] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_140 bl[140] br[140] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_141 bl[141] br[141] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_142 bl[142] br[142] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_143 bl[143] br[143] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_144 bl[144] br[144] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_145 bl[145] br[145] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_146 bl[146] br[146] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_147 bl[147] br[147] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_148 bl[148] br[148] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_149 bl[149] br[149] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_150 bl[150] br[150] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_151 bl[151] br[151] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_152 bl[152] br[152] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_153 bl[153] br[153] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_154 bl[154] br[154] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_155 bl[155] br[155] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_156 bl[156] br[156] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_157 bl[157] br[157] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_158 bl[158] br[158] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_159 bl[159] br[159] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_160 bl[160] br[160] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_161 bl[161] br[161] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_162 bl[162] br[162] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_163 bl[163] br[163] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_164 bl[164] br[164] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_165 bl[165] br[165] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_166 bl[166] br[166] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_167 bl[167] br[167] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_168 bl[168] br[168] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_169 bl[169] br[169] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_170 bl[170] br[170] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_171 bl[171] br[171] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_172 bl[172] br[172] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_173 bl[173] br[173] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_174 bl[174] br[174] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_175 bl[175] br[175] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_176 bl[176] br[176] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_177 bl[177] br[177] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_178 bl[178] br[178] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_179 bl[179] br[179] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_180 bl[180] br[180] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_181 bl[181] br[181] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_182 bl[182] br[182] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_183 bl[183] br[183] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_184 bl[184] br[184] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_185 bl[185] br[185] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_186 bl[186] br[186] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_187 bl[187] br[187] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_188 bl[188] br[188] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_189 bl[189] br[189] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_190 bl[190] br[190] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_191 bl[191] br[191] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_192 bl[192] br[192] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_193 bl[193] br[193] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_194 bl[194] br[194] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_195 bl[195] br[195] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_196 bl[196] br[196] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_197 bl[197] br[197] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_198 bl[198] br[198] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_199 bl[199] br[199] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_200 bl[200] br[200] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_201 bl[201] br[201] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_202 bl[202] br[202] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_203 bl[203] br[203] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_204 bl[204] br[204] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_205 bl[205] br[205] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_206 bl[206] br[206] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_207 bl[207] br[207] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_208 bl[208] br[208] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_209 bl[209] br[209] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_210 bl[210] br[210] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_211 bl[211] br[211] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_212 bl[212] br[212] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_213 bl[213] br[213] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_214 bl[214] br[214] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_215 bl[215] br[215] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_216 bl[216] br[216] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_217 bl[217] br[217] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_218 bl[218] br[218] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_219 bl[219] br[219] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_220 bl[220] br[220] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_221 bl[221] br[221] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_222 bl[222] br[222] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_223 bl[223] br[223] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_224 bl[224] br[224] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_225 bl[225] br[225] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_226 bl[226] br[226] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_227 bl[227] br[227] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_228 bl[228] br[228] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_229 bl[229] br[229] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_230 bl[230] br[230] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_231 bl[231] br[231] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_232 bl[232] br[232] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_233 bl[233] br[233] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_234 bl[234] br[234] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_235 bl[235] br[235] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_236 bl[236] br[236] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_237 bl[237] br[237] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_238 bl[238] br[238] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_239 bl[239] br[239] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_240 bl[240] br[240] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_241 bl[241] br[241] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_242 bl[242] br[242] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_243 bl[243] br[243] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_244 bl[244] br[244] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_245 bl[245] br[245] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_246 bl[246] br[246] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_247 bl[247] br[247] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_248 bl[248] br[248] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_249 bl[249] br[249] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_250 bl[250] br[250] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_251 bl[251] br[251] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_252 bl[252] br[252] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_253 bl[253] br[253] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_254 bl[254] br[254] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_255 bl[255] br[255] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_256 bl[256] br[256] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_257 bl[257] br[257] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_258 bl[258] br[258] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_259 bl[259] br[259] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_260 bl[260] br[260] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_261 bl[261] br[261] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_262 bl[262] br[262] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_263 bl[263] br[263] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_264 bl[264] br[264] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_265 bl[265] br[265] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_266 bl[266] br[266] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_267 bl[267] br[267] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_268 bl[268] br[268] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_269 bl[269] br[269] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_270 bl[270] br[270] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_271 bl[271] br[271] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_272 bl[272] br[272] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_273 bl[273] br[273] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_274 bl[274] br[274] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_275 bl[275] br[275] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_276 bl[276] br[276] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_277 bl[277] br[277] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_278 bl[278] br[278] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_279 bl[279] br[279] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_280 bl[280] br[280] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_281 bl[281] br[281] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_282 bl[282] br[282] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_283 bl[283] br[283] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_284 bl[284] br[284] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_285 bl[285] br[285] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_286 bl[286] br[286] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_287 bl[287] br[287] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_288 bl[288] br[288] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_289 bl[289] br[289] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_290 bl[290] br[290] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_291 bl[291] br[291] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_292 bl[292] br[292] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_293 bl[293] br[293] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_294 bl[294] br[294] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_295 bl[295] br[295] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_296 bl[296] br[296] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_297 bl[297] br[297] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_298 bl[298] br[298] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_299 bl[299] br[299] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_300 bl[300] br[300] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_301 bl[301] br[301] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_302 bl[302] br[302] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_303 bl[303] br[303] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_304 bl[304] br[304] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_305 bl[305] br[305] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_306 bl[306] br[306] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_307 bl[307] br[307] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_308 bl[308] br[308] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_309 bl[309] br[309] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_310 bl[310] br[310] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_311 bl[311] br[311] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_312 bl[312] br[312] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_313 bl[313] br[313] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_314 bl[314] br[314] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_315 bl[315] br[315] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_316 bl[316] br[316] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_317 bl[317] br[317] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_318 bl[318] br[318] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_319 bl[319] br[319] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_320 bl[320] br[320] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_321 bl[321] br[321] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_322 bl[322] br[322] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_323 bl[323] br[323] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_324 bl[324] br[324] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_325 bl[325] br[325] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_326 bl[326] br[326] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_327 bl[327] br[327] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_328 bl[328] br[328] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_329 bl[329] br[329] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_330 bl[330] br[330] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_331 bl[331] br[331] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_332 bl[332] br[332] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_333 bl[333] br[333] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_334 bl[334] br[334] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_335 bl[335] br[335] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_336 bl[336] br[336] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_337 bl[337] br[337] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_338 bl[338] br[338] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_339 bl[339] br[339] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_340 bl[340] br[340] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_341 bl[341] br[341] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_342 bl[342] br[342] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_343 bl[343] br[343] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_344 bl[344] br[344] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_345 bl[345] br[345] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_346 bl[346] br[346] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_347 bl[347] br[347] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_348 bl[348] br[348] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_349 bl[349] br[349] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_350 bl[350] br[350] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_351 bl[351] br[351] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_352 bl[352] br[352] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_353 bl[353] br[353] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_354 bl[354] br[354] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_355 bl[355] br[355] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_356 bl[356] br[356] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_357 bl[357] br[357] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_358 bl[358] br[358] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_359 bl[359] br[359] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_360 bl[360] br[360] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_361 bl[361] br[361] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_362 bl[362] br[362] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_363 bl[363] br[363] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_364 bl[364] br[364] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_365 bl[365] br[365] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_366 bl[366] br[366] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_367 bl[367] br[367] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_368 bl[368] br[368] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_369 bl[369] br[369] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_370 bl[370] br[370] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_371 bl[371] br[371] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_372 bl[372] br[372] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_373 bl[373] br[373] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_374 bl[374] br[374] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_375 bl[375] br[375] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_376 bl[376] br[376] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_377 bl[377] br[377] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_378 bl[378] br[378] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_379 bl[379] br[379] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_380 bl[380] br[380] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_381 bl[381] br[381] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_382 bl[382] br[382] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_383 bl[383] br[383] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_384 bl[384] br[384] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_385 bl[385] br[385] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_386 bl[386] br[386] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_387 bl[387] br[387] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_388 bl[388] br[388] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_389 bl[389] br[389] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_390 bl[390] br[390] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_391 bl[391] br[391] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_392 bl[392] br[392] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_393 bl[393] br[393] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_394 bl[394] br[394] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_395 bl[395] br[395] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_396 bl[396] br[396] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_397 bl[397] br[397] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_398 bl[398] br[398] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_399 bl[399] br[399] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_400 bl[400] br[400] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_401 bl[401] br[401] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_402 bl[402] br[402] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_403 bl[403] br[403] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_404 bl[404] br[404] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_405 bl[405] br[405] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_406 bl[406] br[406] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_407 bl[407] br[407] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_408 bl[408] br[408] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_409 bl[409] br[409] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_410 bl[410] br[410] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_411 bl[411] br[411] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_412 bl[412] br[412] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_413 bl[413] br[413] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_414 bl[414] br[414] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_415 bl[415] br[415] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_416 bl[416] br[416] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_417 bl[417] br[417] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_418 bl[418] br[418] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_419 bl[419] br[419] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_420 bl[420] br[420] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_421 bl[421] br[421] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_422 bl[422] br[422] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_423 bl[423] br[423] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_424 bl[424] br[424] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_425 bl[425] br[425] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_426 bl[426] br[426] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_427 bl[427] br[427] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_428 bl[428] br[428] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_429 bl[429] br[429] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_430 bl[430] br[430] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_431 bl[431] br[431] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_432 bl[432] br[432] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_433 bl[433] br[433] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_434 bl[434] br[434] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_435 bl[435] br[435] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_436 bl[436] br[436] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_437 bl[437] br[437] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_438 bl[438] br[438] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_439 bl[439] br[439] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_440 bl[440] br[440] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_441 bl[441] br[441] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_442 bl[442] br[442] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_443 bl[443] br[443] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_444 bl[444] br[444] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_445 bl[445] br[445] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_446 bl[446] br[446] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_447 bl[447] br[447] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_448 bl[448] br[448] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_449 bl[449] br[449] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_450 bl[450] br[450] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_451 bl[451] br[451] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_452 bl[452] br[452] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_453 bl[453] br[453] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_454 bl[454] br[454] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_455 bl[455] br[455] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_456 bl[456] br[456] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_457 bl[457] br[457] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_458 bl[458] br[458] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_459 bl[459] br[459] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_460 bl[460] br[460] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_461 bl[461] br[461] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_462 bl[462] br[462] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_463 bl[463] br[463] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_464 bl[464] br[464] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_465 bl[465] br[465] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_466 bl[466] br[466] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_467 bl[467] br[467] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_468 bl[468] br[468] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_469 bl[469] br[469] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_470 bl[470] br[470] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_471 bl[471] br[471] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_472 bl[472] br[472] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_473 bl[473] br[473] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_474 bl[474] br[474] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_475 bl[475] br[475] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_476 bl[476] br[476] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_477 bl[477] br[477] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_478 bl[478] br[478] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_479 bl[479] br[479] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_480 bl[480] br[480] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_481 bl[481] br[481] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_482 bl[482] br[482] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_483 bl[483] br[483] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_484 bl[484] br[484] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_485 bl[485] br[485] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_486 bl[486] br[486] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_487 bl[487] br[487] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_488 bl[488] br[488] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_489 bl[489] br[489] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_490 bl[490] br[490] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_491 bl[491] br[491] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_492 bl[492] br[492] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_493 bl[493] br[493] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_494 bl[494] br[494] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_495 bl[495] br[495] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_496 bl[496] br[496] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_497 bl[497] br[497] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_498 bl[498] br[498] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_499 bl[499] br[499] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_500 bl[500] br[500] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_501 bl[501] br[501] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_502 bl[502] br[502] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_503 bl[503] br[503] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_504 bl[504] br[504] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_505 bl[505] br[505] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_506 bl[506] br[506] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_507 bl[507] br[507] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_508 bl[508] br[508] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_509 bl[509] br[509] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_510 bl[510] br[510] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_20_511 bl[511] br[511] vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xcell_21_0 bl[0] br[0] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_1 bl[1] br[1] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_2 bl[2] br[2] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_3 bl[3] br[3] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_4 bl[4] br[4] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_5 bl[5] br[5] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_6 bl[6] br[6] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_7 bl[7] br[7] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_8 bl[8] br[8] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_9 bl[9] br[9] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_10 bl[10] br[10] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_11 bl[11] br[11] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_12 bl[12] br[12] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_13 bl[13] br[13] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_14 bl[14] br[14] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_15 bl[15] br[15] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_16 bl[16] br[16] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_17 bl[17] br[17] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_18 bl[18] br[18] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_19 bl[19] br[19] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_20 bl[20] br[20] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_21 bl[21] br[21] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_22 bl[22] br[22] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_23 bl[23] br[23] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_24 bl[24] br[24] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_25 bl[25] br[25] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_26 bl[26] br[26] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_27 bl[27] br[27] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_28 bl[28] br[28] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_29 bl[29] br[29] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_30 bl[30] br[30] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_31 bl[31] br[31] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_32 bl[32] br[32] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_33 bl[33] br[33] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_34 bl[34] br[34] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_35 bl[35] br[35] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_36 bl[36] br[36] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_37 bl[37] br[37] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_38 bl[38] br[38] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_39 bl[39] br[39] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_40 bl[40] br[40] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_41 bl[41] br[41] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_42 bl[42] br[42] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_43 bl[43] br[43] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_44 bl[44] br[44] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_45 bl[45] br[45] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_46 bl[46] br[46] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_47 bl[47] br[47] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_48 bl[48] br[48] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_49 bl[49] br[49] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_50 bl[50] br[50] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_51 bl[51] br[51] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_52 bl[52] br[52] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_53 bl[53] br[53] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_54 bl[54] br[54] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_55 bl[55] br[55] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_56 bl[56] br[56] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_57 bl[57] br[57] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_58 bl[58] br[58] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_59 bl[59] br[59] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_60 bl[60] br[60] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_61 bl[61] br[61] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_62 bl[62] br[62] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_63 bl[63] br[63] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_64 bl[64] br[64] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_65 bl[65] br[65] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_66 bl[66] br[66] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_67 bl[67] br[67] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_68 bl[68] br[68] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_69 bl[69] br[69] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_70 bl[70] br[70] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_71 bl[71] br[71] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_72 bl[72] br[72] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_73 bl[73] br[73] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_74 bl[74] br[74] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_75 bl[75] br[75] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_76 bl[76] br[76] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_77 bl[77] br[77] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_78 bl[78] br[78] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_79 bl[79] br[79] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_80 bl[80] br[80] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_81 bl[81] br[81] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_82 bl[82] br[82] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_83 bl[83] br[83] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_84 bl[84] br[84] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_85 bl[85] br[85] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_86 bl[86] br[86] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_87 bl[87] br[87] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_88 bl[88] br[88] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_89 bl[89] br[89] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_90 bl[90] br[90] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_91 bl[91] br[91] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_92 bl[92] br[92] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_93 bl[93] br[93] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_94 bl[94] br[94] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_95 bl[95] br[95] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_96 bl[96] br[96] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_97 bl[97] br[97] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_98 bl[98] br[98] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_99 bl[99] br[99] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_100 bl[100] br[100] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_101 bl[101] br[101] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_102 bl[102] br[102] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_103 bl[103] br[103] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_104 bl[104] br[104] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_105 bl[105] br[105] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_106 bl[106] br[106] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_107 bl[107] br[107] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_108 bl[108] br[108] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_109 bl[109] br[109] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_110 bl[110] br[110] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_111 bl[111] br[111] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_112 bl[112] br[112] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_113 bl[113] br[113] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_114 bl[114] br[114] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_115 bl[115] br[115] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_116 bl[116] br[116] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_117 bl[117] br[117] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_118 bl[118] br[118] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_119 bl[119] br[119] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_120 bl[120] br[120] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_121 bl[121] br[121] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_122 bl[122] br[122] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_123 bl[123] br[123] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_124 bl[124] br[124] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_125 bl[125] br[125] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_126 bl[126] br[126] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_127 bl[127] br[127] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_128 bl[128] br[128] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_129 bl[129] br[129] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_130 bl[130] br[130] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_131 bl[131] br[131] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_132 bl[132] br[132] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_133 bl[133] br[133] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_134 bl[134] br[134] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_135 bl[135] br[135] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_136 bl[136] br[136] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_137 bl[137] br[137] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_138 bl[138] br[138] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_139 bl[139] br[139] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_140 bl[140] br[140] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_141 bl[141] br[141] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_142 bl[142] br[142] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_143 bl[143] br[143] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_144 bl[144] br[144] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_145 bl[145] br[145] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_146 bl[146] br[146] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_147 bl[147] br[147] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_148 bl[148] br[148] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_149 bl[149] br[149] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_150 bl[150] br[150] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_151 bl[151] br[151] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_152 bl[152] br[152] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_153 bl[153] br[153] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_154 bl[154] br[154] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_155 bl[155] br[155] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_156 bl[156] br[156] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_157 bl[157] br[157] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_158 bl[158] br[158] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_159 bl[159] br[159] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_160 bl[160] br[160] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_161 bl[161] br[161] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_162 bl[162] br[162] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_163 bl[163] br[163] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_164 bl[164] br[164] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_165 bl[165] br[165] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_166 bl[166] br[166] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_167 bl[167] br[167] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_168 bl[168] br[168] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_169 bl[169] br[169] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_170 bl[170] br[170] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_171 bl[171] br[171] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_172 bl[172] br[172] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_173 bl[173] br[173] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_174 bl[174] br[174] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_175 bl[175] br[175] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_176 bl[176] br[176] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_177 bl[177] br[177] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_178 bl[178] br[178] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_179 bl[179] br[179] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_180 bl[180] br[180] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_181 bl[181] br[181] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_182 bl[182] br[182] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_183 bl[183] br[183] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_184 bl[184] br[184] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_185 bl[185] br[185] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_186 bl[186] br[186] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_187 bl[187] br[187] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_188 bl[188] br[188] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_189 bl[189] br[189] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_190 bl[190] br[190] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_191 bl[191] br[191] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_192 bl[192] br[192] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_193 bl[193] br[193] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_194 bl[194] br[194] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_195 bl[195] br[195] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_196 bl[196] br[196] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_197 bl[197] br[197] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_198 bl[198] br[198] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_199 bl[199] br[199] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_200 bl[200] br[200] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_201 bl[201] br[201] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_202 bl[202] br[202] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_203 bl[203] br[203] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_204 bl[204] br[204] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_205 bl[205] br[205] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_206 bl[206] br[206] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_207 bl[207] br[207] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_208 bl[208] br[208] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_209 bl[209] br[209] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_210 bl[210] br[210] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_211 bl[211] br[211] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_212 bl[212] br[212] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_213 bl[213] br[213] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_214 bl[214] br[214] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_215 bl[215] br[215] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_216 bl[216] br[216] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_217 bl[217] br[217] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_218 bl[218] br[218] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_219 bl[219] br[219] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_220 bl[220] br[220] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_221 bl[221] br[221] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_222 bl[222] br[222] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_223 bl[223] br[223] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_224 bl[224] br[224] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_225 bl[225] br[225] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_226 bl[226] br[226] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_227 bl[227] br[227] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_228 bl[228] br[228] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_229 bl[229] br[229] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_230 bl[230] br[230] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_231 bl[231] br[231] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_232 bl[232] br[232] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_233 bl[233] br[233] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_234 bl[234] br[234] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_235 bl[235] br[235] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_236 bl[236] br[236] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_237 bl[237] br[237] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_238 bl[238] br[238] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_239 bl[239] br[239] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_240 bl[240] br[240] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_241 bl[241] br[241] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_242 bl[242] br[242] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_243 bl[243] br[243] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_244 bl[244] br[244] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_245 bl[245] br[245] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_246 bl[246] br[246] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_247 bl[247] br[247] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_248 bl[248] br[248] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_249 bl[249] br[249] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_250 bl[250] br[250] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_251 bl[251] br[251] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_252 bl[252] br[252] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_253 bl[253] br[253] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_254 bl[254] br[254] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_255 bl[255] br[255] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_256 bl[256] br[256] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_257 bl[257] br[257] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_258 bl[258] br[258] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_259 bl[259] br[259] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_260 bl[260] br[260] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_261 bl[261] br[261] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_262 bl[262] br[262] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_263 bl[263] br[263] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_264 bl[264] br[264] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_265 bl[265] br[265] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_266 bl[266] br[266] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_267 bl[267] br[267] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_268 bl[268] br[268] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_269 bl[269] br[269] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_270 bl[270] br[270] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_271 bl[271] br[271] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_272 bl[272] br[272] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_273 bl[273] br[273] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_274 bl[274] br[274] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_275 bl[275] br[275] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_276 bl[276] br[276] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_277 bl[277] br[277] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_278 bl[278] br[278] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_279 bl[279] br[279] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_280 bl[280] br[280] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_281 bl[281] br[281] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_282 bl[282] br[282] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_283 bl[283] br[283] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_284 bl[284] br[284] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_285 bl[285] br[285] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_286 bl[286] br[286] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_287 bl[287] br[287] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_288 bl[288] br[288] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_289 bl[289] br[289] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_290 bl[290] br[290] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_291 bl[291] br[291] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_292 bl[292] br[292] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_293 bl[293] br[293] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_294 bl[294] br[294] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_295 bl[295] br[295] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_296 bl[296] br[296] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_297 bl[297] br[297] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_298 bl[298] br[298] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_299 bl[299] br[299] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_300 bl[300] br[300] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_301 bl[301] br[301] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_302 bl[302] br[302] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_303 bl[303] br[303] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_304 bl[304] br[304] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_305 bl[305] br[305] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_306 bl[306] br[306] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_307 bl[307] br[307] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_308 bl[308] br[308] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_309 bl[309] br[309] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_310 bl[310] br[310] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_311 bl[311] br[311] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_312 bl[312] br[312] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_313 bl[313] br[313] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_314 bl[314] br[314] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_315 bl[315] br[315] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_316 bl[316] br[316] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_317 bl[317] br[317] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_318 bl[318] br[318] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_319 bl[319] br[319] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_320 bl[320] br[320] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_321 bl[321] br[321] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_322 bl[322] br[322] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_323 bl[323] br[323] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_324 bl[324] br[324] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_325 bl[325] br[325] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_326 bl[326] br[326] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_327 bl[327] br[327] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_328 bl[328] br[328] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_329 bl[329] br[329] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_330 bl[330] br[330] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_331 bl[331] br[331] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_332 bl[332] br[332] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_333 bl[333] br[333] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_334 bl[334] br[334] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_335 bl[335] br[335] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_336 bl[336] br[336] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_337 bl[337] br[337] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_338 bl[338] br[338] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_339 bl[339] br[339] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_340 bl[340] br[340] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_341 bl[341] br[341] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_342 bl[342] br[342] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_343 bl[343] br[343] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_344 bl[344] br[344] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_345 bl[345] br[345] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_346 bl[346] br[346] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_347 bl[347] br[347] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_348 bl[348] br[348] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_349 bl[349] br[349] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_350 bl[350] br[350] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_351 bl[351] br[351] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_352 bl[352] br[352] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_353 bl[353] br[353] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_354 bl[354] br[354] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_355 bl[355] br[355] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_356 bl[356] br[356] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_357 bl[357] br[357] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_358 bl[358] br[358] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_359 bl[359] br[359] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_360 bl[360] br[360] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_361 bl[361] br[361] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_362 bl[362] br[362] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_363 bl[363] br[363] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_364 bl[364] br[364] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_365 bl[365] br[365] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_366 bl[366] br[366] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_367 bl[367] br[367] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_368 bl[368] br[368] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_369 bl[369] br[369] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_370 bl[370] br[370] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_371 bl[371] br[371] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_372 bl[372] br[372] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_373 bl[373] br[373] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_374 bl[374] br[374] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_375 bl[375] br[375] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_376 bl[376] br[376] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_377 bl[377] br[377] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_378 bl[378] br[378] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_379 bl[379] br[379] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_380 bl[380] br[380] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_381 bl[381] br[381] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_382 bl[382] br[382] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_383 bl[383] br[383] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_384 bl[384] br[384] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_385 bl[385] br[385] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_386 bl[386] br[386] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_387 bl[387] br[387] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_388 bl[388] br[388] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_389 bl[389] br[389] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_390 bl[390] br[390] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_391 bl[391] br[391] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_392 bl[392] br[392] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_393 bl[393] br[393] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_394 bl[394] br[394] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_395 bl[395] br[395] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_396 bl[396] br[396] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_397 bl[397] br[397] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_398 bl[398] br[398] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_399 bl[399] br[399] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_400 bl[400] br[400] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_401 bl[401] br[401] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_402 bl[402] br[402] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_403 bl[403] br[403] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_404 bl[404] br[404] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_405 bl[405] br[405] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_406 bl[406] br[406] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_407 bl[407] br[407] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_408 bl[408] br[408] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_409 bl[409] br[409] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_410 bl[410] br[410] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_411 bl[411] br[411] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_412 bl[412] br[412] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_413 bl[413] br[413] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_414 bl[414] br[414] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_415 bl[415] br[415] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_416 bl[416] br[416] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_417 bl[417] br[417] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_418 bl[418] br[418] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_419 bl[419] br[419] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_420 bl[420] br[420] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_421 bl[421] br[421] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_422 bl[422] br[422] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_423 bl[423] br[423] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_424 bl[424] br[424] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_425 bl[425] br[425] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_426 bl[426] br[426] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_427 bl[427] br[427] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_428 bl[428] br[428] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_429 bl[429] br[429] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_430 bl[430] br[430] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_431 bl[431] br[431] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_432 bl[432] br[432] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_433 bl[433] br[433] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_434 bl[434] br[434] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_435 bl[435] br[435] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_436 bl[436] br[436] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_437 bl[437] br[437] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_438 bl[438] br[438] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_439 bl[439] br[439] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_440 bl[440] br[440] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_441 bl[441] br[441] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_442 bl[442] br[442] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_443 bl[443] br[443] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_444 bl[444] br[444] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_445 bl[445] br[445] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_446 bl[446] br[446] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_447 bl[447] br[447] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_448 bl[448] br[448] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_449 bl[449] br[449] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_450 bl[450] br[450] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_451 bl[451] br[451] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_452 bl[452] br[452] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_453 bl[453] br[453] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_454 bl[454] br[454] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_455 bl[455] br[455] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_456 bl[456] br[456] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_457 bl[457] br[457] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_458 bl[458] br[458] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_459 bl[459] br[459] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_460 bl[460] br[460] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_461 bl[461] br[461] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_462 bl[462] br[462] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_463 bl[463] br[463] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_464 bl[464] br[464] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_465 bl[465] br[465] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_466 bl[466] br[466] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_467 bl[467] br[467] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_468 bl[468] br[468] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_469 bl[469] br[469] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_470 bl[470] br[470] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_471 bl[471] br[471] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_472 bl[472] br[472] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_473 bl[473] br[473] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_474 bl[474] br[474] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_475 bl[475] br[475] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_476 bl[476] br[476] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_477 bl[477] br[477] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_478 bl[478] br[478] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_479 bl[479] br[479] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_480 bl[480] br[480] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_481 bl[481] br[481] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_482 bl[482] br[482] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_483 bl[483] br[483] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_484 bl[484] br[484] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_485 bl[485] br[485] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_486 bl[486] br[486] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_487 bl[487] br[487] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_488 bl[488] br[488] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_489 bl[489] br[489] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_490 bl[490] br[490] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_491 bl[491] br[491] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_492 bl[492] br[492] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_493 bl[493] br[493] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_494 bl[494] br[494] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_495 bl[495] br[495] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_496 bl[496] br[496] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_497 bl[497] br[497] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_498 bl[498] br[498] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_499 bl[499] br[499] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_500 bl[500] br[500] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_501 bl[501] br[501] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_502 bl[502] br[502] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_503 bl[503] br[503] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_504 bl[504] br[504] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_505 bl[505] br[505] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_506 bl[506] br[506] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_507 bl[507] br[507] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_508 bl[508] br[508] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_509 bl[509] br[509] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_510 bl[510] br[510] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_21_511 bl[511] br[511] vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xcell_22_0 bl[0] br[0] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_1 bl[1] br[1] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_2 bl[2] br[2] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_3 bl[3] br[3] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_4 bl[4] br[4] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_5 bl[5] br[5] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_6 bl[6] br[6] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_7 bl[7] br[7] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_8 bl[8] br[8] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_9 bl[9] br[9] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_10 bl[10] br[10] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_11 bl[11] br[11] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_12 bl[12] br[12] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_13 bl[13] br[13] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_14 bl[14] br[14] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_15 bl[15] br[15] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_16 bl[16] br[16] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_17 bl[17] br[17] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_18 bl[18] br[18] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_19 bl[19] br[19] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_20 bl[20] br[20] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_21 bl[21] br[21] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_22 bl[22] br[22] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_23 bl[23] br[23] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_24 bl[24] br[24] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_25 bl[25] br[25] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_26 bl[26] br[26] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_27 bl[27] br[27] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_28 bl[28] br[28] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_29 bl[29] br[29] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_30 bl[30] br[30] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_31 bl[31] br[31] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_32 bl[32] br[32] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_33 bl[33] br[33] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_34 bl[34] br[34] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_35 bl[35] br[35] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_36 bl[36] br[36] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_37 bl[37] br[37] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_38 bl[38] br[38] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_39 bl[39] br[39] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_40 bl[40] br[40] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_41 bl[41] br[41] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_42 bl[42] br[42] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_43 bl[43] br[43] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_44 bl[44] br[44] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_45 bl[45] br[45] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_46 bl[46] br[46] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_47 bl[47] br[47] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_48 bl[48] br[48] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_49 bl[49] br[49] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_50 bl[50] br[50] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_51 bl[51] br[51] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_52 bl[52] br[52] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_53 bl[53] br[53] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_54 bl[54] br[54] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_55 bl[55] br[55] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_56 bl[56] br[56] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_57 bl[57] br[57] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_58 bl[58] br[58] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_59 bl[59] br[59] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_60 bl[60] br[60] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_61 bl[61] br[61] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_62 bl[62] br[62] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_63 bl[63] br[63] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_64 bl[64] br[64] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_65 bl[65] br[65] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_66 bl[66] br[66] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_67 bl[67] br[67] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_68 bl[68] br[68] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_69 bl[69] br[69] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_70 bl[70] br[70] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_71 bl[71] br[71] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_72 bl[72] br[72] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_73 bl[73] br[73] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_74 bl[74] br[74] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_75 bl[75] br[75] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_76 bl[76] br[76] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_77 bl[77] br[77] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_78 bl[78] br[78] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_79 bl[79] br[79] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_80 bl[80] br[80] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_81 bl[81] br[81] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_82 bl[82] br[82] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_83 bl[83] br[83] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_84 bl[84] br[84] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_85 bl[85] br[85] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_86 bl[86] br[86] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_87 bl[87] br[87] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_88 bl[88] br[88] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_89 bl[89] br[89] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_90 bl[90] br[90] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_91 bl[91] br[91] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_92 bl[92] br[92] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_93 bl[93] br[93] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_94 bl[94] br[94] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_95 bl[95] br[95] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_96 bl[96] br[96] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_97 bl[97] br[97] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_98 bl[98] br[98] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_99 bl[99] br[99] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_100 bl[100] br[100] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_101 bl[101] br[101] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_102 bl[102] br[102] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_103 bl[103] br[103] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_104 bl[104] br[104] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_105 bl[105] br[105] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_106 bl[106] br[106] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_107 bl[107] br[107] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_108 bl[108] br[108] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_109 bl[109] br[109] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_110 bl[110] br[110] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_111 bl[111] br[111] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_112 bl[112] br[112] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_113 bl[113] br[113] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_114 bl[114] br[114] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_115 bl[115] br[115] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_116 bl[116] br[116] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_117 bl[117] br[117] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_118 bl[118] br[118] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_119 bl[119] br[119] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_120 bl[120] br[120] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_121 bl[121] br[121] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_122 bl[122] br[122] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_123 bl[123] br[123] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_124 bl[124] br[124] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_125 bl[125] br[125] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_126 bl[126] br[126] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_127 bl[127] br[127] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_128 bl[128] br[128] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_129 bl[129] br[129] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_130 bl[130] br[130] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_131 bl[131] br[131] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_132 bl[132] br[132] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_133 bl[133] br[133] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_134 bl[134] br[134] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_135 bl[135] br[135] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_136 bl[136] br[136] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_137 bl[137] br[137] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_138 bl[138] br[138] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_139 bl[139] br[139] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_140 bl[140] br[140] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_141 bl[141] br[141] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_142 bl[142] br[142] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_143 bl[143] br[143] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_144 bl[144] br[144] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_145 bl[145] br[145] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_146 bl[146] br[146] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_147 bl[147] br[147] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_148 bl[148] br[148] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_149 bl[149] br[149] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_150 bl[150] br[150] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_151 bl[151] br[151] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_152 bl[152] br[152] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_153 bl[153] br[153] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_154 bl[154] br[154] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_155 bl[155] br[155] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_156 bl[156] br[156] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_157 bl[157] br[157] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_158 bl[158] br[158] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_159 bl[159] br[159] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_160 bl[160] br[160] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_161 bl[161] br[161] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_162 bl[162] br[162] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_163 bl[163] br[163] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_164 bl[164] br[164] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_165 bl[165] br[165] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_166 bl[166] br[166] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_167 bl[167] br[167] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_168 bl[168] br[168] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_169 bl[169] br[169] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_170 bl[170] br[170] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_171 bl[171] br[171] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_172 bl[172] br[172] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_173 bl[173] br[173] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_174 bl[174] br[174] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_175 bl[175] br[175] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_176 bl[176] br[176] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_177 bl[177] br[177] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_178 bl[178] br[178] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_179 bl[179] br[179] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_180 bl[180] br[180] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_181 bl[181] br[181] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_182 bl[182] br[182] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_183 bl[183] br[183] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_184 bl[184] br[184] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_185 bl[185] br[185] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_186 bl[186] br[186] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_187 bl[187] br[187] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_188 bl[188] br[188] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_189 bl[189] br[189] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_190 bl[190] br[190] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_191 bl[191] br[191] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_192 bl[192] br[192] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_193 bl[193] br[193] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_194 bl[194] br[194] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_195 bl[195] br[195] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_196 bl[196] br[196] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_197 bl[197] br[197] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_198 bl[198] br[198] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_199 bl[199] br[199] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_200 bl[200] br[200] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_201 bl[201] br[201] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_202 bl[202] br[202] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_203 bl[203] br[203] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_204 bl[204] br[204] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_205 bl[205] br[205] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_206 bl[206] br[206] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_207 bl[207] br[207] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_208 bl[208] br[208] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_209 bl[209] br[209] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_210 bl[210] br[210] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_211 bl[211] br[211] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_212 bl[212] br[212] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_213 bl[213] br[213] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_214 bl[214] br[214] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_215 bl[215] br[215] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_216 bl[216] br[216] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_217 bl[217] br[217] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_218 bl[218] br[218] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_219 bl[219] br[219] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_220 bl[220] br[220] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_221 bl[221] br[221] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_222 bl[222] br[222] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_223 bl[223] br[223] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_224 bl[224] br[224] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_225 bl[225] br[225] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_226 bl[226] br[226] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_227 bl[227] br[227] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_228 bl[228] br[228] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_229 bl[229] br[229] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_230 bl[230] br[230] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_231 bl[231] br[231] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_232 bl[232] br[232] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_233 bl[233] br[233] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_234 bl[234] br[234] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_235 bl[235] br[235] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_236 bl[236] br[236] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_237 bl[237] br[237] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_238 bl[238] br[238] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_239 bl[239] br[239] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_240 bl[240] br[240] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_241 bl[241] br[241] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_242 bl[242] br[242] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_243 bl[243] br[243] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_244 bl[244] br[244] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_245 bl[245] br[245] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_246 bl[246] br[246] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_247 bl[247] br[247] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_248 bl[248] br[248] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_249 bl[249] br[249] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_250 bl[250] br[250] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_251 bl[251] br[251] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_252 bl[252] br[252] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_253 bl[253] br[253] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_254 bl[254] br[254] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_255 bl[255] br[255] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_256 bl[256] br[256] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_257 bl[257] br[257] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_258 bl[258] br[258] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_259 bl[259] br[259] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_260 bl[260] br[260] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_261 bl[261] br[261] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_262 bl[262] br[262] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_263 bl[263] br[263] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_264 bl[264] br[264] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_265 bl[265] br[265] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_266 bl[266] br[266] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_267 bl[267] br[267] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_268 bl[268] br[268] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_269 bl[269] br[269] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_270 bl[270] br[270] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_271 bl[271] br[271] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_272 bl[272] br[272] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_273 bl[273] br[273] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_274 bl[274] br[274] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_275 bl[275] br[275] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_276 bl[276] br[276] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_277 bl[277] br[277] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_278 bl[278] br[278] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_279 bl[279] br[279] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_280 bl[280] br[280] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_281 bl[281] br[281] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_282 bl[282] br[282] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_283 bl[283] br[283] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_284 bl[284] br[284] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_285 bl[285] br[285] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_286 bl[286] br[286] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_287 bl[287] br[287] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_288 bl[288] br[288] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_289 bl[289] br[289] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_290 bl[290] br[290] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_291 bl[291] br[291] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_292 bl[292] br[292] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_293 bl[293] br[293] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_294 bl[294] br[294] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_295 bl[295] br[295] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_296 bl[296] br[296] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_297 bl[297] br[297] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_298 bl[298] br[298] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_299 bl[299] br[299] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_300 bl[300] br[300] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_301 bl[301] br[301] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_302 bl[302] br[302] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_303 bl[303] br[303] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_304 bl[304] br[304] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_305 bl[305] br[305] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_306 bl[306] br[306] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_307 bl[307] br[307] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_308 bl[308] br[308] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_309 bl[309] br[309] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_310 bl[310] br[310] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_311 bl[311] br[311] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_312 bl[312] br[312] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_313 bl[313] br[313] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_314 bl[314] br[314] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_315 bl[315] br[315] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_316 bl[316] br[316] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_317 bl[317] br[317] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_318 bl[318] br[318] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_319 bl[319] br[319] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_320 bl[320] br[320] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_321 bl[321] br[321] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_322 bl[322] br[322] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_323 bl[323] br[323] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_324 bl[324] br[324] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_325 bl[325] br[325] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_326 bl[326] br[326] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_327 bl[327] br[327] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_328 bl[328] br[328] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_329 bl[329] br[329] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_330 bl[330] br[330] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_331 bl[331] br[331] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_332 bl[332] br[332] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_333 bl[333] br[333] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_334 bl[334] br[334] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_335 bl[335] br[335] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_336 bl[336] br[336] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_337 bl[337] br[337] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_338 bl[338] br[338] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_339 bl[339] br[339] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_340 bl[340] br[340] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_341 bl[341] br[341] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_342 bl[342] br[342] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_343 bl[343] br[343] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_344 bl[344] br[344] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_345 bl[345] br[345] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_346 bl[346] br[346] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_347 bl[347] br[347] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_348 bl[348] br[348] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_349 bl[349] br[349] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_350 bl[350] br[350] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_351 bl[351] br[351] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_352 bl[352] br[352] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_353 bl[353] br[353] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_354 bl[354] br[354] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_355 bl[355] br[355] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_356 bl[356] br[356] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_357 bl[357] br[357] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_358 bl[358] br[358] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_359 bl[359] br[359] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_360 bl[360] br[360] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_361 bl[361] br[361] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_362 bl[362] br[362] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_363 bl[363] br[363] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_364 bl[364] br[364] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_365 bl[365] br[365] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_366 bl[366] br[366] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_367 bl[367] br[367] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_368 bl[368] br[368] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_369 bl[369] br[369] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_370 bl[370] br[370] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_371 bl[371] br[371] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_372 bl[372] br[372] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_373 bl[373] br[373] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_374 bl[374] br[374] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_375 bl[375] br[375] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_376 bl[376] br[376] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_377 bl[377] br[377] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_378 bl[378] br[378] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_379 bl[379] br[379] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_380 bl[380] br[380] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_381 bl[381] br[381] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_382 bl[382] br[382] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_383 bl[383] br[383] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_384 bl[384] br[384] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_385 bl[385] br[385] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_386 bl[386] br[386] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_387 bl[387] br[387] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_388 bl[388] br[388] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_389 bl[389] br[389] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_390 bl[390] br[390] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_391 bl[391] br[391] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_392 bl[392] br[392] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_393 bl[393] br[393] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_394 bl[394] br[394] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_395 bl[395] br[395] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_396 bl[396] br[396] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_397 bl[397] br[397] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_398 bl[398] br[398] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_399 bl[399] br[399] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_400 bl[400] br[400] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_401 bl[401] br[401] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_402 bl[402] br[402] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_403 bl[403] br[403] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_404 bl[404] br[404] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_405 bl[405] br[405] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_406 bl[406] br[406] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_407 bl[407] br[407] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_408 bl[408] br[408] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_409 bl[409] br[409] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_410 bl[410] br[410] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_411 bl[411] br[411] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_412 bl[412] br[412] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_413 bl[413] br[413] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_414 bl[414] br[414] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_415 bl[415] br[415] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_416 bl[416] br[416] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_417 bl[417] br[417] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_418 bl[418] br[418] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_419 bl[419] br[419] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_420 bl[420] br[420] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_421 bl[421] br[421] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_422 bl[422] br[422] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_423 bl[423] br[423] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_424 bl[424] br[424] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_425 bl[425] br[425] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_426 bl[426] br[426] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_427 bl[427] br[427] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_428 bl[428] br[428] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_429 bl[429] br[429] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_430 bl[430] br[430] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_431 bl[431] br[431] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_432 bl[432] br[432] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_433 bl[433] br[433] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_434 bl[434] br[434] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_435 bl[435] br[435] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_436 bl[436] br[436] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_437 bl[437] br[437] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_438 bl[438] br[438] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_439 bl[439] br[439] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_440 bl[440] br[440] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_441 bl[441] br[441] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_442 bl[442] br[442] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_443 bl[443] br[443] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_444 bl[444] br[444] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_445 bl[445] br[445] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_446 bl[446] br[446] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_447 bl[447] br[447] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_448 bl[448] br[448] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_449 bl[449] br[449] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_450 bl[450] br[450] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_451 bl[451] br[451] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_452 bl[452] br[452] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_453 bl[453] br[453] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_454 bl[454] br[454] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_455 bl[455] br[455] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_456 bl[456] br[456] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_457 bl[457] br[457] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_458 bl[458] br[458] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_459 bl[459] br[459] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_460 bl[460] br[460] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_461 bl[461] br[461] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_462 bl[462] br[462] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_463 bl[463] br[463] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_464 bl[464] br[464] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_465 bl[465] br[465] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_466 bl[466] br[466] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_467 bl[467] br[467] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_468 bl[468] br[468] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_469 bl[469] br[469] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_470 bl[470] br[470] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_471 bl[471] br[471] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_472 bl[472] br[472] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_473 bl[473] br[473] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_474 bl[474] br[474] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_475 bl[475] br[475] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_476 bl[476] br[476] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_477 bl[477] br[477] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_478 bl[478] br[478] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_479 bl[479] br[479] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_480 bl[480] br[480] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_481 bl[481] br[481] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_482 bl[482] br[482] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_483 bl[483] br[483] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_484 bl[484] br[484] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_485 bl[485] br[485] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_486 bl[486] br[486] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_487 bl[487] br[487] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_488 bl[488] br[488] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_489 bl[489] br[489] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_490 bl[490] br[490] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_491 bl[491] br[491] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_492 bl[492] br[492] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_493 bl[493] br[493] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_494 bl[494] br[494] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_495 bl[495] br[495] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_496 bl[496] br[496] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_497 bl[497] br[497] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_498 bl[498] br[498] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_499 bl[499] br[499] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_500 bl[500] br[500] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_501 bl[501] br[501] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_502 bl[502] br[502] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_503 bl[503] br[503] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_504 bl[504] br[504] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_505 bl[505] br[505] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_506 bl[506] br[506] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_507 bl[507] br[507] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_508 bl[508] br[508] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_509 bl[509] br[509] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_510 bl[510] br[510] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_22_511 bl[511] br[511] vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xcell_23_0 bl[0] br[0] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_1 bl[1] br[1] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_2 bl[2] br[2] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_3 bl[3] br[3] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_4 bl[4] br[4] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_5 bl[5] br[5] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_6 bl[6] br[6] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_7 bl[7] br[7] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_8 bl[8] br[8] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_9 bl[9] br[9] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_10 bl[10] br[10] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_11 bl[11] br[11] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_12 bl[12] br[12] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_13 bl[13] br[13] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_14 bl[14] br[14] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_15 bl[15] br[15] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_16 bl[16] br[16] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_17 bl[17] br[17] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_18 bl[18] br[18] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_19 bl[19] br[19] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_20 bl[20] br[20] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_21 bl[21] br[21] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_22 bl[22] br[22] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_23 bl[23] br[23] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_24 bl[24] br[24] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_25 bl[25] br[25] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_26 bl[26] br[26] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_27 bl[27] br[27] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_28 bl[28] br[28] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_29 bl[29] br[29] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_30 bl[30] br[30] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_31 bl[31] br[31] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_32 bl[32] br[32] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_33 bl[33] br[33] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_34 bl[34] br[34] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_35 bl[35] br[35] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_36 bl[36] br[36] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_37 bl[37] br[37] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_38 bl[38] br[38] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_39 bl[39] br[39] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_40 bl[40] br[40] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_41 bl[41] br[41] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_42 bl[42] br[42] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_43 bl[43] br[43] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_44 bl[44] br[44] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_45 bl[45] br[45] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_46 bl[46] br[46] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_47 bl[47] br[47] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_48 bl[48] br[48] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_49 bl[49] br[49] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_50 bl[50] br[50] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_51 bl[51] br[51] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_52 bl[52] br[52] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_53 bl[53] br[53] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_54 bl[54] br[54] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_55 bl[55] br[55] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_56 bl[56] br[56] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_57 bl[57] br[57] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_58 bl[58] br[58] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_59 bl[59] br[59] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_60 bl[60] br[60] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_61 bl[61] br[61] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_62 bl[62] br[62] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_63 bl[63] br[63] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_64 bl[64] br[64] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_65 bl[65] br[65] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_66 bl[66] br[66] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_67 bl[67] br[67] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_68 bl[68] br[68] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_69 bl[69] br[69] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_70 bl[70] br[70] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_71 bl[71] br[71] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_72 bl[72] br[72] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_73 bl[73] br[73] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_74 bl[74] br[74] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_75 bl[75] br[75] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_76 bl[76] br[76] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_77 bl[77] br[77] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_78 bl[78] br[78] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_79 bl[79] br[79] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_80 bl[80] br[80] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_81 bl[81] br[81] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_82 bl[82] br[82] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_83 bl[83] br[83] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_84 bl[84] br[84] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_85 bl[85] br[85] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_86 bl[86] br[86] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_87 bl[87] br[87] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_88 bl[88] br[88] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_89 bl[89] br[89] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_90 bl[90] br[90] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_91 bl[91] br[91] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_92 bl[92] br[92] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_93 bl[93] br[93] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_94 bl[94] br[94] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_95 bl[95] br[95] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_96 bl[96] br[96] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_97 bl[97] br[97] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_98 bl[98] br[98] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_99 bl[99] br[99] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_100 bl[100] br[100] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_101 bl[101] br[101] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_102 bl[102] br[102] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_103 bl[103] br[103] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_104 bl[104] br[104] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_105 bl[105] br[105] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_106 bl[106] br[106] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_107 bl[107] br[107] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_108 bl[108] br[108] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_109 bl[109] br[109] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_110 bl[110] br[110] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_111 bl[111] br[111] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_112 bl[112] br[112] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_113 bl[113] br[113] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_114 bl[114] br[114] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_115 bl[115] br[115] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_116 bl[116] br[116] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_117 bl[117] br[117] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_118 bl[118] br[118] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_119 bl[119] br[119] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_120 bl[120] br[120] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_121 bl[121] br[121] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_122 bl[122] br[122] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_123 bl[123] br[123] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_124 bl[124] br[124] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_125 bl[125] br[125] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_126 bl[126] br[126] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_127 bl[127] br[127] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_128 bl[128] br[128] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_129 bl[129] br[129] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_130 bl[130] br[130] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_131 bl[131] br[131] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_132 bl[132] br[132] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_133 bl[133] br[133] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_134 bl[134] br[134] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_135 bl[135] br[135] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_136 bl[136] br[136] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_137 bl[137] br[137] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_138 bl[138] br[138] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_139 bl[139] br[139] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_140 bl[140] br[140] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_141 bl[141] br[141] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_142 bl[142] br[142] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_143 bl[143] br[143] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_144 bl[144] br[144] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_145 bl[145] br[145] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_146 bl[146] br[146] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_147 bl[147] br[147] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_148 bl[148] br[148] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_149 bl[149] br[149] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_150 bl[150] br[150] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_151 bl[151] br[151] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_152 bl[152] br[152] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_153 bl[153] br[153] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_154 bl[154] br[154] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_155 bl[155] br[155] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_156 bl[156] br[156] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_157 bl[157] br[157] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_158 bl[158] br[158] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_159 bl[159] br[159] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_160 bl[160] br[160] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_161 bl[161] br[161] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_162 bl[162] br[162] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_163 bl[163] br[163] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_164 bl[164] br[164] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_165 bl[165] br[165] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_166 bl[166] br[166] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_167 bl[167] br[167] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_168 bl[168] br[168] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_169 bl[169] br[169] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_170 bl[170] br[170] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_171 bl[171] br[171] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_172 bl[172] br[172] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_173 bl[173] br[173] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_174 bl[174] br[174] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_175 bl[175] br[175] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_176 bl[176] br[176] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_177 bl[177] br[177] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_178 bl[178] br[178] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_179 bl[179] br[179] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_180 bl[180] br[180] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_181 bl[181] br[181] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_182 bl[182] br[182] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_183 bl[183] br[183] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_184 bl[184] br[184] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_185 bl[185] br[185] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_186 bl[186] br[186] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_187 bl[187] br[187] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_188 bl[188] br[188] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_189 bl[189] br[189] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_190 bl[190] br[190] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_191 bl[191] br[191] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_192 bl[192] br[192] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_193 bl[193] br[193] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_194 bl[194] br[194] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_195 bl[195] br[195] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_196 bl[196] br[196] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_197 bl[197] br[197] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_198 bl[198] br[198] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_199 bl[199] br[199] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_200 bl[200] br[200] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_201 bl[201] br[201] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_202 bl[202] br[202] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_203 bl[203] br[203] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_204 bl[204] br[204] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_205 bl[205] br[205] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_206 bl[206] br[206] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_207 bl[207] br[207] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_208 bl[208] br[208] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_209 bl[209] br[209] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_210 bl[210] br[210] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_211 bl[211] br[211] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_212 bl[212] br[212] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_213 bl[213] br[213] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_214 bl[214] br[214] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_215 bl[215] br[215] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_216 bl[216] br[216] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_217 bl[217] br[217] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_218 bl[218] br[218] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_219 bl[219] br[219] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_220 bl[220] br[220] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_221 bl[221] br[221] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_222 bl[222] br[222] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_223 bl[223] br[223] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_224 bl[224] br[224] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_225 bl[225] br[225] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_226 bl[226] br[226] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_227 bl[227] br[227] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_228 bl[228] br[228] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_229 bl[229] br[229] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_230 bl[230] br[230] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_231 bl[231] br[231] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_232 bl[232] br[232] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_233 bl[233] br[233] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_234 bl[234] br[234] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_235 bl[235] br[235] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_236 bl[236] br[236] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_237 bl[237] br[237] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_238 bl[238] br[238] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_239 bl[239] br[239] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_240 bl[240] br[240] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_241 bl[241] br[241] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_242 bl[242] br[242] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_243 bl[243] br[243] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_244 bl[244] br[244] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_245 bl[245] br[245] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_246 bl[246] br[246] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_247 bl[247] br[247] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_248 bl[248] br[248] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_249 bl[249] br[249] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_250 bl[250] br[250] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_251 bl[251] br[251] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_252 bl[252] br[252] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_253 bl[253] br[253] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_254 bl[254] br[254] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_255 bl[255] br[255] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_256 bl[256] br[256] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_257 bl[257] br[257] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_258 bl[258] br[258] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_259 bl[259] br[259] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_260 bl[260] br[260] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_261 bl[261] br[261] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_262 bl[262] br[262] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_263 bl[263] br[263] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_264 bl[264] br[264] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_265 bl[265] br[265] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_266 bl[266] br[266] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_267 bl[267] br[267] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_268 bl[268] br[268] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_269 bl[269] br[269] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_270 bl[270] br[270] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_271 bl[271] br[271] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_272 bl[272] br[272] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_273 bl[273] br[273] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_274 bl[274] br[274] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_275 bl[275] br[275] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_276 bl[276] br[276] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_277 bl[277] br[277] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_278 bl[278] br[278] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_279 bl[279] br[279] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_280 bl[280] br[280] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_281 bl[281] br[281] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_282 bl[282] br[282] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_283 bl[283] br[283] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_284 bl[284] br[284] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_285 bl[285] br[285] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_286 bl[286] br[286] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_287 bl[287] br[287] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_288 bl[288] br[288] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_289 bl[289] br[289] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_290 bl[290] br[290] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_291 bl[291] br[291] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_292 bl[292] br[292] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_293 bl[293] br[293] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_294 bl[294] br[294] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_295 bl[295] br[295] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_296 bl[296] br[296] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_297 bl[297] br[297] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_298 bl[298] br[298] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_299 bl[299] br[299] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_300 bl[300] br[300] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_301 bl[301] br[301] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_302 bl[302] br[302] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_303 bl[303] br[303] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_304 bl[304] br[304] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_305 bl[305] br[305] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_306 bl[306] br[306] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_307 bl[307] br[307] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_308 bl[308] br[308] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_309 bl[309] br[309] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_310 bl[310] br[310] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_311 bl[311] br[311] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_312 bl[312] br[312] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_313 bl[313] br[313] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_314 bl[314] br[314] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_315 bl[315] br[315] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_316 bl[316] br[316] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_317 bl[317] br[317] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_318 bl[318] br[318] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_319 bl[319] br[319] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_320 bl[320] br[320] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_321 bl[321] br[321] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_322 bl[322] br[322] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_323 bl[323] br[323] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_324 bl[324] br[324] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_325 bl[325] br[325] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_326 bl[326] br[326] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_327 bl[327] br[327] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_328 bl[328] br[328] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_329 bl[329] br[329] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_330 bl[330] br[330] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_331 bl[331] br[331] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_332 bl[332] br[332] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_333 bl[333] br[333] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_334 bl[334] br[334] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_335 bl[335] br[335] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_336 bl[336] br[336] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_337 bl[337] br[337] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_338 bl[338] br[338] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_339 bl[339] br[339] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_340 bl[340] br[340] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_341 bl[341] br[341] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_342 bl[342] br[342] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_343 bl[343] br[343] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_344 bl[344] br[344] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_345 bl[345] br[345] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_346 bl[346] br[346] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_347 bl[347] br[347] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_348 bl[348] br[348] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_349 bl[349] br[349] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_350 bl[350] br[350] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_351 bl[351] br[351] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_352 bl[352] br[352] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_353 bl[353] br[353] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_354 bl[354] br[354] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_355 bl[355] br[355] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_356 bl[356] br[356] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_357 bl[357] br[357] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_358 bl[358] br[358] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_359 bl[359] br[359] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_360 bl[360] br[360] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_361 bl[361] br[361] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_362 bl[362] br[362] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_363 bl[363] br[363] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_364 bl[364] br[364] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_365 bl[365] br[365] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_366 bl[366] br[366] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_367 bl[367] br[367] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_368 bl[368] br[368] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_369 bl[369] br[369] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_370 bl[370] br[370] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_371 bl[371] br[371] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_372 bl[372] br[372] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_373 bl[373] br[373] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_374 bl[374] br[374] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_375 bl[375] br[375] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_376 bl[376] br[376] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_377 bl[377] br[377] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_378 bl[378] br[378] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_379 bl[379] br[379] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_380 bl[380] br[380] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_381 bl[381] br[381] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_382 bl[382] br[382] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_383 bl[383] br[383] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_384 bl[384] br[384] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_385 bl[385] br[385] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_386 bl[386] br[386] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_387 bl[387] br[387] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_388 bl[388] br[388] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_389 bl[389] br[389] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_390 bl[390] br[390] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_391 bl[391] br[391] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_392 bl[392] br[392] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_393 bl[393] br[393] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_394 bl[394] br[394] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_395 bl[395] br[395] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_396 bl[396] br[396] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_397 bl[397] br[397] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_398 bl[398] br[398] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_399 bl[399] br[399] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_400 bl[400] br[400] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_401 bl[401] br[401] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_402 bl[402] br[402] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_403 bl[403] br[403] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_404 bl[404] br[404] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_405 bl[405] br[405] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_406 bl[406] br[406] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_407 bl[407] br[407] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_408 bl[408] br[408] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_409 bl[409] br[409] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_410 bl[410] br[410] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_411 bl[411] br[411] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_412 bl[412] br[412] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_413 bl[413] br[413] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_414 bl[414] br[414] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_415 bl[415] br[415] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_416 bl[416] br[416] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_417 bl[417] br[417] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_418 bl[418] br[418] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_419 bl[419] br[419] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_420 bl[420] br[420] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_421 bl[421] br[421] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_422 bl[422] br[422] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_423 bl[423] br[423] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_424 bl[424] br[424] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_425 bl[425] br[425] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_426 bl[426] br[426] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_427 bl[427] br[427] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_428 bl[428] br[428] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_429 bl[429] br[429] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_430 bl[430] br[430] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_431 bl[431] br[431] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_432 bl[432] br[432] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_433 bl[433] br[433] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_434 bl[434] br[434] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_435 bl[435] br[435] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_436 bl[436] br[436] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_437 bl[437] br[437] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_438 bl[438] br[438] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_439 bl[439] br[439] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_440 bl[440] br[440] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_441 bl[441] br[441] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_442 bl[442] br[442] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_443 bl[443] br[443] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_444 bl[444] br[444] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_445 bl[445] br[445] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_446 bl[446] br[446] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_447 bl[447] br[447] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_448 bl[448] br[448] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_449 bl[449] br[449] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_450 bl[450] br[450] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_451 bl[451] br[451] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_452 bl[452] br[452] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_453 bl[453] br[453] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_454 bl[454] br[454] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_455 bl[455] br[455] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_456 bl[456] br[456] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_457 bl[457] br[457] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_458 bl[458] br[458] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_459 bl[459] br[459] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_460 bl[460] br[460] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_461 bl[461] br[461] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_462 bl[462] br[462] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_463 bl[463] br[463] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_464 bl[464] br[464] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_465 bl[465] br[465] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_466 bl[466] br[466] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_467 bl[467] br[467] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_468 bl[468] br[468] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_469 bl[469] br[469] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_470 bl[470] br[470] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_471 bl[471] br[471] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_472 bl[472] br[472] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_473 bl[473] br[473] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_474 bl[474] br[474] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_475 bl[475] br[475] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_476 bl[476] br[476] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_477 bl[477] br[477] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_478 bl[478] br[478] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_479 bl[479] br[479] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_480 bl[480] br[480] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_481 bl[481] br[481] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_482 bl[482] br[482] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_483 bl[483] br[483] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_484 bl[484] br[484] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_485 bl[485] br[485] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_486 bl[486] br[486] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_487 bl[487] br[487] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_488 bl[488] br[488] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_489 bl[489] br[489] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_490 bl[490] br[490] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_491 bl[491] br[491] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_492 bl[492] br[492] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_493 bl[493] br[493] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_494 bl[494] br[494] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_495 bl[495] br[495] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_496 bl[496] br[496] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_497 bl[497] br[497] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_498 bl[498] br[498] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_499 bl[499] br[499] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_500 bl[500] br[500] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_501 bl[501] br[501] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_502 bl[502] br[502] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_503 bl[503] br[503] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_504 bl[504] br[504] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_505 bl[505] br[505] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_506 bl[506] br[506] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_507 bl[507] br[507] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_508 bl[508] br[508] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_509 bl[509] br[509] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_510 bl[510] br[510] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_23_511 bl[511] br[511] vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xcell_24_0 bl[0] br[0] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_1 bl[1] br[1] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_2 bl[2] br[2] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_3 bl[3] br[3] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_4 bl[4] br[4] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_5 bl[5] br[5] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_6 bl[6] br[6] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_7 bl[7] br[7] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_8 bl[8] br[8] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_9 bl[9] br[9] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_10 bl[10] br[10] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_11 bl[11] br[11] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_12 bl[12] br[12] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_13 bl[13] br[13] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_14 bl[14] br[14] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_15 bl[15] br[15] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_16 bl[16] br[16] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_17 bl[17] br[17] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_18 bl[18] br[18] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_19 bl[19] br[19] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_20 bl[20] br[20] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_21 bl[21] br[21] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_22 bl[22] br[22] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_23 bl[23] br[23] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_24 bl[24] br[24] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_25 bl[25] br[25] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_26 bl[26] br[26] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_27 bl[27] br[27] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_28 bl[28] br[28] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_29 bl[29] br[29] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_30 bl[30] br[30] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_31 bl[31] br[31] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_32 bl[32] br[32] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_33 bl[33] br[33] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_34 bl[34] br[34] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_35 bl[35] br[35] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_36 bl[36] br[36] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_37 bl[37] br[37] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_38 bl[38] br[38] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_39 bl[39] br[39] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_40 bl[40] br[40] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_41 bl[41] br[41] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_42 bl[42] br[42] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_43 bl[43] br[43] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_44 bl[44] br[44] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_45 bl[45] br[45] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_46 bl[46] br[46] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_47 bl[47] br[47] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_48 bl[48] br[48] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_49 bl[49] br[49] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_50 bl[50] br[50] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_51 bl[51] br[51] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_52 bl[52] br[52] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_53 bl[53] br[53] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_54 bl[54] br[54] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_55 bl[55] br[55] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_56 bl[56] br[56] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_57 bl[57] br[57] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_58 bl[58] br[58] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_59 bl[59] br[59] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_60 bl[60] br[60] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_61 bl[61] br[61] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_62 bl[62] br[62] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_63 bl[63] br[63] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_64 bl[64] br[64] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_65 bl[65] br[65] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_66 bl[66] br[66] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_67 bl[67] br[67] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_68 bl[68] br[68] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_69 bl[69] br[69] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_70 bl[70] br[70] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_71 bl[71] br[71] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_72 bl[72] br[72] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_73 bl[73] br[73] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_74 bl[74] br[74] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_75 bl[75] br[75] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_76 bl[76] br[76] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_77 bl[77] br[77] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_78 bl[78] br[78] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_79 bl[79] br[79] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_80 bl[80] br[80] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_81 bl[81] br[81] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_82 bl[82] br[82] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_83 bl[83] br[83] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_84 bl[84] br[84] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_85 bl[85] br[85] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_86 bl[86] br[86] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_87 bl[87] br[87] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_88 bl[88] br[88] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_89 bl[89] br[89] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_90 bl[90] br[90] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_91 bl[91] br[91] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_92 bl[92] br[92] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_93 bl[93] br[93] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_94 bl[94] br[94] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_95 bl[95] br[95] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_96 bl[96] br[96] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_97 bl[97] br[97] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_98 bl[98] br[98] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_99 bl[99] br[99] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_100 bl[100] br[100] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_101 bl[101] br[101] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_102 bl[102] br[102] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_103 bl[103] br[103] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_104 bl[104] br[104] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_105 bl[105] br[105] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_106 bl[106] br[106] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_107 bl[107] br[107] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_108 bl[108] br[108] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_109 bl[109] br[109] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_110 bl[110] br[110] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_111 bl[111] br[111] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_112 bl[112] br[112] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_113 bl[113] br[113] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_114 bl[114] br[114] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_115 bl[115] br[115] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_116 bl[116] br[116] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_117 bl[117] br[117] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_118 bl[118] br[118] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_119 bl[119] br[119] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_120 bl[120] br[120] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_121 bl[121] br[121] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_122 bl[122] br[122] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_123 bl[123] br[123] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_124 bl[124] br[124] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_125 bl[125] br[125] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_126 bl[126] br[126] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_127 bl[127] br[127] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_128 bl[128] br[128] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_129 bl[129] br[129] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_130 bl[130] br[130] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_131 bl[131] br[131] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_132 bl[132] br[132] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_133 bl[133] br[133] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_134 bl[134] br[134] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_135 bl[135] br[135] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_136 bl[136] br[136] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_137 bl[137] br[137] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_138 bl[138] br[138] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_139 bl[139] br[139] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_140 bl[140] br[140] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_141 bl[141] br[141] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_142 bl[142] br[142] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_143 bl[143] br[143] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_144 bl[144] br[144] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_145 bl[145] br[145] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_146 bl[146] br[146] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_147 bl[147] br[147] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_148 bl[148] br[148] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_149 bl[149] br[149] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_150 bl[150] br[150] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_151 bl[151] br[151] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_152 bl[152] br[152] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_153 bl[153] br[153] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_154 bl[154] br[154] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_155 bl[155] br[155] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_156 bl[156] br[156] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_157 bl[157] br[157] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_158 bl[158] br[158] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_159 bl[159] br[159] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_160 bl[160] br[160] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_161 bl[161] br[161] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_162 bl[162] br[162] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_163 bl[163] br[163] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_164 bl[164] br[164] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_165 bl[165] br[165] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_166 bl[166] br[166] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_167 bl[167] br[167] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_168 bl[168] br[168] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_169 bl[169] br[169] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_170 bl[170] br[170] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_171 bl[171] br[171] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_172 bl[172] br[172] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_173 bl[173] br[173] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_174 bl[174] br[174] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_175 bl[175] br[175] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_176 bl[176] br[176] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_177 bl[177] br[177] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_178 bl[178] br[178] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_179 bl[179] br[179] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_180 bl[180] br[180] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_181 bl[181] br[181] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_182 bl[182] br[182] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_183 bl[183] br[183] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_184 bl[184] br[184] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_185 bl[185] br[185] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_186 bl[186] br[186] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_187 bl[187] br[187] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_188 bl[188] br[188] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_189 bl[189] br[189] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_190 bl[190] br[190] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_191 bl[191] br[191] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_192 bl[192] br[192] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_193 bl[193] br[193] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_194 bl[194] br[194] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_195 bl[195] br[195] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_196 bl[196] br[196] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_197 bl[197] br[197] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_198 bl[198] br[198] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_199 bl[199] br[199] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_200 bl[200] br[200] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_201 bl[201] br[201] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_202 bl[202] br[202] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_203 bl[203] br[203] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_204 bl[204] br[204] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_205 bl[205] br[205] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_206 bl[206] br[206] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_207 bl[207] br[207] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_208 bl[208] br[208] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_209 bl[209] br[209] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_210 bl[210] br[210] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_211 bl[211] br[211] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_212 bl[212] br[212] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_213 bl[213] br[213] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_214 bl[214] br[214] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_215 bl[215] br[215] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_216 bl[216] br[216] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_217 bl[217] br[217] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_218 bl[218] br[218] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_219 bl[219] br[219] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_220 bl[220] br[220] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_221 bl[221] br[221] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_222 bl[222] br[222] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_223 bl[223] br[223] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_224 bl[224] br[224] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_225 bl[225] br[225] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_226 bl[226] br[226] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_227 bl[227] br[227] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_228 bl[228] br[228] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_229 bl[229] br[229] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_230 bl[230] br[230] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_231 bl[231] br[231] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_232 bl[232] br[232] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_233 bl[233] br[233] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_234 bl[234] br[234] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_235 bl[235] br[235] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_236 bl[236] br[236] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_237 bl[237] br[237] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_238 bl[238] br[238] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_239 bl[239] br[239] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_240 bl[240] br[240] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_241 bl[241] br[241] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_242 bl[242] br[242] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_243 bl[243] br[243] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_244 bl[244] br[244] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_245 bl[245] br[245] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_246 bl[246] br[246] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_247 bl[247] br[247] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_248 bl[248] br[248] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_249 bl[249] br[249] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_250 bl[250] br[250] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_251 bl[251] br[251] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_252 bl[252] br[252] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_253 bl[253] br[253] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_254 bl[254] br[254] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_255 bl[255] br[255] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_256 bl[256] br[256] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_257 bl[257] br[257] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_258 bl[258] br[258] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_259 bl[259] br[259] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_260 bl[260] br[260] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_261 bl[261] br[261] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_262 bl[262] br[262] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_263 bl[263] br[263] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_264 bl[264] br[264] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_265 bl[265] br[265] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_266 bl[266] br[266] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_267 bl[267] br[267] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_268 bl[268] br[268] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_269 bl[269] br[269] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_270 bl[270] br[270] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_271 bl[271] br[271] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_272 bl[272] br[272] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_273 bl[273] br[273] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_274 bl[274] br[274] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_275 bl[275] br[275] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_276 bl[276] br[276] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_277 bl[277] br[277] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_278 bl[278] br[278] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_279 bl[279] br[279] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_280 bl[280] br[280] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_281 bl[281] br[281] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_282 bl[282] br[282] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_283 bl[283] br[283] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_284 bl[284] br[284] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_285 bl[285] br[285] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_286 bl[286] br[286] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_287 bl[287] br[287] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_288 bl[288] br[288] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_289 bl[289] br[289] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_290 bl[290] br[290] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_291 bl[291] br[291] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_292 bl[292] br[292] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_293 bl[293] br[293] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_294 bl[294] br[294] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_295 bl[295] br[295] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_296 bl[296] br[296] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_297 bl[297] br[297] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_298 bl[298] br[298] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_299 bl[299] br[299] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_300 bl[300] br[300] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_301 bl[301] br[301] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_302 bl[302] br[302] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_303 bl[303] br[303] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_304 bl[304] br[304] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_305 bl[305] br[305] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_306 bl[306] br[306] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_307 bl[307] br[307] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_308 bl[308] br[308] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_309 bl[309] br[309] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_310 bl[310] br[310] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_311 bl[311] br[311] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_312 bl[312] br[312] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_313 bl[313] br[313] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_314 bl[314] br[314] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_315 bl[315] br[315] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_316 bl[316] br[316] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_317 bl[317] br[317] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_318 bl[318] br[318] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_319 bl[319] br[319] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_320 bl[320] br[320] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_321 bl[321] br[321] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_322 bl[322] br[322] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_323 bl[323] br[323] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_324 bl[324] br[324] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_325 bl[325] br[325] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_326 bl[326] br[326] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_327 bl[327] br[327] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_328 bl[328] br[328] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_329 bl[329] br[329] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_330 bl[330] br[330] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_331 bl[331] br[331] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_332 bl[332] br[332] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_333 bl[333] br[333] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_334 bl[334] br[334] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_335 bl[335] br[335] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_336 bl[336] br[336] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_337 bl[337] br[337] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_338 bl[338] br[338] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_339 bl[339] br[339] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_340 bl[340] br[340] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_341 bl[341] br[341] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_342 bl[342] br[342] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_343 bl[343] br[343] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_344 bl[344] br[344] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_345 bl[345] br[345] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_346 bl[346] br[346] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_347 bl[347] br[347] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_348 bl[348] br[348] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_349 bl[349] br[349] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_350 bl[350] br[350] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_351 bl[351] br[351] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_352 bl[352] br[352] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_353 bl[353] br[353] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_354 bl[354] br[354] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_355 bl[355] br[355] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_356 bl[356] br[356] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_357 bl[357] br[357] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_358 bl[358] br[358] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_359 bl[359] br[359] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_360 bl[360] br[360] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_361 bl[361] br[361] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_362 bl[362] br[362] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_363 bl[363] br[363] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_364 bl[364] br[364] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_365 bl[365] br[365] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_366 bl[366] br[366] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_367 bl[367] br[367] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_368 bl[368] br[368] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_369 bl[369] br[369] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_370 bl[370] br[370] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_371 bl[371] br[371] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_372 bl[372] br[372] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_373 bl[373] br[373] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_374 bl[374] br[374] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_375 bl[375] br[375] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_376 bl[376] br[376] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_377 bl[377] br[377] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_378 bl[378] br[378] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_379 bl[379] br[379] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_380 bl[380] br[380] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_381 bl[381] br[381] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_382 bl[382] br[382] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_383 bl[383] br[383] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_384 bl[384] br[384] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_385 bl[385] br[385] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_386 bl[386] br[386] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_387 bl[387] br[387] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_388 bl[388] br[388] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_389 bl[389] br[389] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_390 bl[390] br[390] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_391 bl[391] br[391] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_392 bl[392] br[392] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_393 bl[393] br[393] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_394 bl[394] br[394] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_395 bl[395] br[395] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_396 bl[396] br[396] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_397 bl[397] br[397] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_398 bl[398] br[398] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_399 bl[399] br[399] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_400 bl[400] br[400] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_401 bl[401] br[401] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_402 bl[402] br[402] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_403 bl[403] br[403] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_404 bl[404] br[404] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_405 bl[405] br[405] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_406 bl[406] br[406] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_407 bl[407] br[407] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_408 bl[408] br[408] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_409 bl[409] br[409] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_410 bl[410] br[410] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_411 bl[411] br[411] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_412 bl[412] br[412] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_413 bl[413] br[413] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_414 bl[414] br[414] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_415 bl[415] br[415] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_416 bl[416] br[416] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_417 bl[417] br[417] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_418 bl[418] br[418] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_419 bl[419] br[419] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_420 bl[420] br[420] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_421 bl[421] br[421] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_422 bl[422] br[422] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_423 bl[423] br[423] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_424 bl[424] br[424] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_425 bl[425] br[425] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_426 bl[426] br[426] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_427 bl[427] br[427] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_428 bl[428] br[428] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_429 bl[429] br[429] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_430 bl[430] br[430] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_431 bl[431] br[431] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_432 bl[432] br[432] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_433 bl[433] br[433] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_434 bl[434] br[434] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_435 bl[435] br[435] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_436 bl[436] br[436] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_437 bl[437] br[437] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_438 bl[438] br[438] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_439 bl[439] br[439] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_440 bl[440] br[440] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_441 bl[441] br[441] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_442 bl[442] br[442] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_443 bl[443] br[443] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_444 bl[444] br[444] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_445 bl[445] br[445] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_446 bl[446] br[446] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_447 bl[447] br[447] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_448 bl[448] br[448] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_449 bl[449] br[449] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_450 bl[450] br[450] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_451 bl[451] br[451] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_452 bl[452] br[452] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_453 bl[453] br[453] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_454 bl[454] br[454] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_455 bl[455] br[455] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_456 bl[456] br[456] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_457 bl[457] br[457] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_458 bl[458] br[458] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_459 bl[459] br[459] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_460 bl[460] br[460] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_461 bl[461] br[461] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_462 bl[462] br[462] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_463 bl[463] br[463] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_464 bl[464] br[464] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_465 bl[465] br[465] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_466 bl[466] br[466] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_467 bl[467] br[467] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_468 bl[468] br[468] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_469 bl[469] br[469] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_470 bl[470] br[470] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_471 bl[471] br[471] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_472 bl[472] br[472] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_473 bl[473] br[473] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_474 bl[474] br[474] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_475 bl[475] br[475] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_476 bl[476] br[476] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_477 bl[477] br[477] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_478 bl[478] br[478] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_479 bl[479] br[479] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_480 bl[480] br[480] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_481 bl[481] br[481] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_482 bl[482] br[482] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_483 bl[483] br[483] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_484 bl[484] br[484] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_485 bl[485] br[485] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_486 bl[486] br[486] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_487 bl[487] br[487] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_488 bl[488] br[488] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_489 bl[489] br[489] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_490 bl[490] br[490] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_491 bl[491] br[491] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_492 bl[492] br[492] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_493 bl[493] br[493] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_494 bl[494] br[494] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_495 bl[495] br[495] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_496 bl[496] br[496] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_497 bl[497] br[497] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_498 bl[498] br[498] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_499 bl[499] br[499] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_500 bl[500] br[500] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_501 bl[501] br[501] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_502 bl[502] br[502] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_503 bl[503] br[503] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_504 bl[504] br[504] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_505 bl[505] br[505] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_506 bl[506] br[506] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_507 bl[507] br[507] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_508 bl[508] br[508] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_509 bl[509] br[509] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_510 bl[510] br[510] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_24_511 bl[511] br[511] vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xcell_25_0 bl[0] br[0] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_1 bl[1] br[1] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_2 bl[2] br[2] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_3 bl[3] br[3] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_4 bl[4] br[4] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_5 bl[5] br[5] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_6 bl[6] br[6] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_7 bl[7] br[7] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_8 bl[8] br[8] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_9 bl[9] br[9] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_10 bl[10] br[10] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_11 bl[11] br[11] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_12 bl[12] br[12] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_13 bl[13] br[13] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_14 bl[14] br[14] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_15 bl[15] br[15] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_16 bl[16] br[16] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_17 bl[17] br[17] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_18 bl[18] br[18] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_19 bl[19] br[19] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_20 bl[20] br[20] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_21 bl[21] br[21] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_22 bl[22] br[22] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_23 bl[23] br[23] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_24 bl[24] br[24] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_25 bl[25] br[25] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_26 bl[26] br[26] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_27 bl[27] br[27] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_28 bl[28] br[28] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_29 bl[29] br[29] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_30 bl[30] br[30] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_31 bl[31] br[31] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_32 bl[32] br[32] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_33 bl[33] br[33] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_34 bl[34] br[34] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_35 bl[35] br[35] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_36 bl[36] br[36] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_37 bl[37] br[37] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_38 bl[38] br[38] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_39 bl[39] br[39] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_40 bl[40] br[40] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_41 bl[41] br[41] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_42 bl[42] br[42] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_43 bl[43] br[43] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_44 bl[44] br[44] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_45 bl[45] br[45] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_46 bl[46] br[46] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_47 bl[47] br[47] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_48 bl[48] br[48] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_49 bl[49] br[49] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_50 bl[50] br[50] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_51 bl[51] br[51] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_52 bl[52] br[52] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_53 bl[53] br[53] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_54 bl[54] br[54] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_55 bl[55] br[55] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_56 bl[56] br[56] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_57 bl[57] br[57] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_58 bl[58] br[58] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_59 bl[59] br[59] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_60 bl[60] br[60] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_61 bl[61] br[61] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_62 bl[62] br[62] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_63 bl[63] br[63] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_64 bl[64] br[64] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_65 bl[65] br[65] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_66 bl[66] br[66] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_67 bl[67] br[67] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_68 bl[68] br[68] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_69 bl[69] br[69] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_70 bl[70] br[70] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_71 bl[71] br[71] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_72 bl[72] br[72] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_73 bl[73] br[73] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_74 bl[74] br[74] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_75 bl[75] br[75] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_76 bl[76] br[76] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_77 bl[77] br[77] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_78 bl[78] br[78] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_79 bl[79] br[79] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_80 bl[80] br[80] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_81 bl[81] br[81] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_82 bl[82] br[82] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_83 bl[83] br[83] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_84 bl[84] br[84] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_85 bl[85] br[85] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_86 bl[86] br[86] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_87 bl[87] br[87] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_88 bl[88] br[88] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_89 bl[89] br[89] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_90 bl[90] br[90] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_91 bl[91] br[91] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_92 bl[92] br[92] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_93 bl[93] br[93] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_94 bl[94] br[94] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_95 bl[95] br[95] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_96 bl[96] br[96] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_97 bl[97] br[97] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_98 bl[98] br[98] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_99 bl[99] br[99] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_100 bl[100] br[100] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_101 bl[101] br[101] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_102 bl[102] br[102] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_103 bl[103] br[103] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_104 bl[104] br[104] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_105 bl[105] br[105] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_106 bl[106] br[106] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_107 bl[107] br[107] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_108 bl[108] br[108] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_109 bl[109] br[109] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_110 bl[110] br[110] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_111 bl[111] br[111] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_112 bl[112] br[112] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_113 bl[113] br[113] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_114 bl[114] br[114] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_115 bl[115] br[115] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_116 bl[116] br[116] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_117 bl[117] br[117] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_118 bl[118] br[118] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_119 bl[119] br[119] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_120 bl[120] br[120] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_121 bl[121] br[121] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_122 bl[122] br[122] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_123 bl[123] br[123] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_124 bl[124] br[124] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_125 bl[125] br[125] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_126 bl[126] br[126] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_127 bl[127] br[127] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_128 bl[128] br[128] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_129 bl[129] br[129] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_130 bl[130] br[130] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_131 bl[131] br[131] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_132 bl[132] br[132] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_133 bl[133] br[133] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_134 bl[134] br[134] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_135 bl[135] br[135] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_136 bl[136] br[136] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_137 bl[137] br[137] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_138 bl[138] br[138] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_139 bl[139] br[139] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_140 bl[140] br[140] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_141 bl[141] br[141] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_142 bl[142] br[142] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_143 bl[143] br[143] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_144 bl[144] br[144] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_145 bl[145] br[145] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_146 bl[146] br[146] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_147 bl[147] br[147] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_148 bl[148] br[148] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_149 bl[149] br[149] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_150 bl[150] br[150] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_151 bl[151] br[151] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_152 bl[152] br[152] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_153 bl[153] br[153] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_154 bl[154] br[154] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_155 bl[155] br[155] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_156 bl[156] br[156] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_157 bl[157] br[157] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_158 bl[158] br[158] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_159 bl[159] br[159] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_160 bl[160] br[160] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_161 bl[161] br[161] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_162 bl[162] br[162] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_163 bl[163] br[163] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_164 bl[164] br[164] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_165 bl[165] br[165] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_166 bl[166] br[166] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_167 bl[167] br[167] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_168 bl[168] br[168] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_169 bl[169] br[169] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_170 bl[170] br[170] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_171 bl[171] br[171] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_172 bl[172] br[172] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_173 bl[173] br[173] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_174 bl[174] br[174] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_175 bl[175] br[175] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_176 bl[176] br[176] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_177 bl[177] br[177] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_178 bl[178] br[178] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_179 bl[179] br[179] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_180 bl[180] br[180] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_181 bl[181] br[181] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_182 bl[182] br[182] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_183 bl[183] br[183] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_184 bl[184] br[184] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_185 bl[185] br[185] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_186 bl[186] br[186] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_187 bl[187] br[187] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_188 bl[188] br[188] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_189 bl[189] br[189] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_190 bl[190] br[190] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_191 bl[191] br[191] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_192 bl[192] br[192] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_193 bl[193] br[193] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_194 bl[194] br[194] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_195 bl[195] br[195] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_196 bl[196] br[196] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_197 bl[197] br[197] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_198 bl[198] br[198] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_199 bl[199] br[199] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_200 bl[200] br[200] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_201 bl[201] br[201] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_202 bl[202] br[202] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_203 bl[203] br[203] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_204 bl[204] br[204] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_205 bl[205] br[205] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_206 bl[206] br[206] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_207 bl[207] br[207] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_208 bl[208] br[208] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_209 bl[209] br[209] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_210 bl[210] br[210] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_211 bl[211] br[211] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_212 bl[212] br[212] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_213 bl[213] br[213] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_214 bl[214] br[214] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_215 bl[215] br[215] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_216 bl[216] br[216] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_217 bl[217] br[217] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_218 bl[218] br[218] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_219 bl[219] br[219] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_220 bl[220] br[220] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_221 bl[221] br[221] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_222 bl[222] br[222] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_223 bl[223] br[223] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_224 bl[224] br[224] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_225 bl[225] br[225] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_226 bl[226] br[226] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_227 bl[227] br[227] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_228 bl[228] br[228] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_229 bl[229] br[229] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_230 bl[230] br[230] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_231 bl[231] br[231] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_232 bl[232] br[232] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_233 bl[233] br[233] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_234 bl[234] br[234] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_235 bl[235] br[235] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_236 bl[236] br[236] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_237 bl[237] br[237] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_238 bl[238] br[238] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_239 bl[239] br[239] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_240 bl[240] br[240] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_241 bl[241] br[241] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_242 bl[242] br[242] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_243 bl[243] br[243] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_244 bl[244] br[244] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_245 bl[245] br[245] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_246 bl[246] br[246] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_247 bl[247] br[247] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_248 bl[248] br[248] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_249 bl[249] br[249] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_250 bl[250] br[250] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_251 bl[251] br[251] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_252 bl[252] br[252] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_253 bl[253] br[253] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_254 bl[254] br[254] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_255 bl[255] br[255] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_256 bl[256] br[256] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_257 bl[257] br[257] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_258 bl[258] br[258] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_259 bl[259] br[259] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_260 bl[260] br[260] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_261 bl[261] br[261] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_262 bl[262] br[262] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_263 bl[263] br[263] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_264 bl[264] br[264] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_265 bl[265] br[265] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_266 bl[266] br[266] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_267 bl[267] br[267] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_268 bl[268] br[268] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_269 bl[269] br[269] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_270 bl[270] br[270] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_271 bl[271] br[271] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_272 bl[272] br[272] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_273 bl[273] br[273] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_274 bl[274] br[274] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_275 bl[275] br[275] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_276 bl[276] br[276] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_277 bl[277] br[277] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_278 bl[278] br[278] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_279 bl[279] br[279] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_280 bl[280] br[280] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_281 bl[281] br[281] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_282 bl[282] br[282] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_283 bl[283] br[283] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_284 bl[284] br[284] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_285 bl[285] br[285] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_286 bl[286] br[286] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_287 bl[287] br[287] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_288 bl[288] br[288] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_289 bl[289] br[289] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_290 bl[290] br[290] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_291 bl[291] br[291] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_292 bl[292] br[292] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_293 bl[293] br[293] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_294 bl[294] br[294] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_295 bl[295] br[295] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_296 bl[296] br[296] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_297 bl[297] br[297] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_298 bl[298] br[298] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_299 bl[299] br[299] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_300 bl[300] br[300] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_301 bl[301] br[301] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_302 bl[302] br[302] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_303 bl[303] br[303] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_304 bl[304] br[304] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_305 bl[305] br[305] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_306 bl[306] br[306] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_307 bl[307] br[307] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_308 bl[308] br[308] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_309 bl[309] br[309] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_310 bl[310] br[310] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_311 bl[311] br[311] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_312 bl[312] br[312] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_313 bl[313] br[313] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_314 bl[314] br[314] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_315 bl[315] br[315] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_316 bl[316] br[316] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_317 bl[317] br[317] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_318 bl[318] br[318] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_319 bl[319] br[319] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_320 bl[320] br[320] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_321 bl[321] br[321] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_322 bl[322] br[322] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_323 bl[323] br[323] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_324 bl[324] br[324] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_325 bl[325] br[325] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_326 bl[326] br[326] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_327 bl[327] br[327] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_328 bl[328] br[328] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_329 bl[329] br[329] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_330 bl[330] br[330] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_331 bl[331] br[331] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_332 bl[332] br[332] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_333 bl[333] br[333] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_334 bl[334] br[334] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_335 bl[335] br[335] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_336 bl[336] br[336] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_337 bl[337] br[337] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_338 bl[338] br[338] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_339 bl[339] br[339] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_340 bl[340] br[340] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_341 bl[341] br[341] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_342 bl[342] br[342] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_343 bl[343] br[343] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_344 bl[344] br[344] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_345 bl[345] br[345] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_346 bl[346] br[346] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_347 bl[347] br[347] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_348 bl[348] br[348] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_349 bl[349] br[349] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_350 bl[350] br[350] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_351 bl[351] br[351] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_352 bl[352] br[352] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_353 bl[353] br[353] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_354 bl[354] br[354] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_355 bl[355] br[355] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_356 bl[356] br[356] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_357 bl[357] br[357] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_358 bl[358] br[358] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_359 bl[359] br[359] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_360 bl[360] br[360] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_361 bl[361] br[361] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_362 bl[362] br[362] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_363 bl[363] br[363] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_364 bl[364] br[364] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_365 bl[365] br[365] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_366 bl[366] br[366] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_367 bl[367] br[367] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_368 bl[368] br[368] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_369 bl[369] br[369] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_370 bl[370] br[370] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_371 bl[371] br[371] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_372 bl[372] br[372] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_373 bl[373] br[373] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_374 bl[374] br[374] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_375 bl[375] br[375] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_376 bl[376] br[376] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_377 bl[377] br[377] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_378 bl[378] br[378] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_379 bl[379] br[379] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_380 bl[380] br[380] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_381 bl[381] br[381] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_382 bl[382] br[382] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_383 bl[383] br[383] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_384 bl[384] br[384] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_385 bl[385] br[385] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_386 bl[386] br[386] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_387 bl[387] br[387] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_388 bl[388] br[388] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_389 bl[389] br[389] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_390 bl[390] br[390] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_391 bl[391] br[391] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_392 bl[392] br[392] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_393 bl[393] br[393] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_394 bl[394] br[394] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_395 bl[395] br[395] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_396 bl[396] br[396] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_397 bl[397] br[397] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_398 bl[398] br[398] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_399 bl[399] br[399] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_400 bl[400] br[400] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_401 bl[401] br[401] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_402 bl[402] br[402] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_403 bl[403] br[403] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_404 bl[404] br[404] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_405 bl[405] br[405] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_406 bl[406] br[406] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_407 bl[407] br[407] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_408 bl[408] br[408] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_409 bl[409] br[409] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_410 bl[410] br[410] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_411 bl[411] br[411] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_412 bl[412] br[412] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_413 bl[413] br[413] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_414 bl[414] br[414] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_415 bl[415] br[415] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_416 bl[416] br[416] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_417 bl[417] br[417] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_418 bl[418] br[418] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_419 bl[419] br[419] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_420 bl[420] br[420] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_421 bl[421] br[421] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_422 bl[422] br[422] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_423 bl[423] br[423] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_424 bl[424] br[424] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_425 bl[425] br[425] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_426 bl[426] br[426] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_427 bl[427] br[427] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_428 bl[428] br[428] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_429 bl[429] br[429] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_430 bl[430] br[430] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_431 bl[431] br[431] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_432 bl[432] br[432] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_433 bl[433] br[433] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_434 bl[434] br[434] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_435 bl[435] br[435] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_436 bl[436] br[436] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_437 bl[437] br[437] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_438 bl[438] br[438] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_439 bl[439] br[439] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_440 bl[440] br[440] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_441 bl[441] br[441] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_442 bl[442] br[442] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_443 bl[443] br[443] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_444 bl[444] br[444] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_445 bl[445] br[445] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_446 bl[446] br[446] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_447 bl[447] br[447] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_448 bl[448] br[448] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_449 bl[449] br[449] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_450 bl[450] br[450] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_451 bl[451] br[451] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_452 bl[452] br[452] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_453 bl[453] br[453] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_454 bl[454] br[454] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_455 bl[455] br[455] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_456 bl[456] br[456] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_457 bl[457] br[457] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_458 bl[458] br[458] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_459 bl[459] br[459] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_460 bl[460] br[460] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_461 bl[461] br[461] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_462 bl[462] br[462] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_463 bl[463] br[463] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_464 bl[464] br[464] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_465 bl[465] br[465] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_466 bl[466] br[466] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_467 bl[467] br[467] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_468 bl[468] br[468] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_469 bl[469] br[469] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_470 bl[470] br[470] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_471 bl[471] br[471] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_472 bl[472] br[472] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_473 bl[473] br[473] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_474 bl[474] br[474] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_475 bl[475] br[475] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_476 bl[476] br[476] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_477 bl[477] br[477] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_478 bl[478] br[478] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_479 bl[479] br[479] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_480 bl[480] br[480] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_481 bl[481] br[481] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_482 bl[482] br[482] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_483 bl[483] br[483] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_484 bl[484] br[484] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_485 bl[485] br[485] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_486 bl[486] br[486] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_487 bl[487] br[487] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_488 bl[488] br[488] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_489 bl[489] br[489] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_490 bl[490] br[490] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_491 bl[491] br[491] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_492 bl[492] br[492] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_493 bl[493] br[493] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_494 bl[494] br[494] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_495 bl[495] br[495] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_496 bl[496] br[496] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_497 bl[497] br[497] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_498 bl[498] br[498] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_499 bl[499] br[499] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_500 bl[500] br[500] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_501 bl[501] br[501] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_502 bl[502] br[502] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_503 bl[503] br[503] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_504 bl[504] br[504] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_505 bl[505] br[505] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_506 bl[506] br[506] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_507 bl[507] br[507] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_508 bl[508] br[508] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_509 bl[509] br[509] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_510 bl[510] br[510] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_25_511 bl[511] br[511] vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xcell_26_0 bl[0] br[0] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_1 bl[1] br[1] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_2 bl[2] br[2] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_3 bl[3] br[3] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_4 bl[4] br[4] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_5 bl[5] br[5] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_6 bl[6] br[6] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_7 bl[7] br[7] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_8 bl[8] br[8] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_9 bl[9] br[9] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_10 bl[10] br[10] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_11 bl[11] br[11] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_12 bl[12] br[12] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_13 bl[13] br[13] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_14 bl[14] br[14] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_15 bl[15] br[15] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_16 bl[16] br[16] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_17 bl[17] br[17] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_18 bl[18] br[18] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_19 bl[19] br[19] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_20 bl[20] br[20] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_21 bl[21] br[21] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_22 bl[22] br[22] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_23 bl[23] br[23] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_24 bl[24] br[24] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_25 bl[25] br[25] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_26 bl[26] br[26] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_27 bl[27] br[27] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_28 bl[28] br[28] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_29 bl[29] br[29] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_30 bl[30] br[30] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_31 bl[31] br[31] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_32 bl[32] br[32] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_33 bl[33] br[33] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_34 bl[34] br[34] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_35 bl[35] br[35] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_36 bl[36] br[36] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_37 bl[37] br[37] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_38 bl[38] br[38] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_39 bl[39] br[39] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_40 bl[40] br[40] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_41 bl[41] br[41] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_42 bl[42] br[42] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_43 bl[43] br[43] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_44 bl[44] br[44] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_45 bl[45] br[45] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_46 bl[46] br[46] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_47 bl[47] br[47] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_48 bl[48] br[48] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_49 bl[49] br[49] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_50 bl[50] br[50] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_51 bl[51] br[51] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_52 bl[52] br[52] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_53 bl[53] br[53] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_54 bl[54] br[54] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_55 bl[55] br[55] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_56 bl[56] br[56] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_57 bl[57] br[57] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_58 bl[58] br[58] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_59 bl[59] br[59] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_60 bl[60] br[60] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_61 bl[61] br[61] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_62 bl[62] br[62] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_63 bl[63] br[63] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_64 bl[64] br[64] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_65 bl[65] br[65] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_66 bl[66] br[66] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_67 bl[67] br[67] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_68 bl[68] br[68] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_69 bl[69] br[69] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_70 bl[70] br[70] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_71 bl[71] br[71] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_72 bl[72] br[72] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_73 bl[73] br[73] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_74 bl[74] br[74] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_75 bl[75] br[75] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_76 bl[76] br[76] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_77 bl[77] br[77] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_78 bl[78] br[78] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_79 bl[79] br[79] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_80 bl[80] br[80] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_81 bl[81] br[81] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_82 bl[82] br[82] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_83 bl[83] br[83] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_84 bl[84] br[84] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_85 bl[85] br[85] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_86 bl[86] br[86] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_87 bl[87] br[87] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_88 bl[88] br[88] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_89 bl[89] br[89] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_90 bl[90] br[90] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_91 bl[91] br[91] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_92 bl[92] br[92] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_93 bl[93] br[93] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_94 bl[94] br[94] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_95 bl[95] br[95] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_96 bl[96] br[96] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_97 bl[97] br[97] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_98 bl[98] br[98] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_99 bl[99] br[99] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_100 bl[100] br[100] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_101 bl[101] br[101] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_102 bl[102] br[102] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_103 bl[103] br[103] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_104 bl[104] br[104] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_105 bl[105] br[105] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_106 bl[106] br[106] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_107 bl[107] br[107] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_108 bl[108] br[108] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_109 bl[109] br[109] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_110 bl[110] br[110] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_111 bl[111] br[111] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_112 bl[112] br[112] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_113 bl[113] br[113] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_114 bl[114] br[114] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_115 bl[115] br[115] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_116 bl[116] br[116] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_117 bl[117] br[117] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_118 bl[118] br[118] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_119 bl[119] br[119] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_120 bl[120] br[120] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_121 bl[121] br[121] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_122 bl[122] br[122] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_123 bl[123] br[123] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_124 bl[124] br[124] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_125 bl[125] br[125] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_126 bl[126] br[126] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_127 bl[127] br[127] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_128 bl[128] br[128] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_129 bl[129] br[129] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_130 bl[130] br[130] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_131 bl[131] br[131] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_132 bl[132] br[132] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_133 bl[133] br[133] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_134 bl[134] br[134] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_135 bl[135] br[135] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_136 bl[136] br[136] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_137 bl[137] br[137] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_138 bl[138] br[138] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_139 bl[139] br[139] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_140 bl[140] br[140] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_141 bl[141] br[141] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_142 bl[142] br[142] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_143 bl[143] br[143] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_144 bl[144] br[144] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_145 bl[145] br[145] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_146 bl[146] br[146] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_147 bl[147] br[147] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_148 bl[148] br[148] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_149 bl[149] br[149] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_150 bl[150] br[150] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_151 bl[151] br[151] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_152 bl[152] br[152] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_153 bl[153] br[153] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_154 bl[154] br[154] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_155 bl[155] br[155] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_156 bl[156] br[156] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_157 bl[157] br[157] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_158 bl[158] br[158] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_159 bl[159] br[159] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_160 bl[160] br[160] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_161 bl[161] br[161] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_162 bl[162] br[162] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_163 bl[163] br[163] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_164 bl[164] br[164] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_165 bl[165] br[165] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_166 bl[166] br[166] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_167 bl[167] br[167] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_168 bl[168] br[168] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_169 bl[169] br[169] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_170 bl[170] br[170] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_171 bl[171] br[171] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_172 bl[172] br[172] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_173 bl[173] br[173] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_174 bl[174] br[174] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_175 bl[175] br[175] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_176 bl[176] br[176] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_177 bl[177] br[177] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_178 bl[178] br[178] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_179 bl[179] br[179] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_180 bl[180] br[180] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_181 bl[181] br[181] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_182 bl[182] br[182] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_183 bl[183] br[183] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_184 bl[184] br[184] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_185 bl[185] br[185] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_186 bl[186] br[186] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_187 bl[187] br[187] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_188 bl[188] br[188] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_189 bl[189] br[189] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_190 bl[190] br[190] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_191 bl[191] br[191] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_192 bl[192] br[192] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_193 bl[193] br[193] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_194 bl[194] br[194] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_195 bl[195] br[195] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_196 bl[196] br[196] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_197 bl[197] br[197] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_198 bl[198] br[198] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_199 bl[199] br[199] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_200 bl[200] br[200] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_201 bl[201] br[201] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_202 bl[202] br[202] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_203 bl[203] br[203] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_204 bl[204] br[204] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_205 bl[205] br[205] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_206 bl[206] br[206] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_207 bl[207] br[207] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_208 bl[208] br[208] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_209 bl[209] br[209] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_210 bl[210] br[210] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_211 bl[211] br[211] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_212 bl[212] br[212] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_213 bl[213] br[213] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_214 bl[214] br[214] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_215 bl[215] br[215] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_216 bl[216] br[216] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_217 bl[217] br[217] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_218 bl[218] br[218] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_219 bl[219] br[219] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_220 bl[220] br[220] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_221 bl[221] br[221] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_222 bl[222] br[222] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_223 bl[223] br[223] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_224 bl[224] br[224] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_225 bl[225] br[225] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_226 bl[226] br[226] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_227 bl[227] br[227] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_228 bl[228] br[228] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_229 bl[229] br[229] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_230 bl[230] br[230] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_231 bl[231] br[231] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_232 bl[232] br[232] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_233 bl[233] br[233] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_234 bl[234] br[234] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_235 bl[235] br[235] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_236 bl[236] br[236] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_237 bl[237] br[237] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_238 bl[238] br[238] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_239 bl[239] br[239] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_240 bl[240] br[240] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_241 bl[241] br[241] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_242 bl[242] br[242] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_243 bl[243] br[243] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_244 bl[244] br[244] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_245 bl[245] br[245] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_246 bl[246] br[246] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_247 bl[247] br[247] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_248 bl[248] br[248] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_249 bl[249] br[249] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_250 bl[250] br[250] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_251 bl[251] br[251] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_252 bl[252] br[252] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_253 bl[253] br[253] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_254 bl[254] br[254] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_255 bl[255] br[255] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_256 bl[256] br[256] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_257 bl[257] br[257] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_258 bl[258] br[258] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_259 bl[259] br[259] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_260 bl[260] br[260] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_261 bl[261] br[261] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_262 bl[262] br[262] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_263 bl[263] br[263] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_264 bl[264] br[264] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_265 bl[265] br[265] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_266 bl[266] br[266] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_267 bl[267] br[267] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_268 bl[268] br[268] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_269 bl[269] br[269] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_270 bl[270] br[270] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_271 bl[271] br[271] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_272 bl[272] br[272] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_273 bl[273] br[273] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_274 bl[274] br[274] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_275 bl[275] br[275] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_276 bl[276] br[276] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_277 bl[277] br[277] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_278 bl[278] br[278] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_279 bl[279] br[279] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_280 bl[280] br[280] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_281 bl[281] br[281] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_282 bl[282] br[282] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_283 bl[283] br[283] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_284 bl[284] br[284] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_285 bl[285] br[285] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_286 bl[286] br[286] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_287 bl[287] br[287] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_288 bl[288] br[288] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_289 bl[289] br[289] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_290 bl[290] br[290] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_291 bl[291] br[291] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_292 bl[292] br[292] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_293 bl[293] br[293] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_294 bl[294] br[294] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_295 bl[295] br[295] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_296 bl[296] br[296] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_297 bl[297] br[297] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_298 bl[298] br[298] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_299 bl[299] br[299] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_300 bl[300] br[300] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_301 bl[301] br[301] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_302 bl[302] br[302] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_303 bl[303] br[303] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_304 bl[304] br[304] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_305 bl[305] br[305] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_306 bl[306] br[306] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_307 bl[307] br[307] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_308 bl[308] br[308] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_309 bl[309] br[309] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_310 bl[310] br[310] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_311 bl[311] br[311] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_312 bl[312] br[312] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_313 bl[313] br[313] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_314 bl[314] br[314] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_315 bl[315] br[315] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_316 bl[316] br[316] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_317 bl[317] br[317] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_318 bl[318] br[318] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_319 bl[319] br[319] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_320 bl[320] br[320] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_321 bl[321] br[321] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_322 bl[322] br[322] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_323 bl[323] br[323] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_324 bl[324] br[324] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_325 bl[325] br[325] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_326 bl[326] br[326] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_327 bl[327] br[327] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_328 bl[328] br[328] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_329 bl[329] br[329] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_330 bl[330] br[330] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_331 bl[331] br[331] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_332 bl[332] br[332] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_333 bl[333] br[333] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_334 bl[334] br[334] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_335 bl[335] br[335] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_336 bl[336] br[336] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_337 bl[337] br[337] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_338 bl[338] br[338] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_339 bl[339] br[339] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_340 bl[340] br[340] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_341 bl[341] br[341] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_342 bl[342] br[342] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_343 bl[343] br[343] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_344 bl[344] br[344] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_345 bl[345] br[345] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_346 bl[346] br[346] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_347 bl[347] br[347] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_348 bl[348] br[348] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_349 bl[349] br[349] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_350 bl[350] br[350] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_351 bl[351] br[351] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_352 bl[352] br[352] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_353 bl[353] br[353] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_354 bl[354] br[354] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_355 bl[355] br[355] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_356 bl[356] br[356] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_357 bl[357] br[357] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_358 bl[358] br[358] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_359 bl[359] br[359] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_360 bl[360] br[360] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_361 bl[361] br[361] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_362 bl[362] br[362] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_363 bl[363] br[363] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_364 bl[364] br[364] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_365 bl[365] br[365] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_366 bl[366] br[366] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_367 bl[367] br[367] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_368 bl[368] br[368] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_369 bl[369] br[369] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_370 bl[370] br[370] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_371 bl[371] br[371] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_372 bl[372] br[372] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_373 bl[373] br[373] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_374 bl[374] br[374] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_375 bl[375] br[375] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_376 bl[376] br[376] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_377 bl[377] br[377] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_378 bl[378] br[378] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_379 bl[379] br[379] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_380 bl[380] br[380] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_381 bl[381] br[381] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_382 bl[382] br[382] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_383 bl[383] br[383] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_384 bl[384] br[384] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_385 bl[385] br[385] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_386 bl[386] br[386] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_387 bl[387] br[387] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_388 bl[388] br[388] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_389 bl[389] br[389] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_390 bl[390] br[390] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_391 bl[391] br[391] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_392 bl[392] br[392] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_393 bl[393] br[393] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_394 bl[394] br[394] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_395 bl[395] br[395] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_396 bl[396] br[396] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_397 bl[397] br[397] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_398 bl[398] br[398] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_399 bl[399] br[399] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_400 bl[400] br[400] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_401 bl[401] br[401] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_402 bl[402] br[402] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_403 bl[403] br[403] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_404 bl[404] br[404] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_405 bl[405] br[405] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_406 bl[406] br[406] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_407 bl[407] br[407] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_408 bl[408] br[408] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_409 bl[409] br[409] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_410 bl[410] br[410] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_411 bl[411] br[411] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_412 bl[412] br[412] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_413 bl[413] br[413] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_414 bl[414] br[414] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_415 bl[415] br[415] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_416 bl[416] br[416] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_417 bl[417] br[417] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_418 bl[418] br[418] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_419 bl[419] br[419] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_420 bl[420] br[420] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_421 bl[421] br[421] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_422 bl[422] br[422] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_423 bl[423] br[423] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_424 bl[424] br[424] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_425 bl[425] br[425] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_426 bl[426] br[426] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_427 bl[427] br[427] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_428 bl[428] br[428] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_429 bl[429] br[429] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_430 bl[430] br[430] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_431 bl[431] br[431] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_432 bl[432] br[432] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_433 bl[433] br[433] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_434 bl[434] br[434] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_435 bl[435] br[435] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_436 bl[436] br[436] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_437 bl[437] br[437] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_438 bl[438] br[438] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_439 bl[439] br[439] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_440 bl[440] br[440] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_441 bl[441] br[441] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_442 bl[442] br[442] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_443 bl[443] br[443] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_444 bl[444] br[444] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_445 bl[445] br[445] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_446 bl[446] br[446] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_447 bl[447] br[447] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_448 bl[448] br[448] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_449 bl[449] br[449] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_450 bl[450] br[450] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_451 bl[451] br[451] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_452 bl[452] br[452] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_453 bl[453] br[453] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_454 bl[454] br[454] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_455 bl[455] br[455] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_456 bl[456] br[456] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_457 bl[457] br[457] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_458 bl[458] br[458] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_459 bl[459] br[459] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_460 bl[460] br[460] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_461 bl[461] br[461] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_462 bl[462] br[462] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_463 bl[463] br[463] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_464 bl[464] br[464] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_465 bl[465] br[465] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_466 bl[466] br[466] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_467 bl[467] br[467] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_468 bl[468] br[468] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_469 bl[469] br[469] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_470 bl[470] br[470] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_471 bl[471] br[471] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_472 bl[472] br[472] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_473 bl[473] br[473] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_474 bl[474] br[474] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_475 bl[475] br[475] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_476 bl[476] br[476] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_477 bl[477] br[477] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_478 bl[478] br[478] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_479 bl[479] br[479] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_480 bl[480] br[480] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_481 bl[481] br[481] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_482 bl[482] br[482] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_483 bl[483] br[483] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_484 bl[484] br[484] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_485 bl[485] br[485] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_486 bl[486] br[486] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_487 bl[487] br[487] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_488 bl[488] br[488] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_489 bl[489] br[489] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_490 bl[490] br[490] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_491 bl[491] br[491] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_492 bl[492] br[492] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_493 bl[493] br[493] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_494 bl[494] br[494] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_495 bl[495] br[495] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_496 bl[496] br[496] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_497 bl[497] br[497] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_498 bl[498] br[498] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_499 bl[499] br[499] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_500 bl[500] br[500] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_501 bl[501] br[501] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_502 bl[502] br[502] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_503 bl[503] br[503] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_504 bl[504] br[504] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_505 bl[505] br[505] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_506 bl[506] br[506] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_507 bl[507] br[507] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_508 bl[508] br[508] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_509 bl[509] br[509] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_510 bl[510] br[510] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_26_511 bl[511] br[511] vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xcell_27_0 bl[0] br[0] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_1 bl[1] br[1] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_2 bl[2] br[2] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_3 bl[3] br[3] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_4 bl[4] br[4] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_5 bl[5] br[5] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_6 bl[6] br[6] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_7 bl[7] br[7] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_8 bl[8] br[8] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_9 bl[9] br[9] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_10 bl[10] br[10] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_11 bl[11] br[11] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_12 bl[12] br[12] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_13 bl[13] br[13] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_14 bl[14] br[14] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_15 bl[15] br[15] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_16 bl[16] br[16] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_17 bl[17] br[17] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_18 bl[18] br[18] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_19 bl[19] br[19] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_20 bl[20] br[20] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_21 bl[21] br[21] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_22 bl[22] br[22] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_23 bl[23] br[23] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_24 bl[24] br[24] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_25 bl[25] br[25] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_26 bl[26] br[26] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_27 bl[27] br[27] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_28 bl[28] br[28] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_29 bl[29] br[29] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_30 bl[30] br[30] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_31 bl[31] br[31] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_32 bl[32] br[32] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_33 bl[33] br[33] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_34 bl[34] br[34] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_35 bl[35] br[35] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_36 bl[36] br[36] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_37 bl[37] br[37] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_38 bl[38] br[38] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_39 bl[39] br[39] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_40 bl[40] br[40] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_41 bl[41] br[41] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_42 bl[42] br[42] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_43 bl[43] br[43] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_44 bl[44] br[44] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_45 bl[45] br[45] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_46 bl[46] br[46] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_47 bl[47] br[47] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_48 bl[48] br[48] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_49 bl[49] br[49] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_50 bl[50] br[50] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_51 bl[51] br[51] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_52 bl[52] br[52] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_53 bl[53] br[53] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_54 bl[54] br[54] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_55 bl[55] br[55] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_56 bl[56] br[56] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_57 bl[57] br[57] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_58 bl[58] br[58] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_59 bl[59] br[59] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_60 bl[60] br[60] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_61 bl[61] br[61] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_62 bl[62] br[62] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_63 bl[63] br[63] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_64 bl[64] br[64] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_65 bl[65] br[65] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_66 bl[66] br[66] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_67 bl[67] br[67] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_68 bl[68] br[68] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_69 bl[69] br[69] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_70 bl[70] br[70] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_71 bl[71] br[71] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_72 bl[72] br[72] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_73 bl[73] br[73] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_74 bl[74] br[74] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_75 bl[75] br[75] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_76 bl[76] br[76] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_77 bl[77] br[77] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_78 bl[78] br[78] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_79 bl[79] br[79] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_80 bl[80] br[80] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_81 bl[81] br[81] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_82 bl[82] br[82] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_83 bl[83] br[83] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_84 bl[84] br[84] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_85 bl[85] br[85] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_86 bl[86] br[86] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_87 bl[87] br[87] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_88 bl[88] br[88] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_89 bl[89] br[89] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_90 bl[90] br[90] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_91 bl[91] br[91] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_92 bl[92] br[92] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_93 bl[93] br[93] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_94 bl[94] br[94] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_95 bl[95] br[95] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_96 bl[96] br[96] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_97 bl[97] br[97] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_98 bl[98] br[98] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_99 bl[99] br[99] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_100 bl[100] br[100] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_101 bl[101] br[101] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_102 bl[102] br[102] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_103 bl[103] br[103] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_104 bl[104] br[104] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_105 bl[105] br[105] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_106 bl[106] br[106] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_107 bl[107] br[107] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_108 bl[108] br[108] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_109 bl[109] br[109] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_110 bl[110] br[110] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_111 bl[111] br[111] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_112 bl[112] br[112] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_113 bl[113] br[113] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_114 bl[114] br[114] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_115 bl[115] br[115] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_116 bl[116] br[116] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_117 bl[117] br[117] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_118 bl[118] br[118] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_119 bl[119] br[119] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_120 bl[120] br[120] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_121 bl[121] br[121] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_122 bl[122] br[122] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_123 bl[123] br[123] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_124 bl[124] br[124] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_125 bl[125] br[125] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_126 bl[126] br[126] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_127 bl[127] br[127] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_128 bl[128] br[128] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_129 bl[129] br[129] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_130 bl[130] br[130] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_131 bl[131] br[131] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_132 bl[132] br[132] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_133 bl[133] br[133] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_134 bl[134] br[134] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_135 bl[135] br[135] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_136 bl[136] br[136] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_137 bl[137] br[137] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_138 bl[138] br[138] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_139 bl[139] br[139] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_140 bl[140] br[140] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_141 bl[141] br[141] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_142 bl[142] br[142] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_143 bl[143] br[143] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_144 bl[144] br[144] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_145 bl[145] br[145] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_146 bl[146] br[146] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_147 bl[147] br[147] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_148 bl[148] br[148] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_149 bl[149] br[149] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_150 bl[150] br[150] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_151 bl[151] br[151] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_152 bl[152] br[152] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_153 bl[153] br[153] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_154 bl[154] br[154] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_155 bl[155] br[155] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_156 bl[156] br[156] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_157 bl[157] br[157] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_158 bl[158] br[158] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_159 bl[159] br[159] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_160 bl[160] br[160] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_161 bl[161] br[161] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_162 bl[162] br[162] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_163 bl[163] br[163] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_164 bl[164] br[164] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_165 bl[165] br[165] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_166 bl[166] br[166] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_167 bl[167] br[167] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_168 bl[168] br[168] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_169 bl[169] br[169] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_170 bl[170] br[170] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_171 bl[171] br[171] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_172 bl[172] br[172] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_173 bl[173] br[173] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_174 bl[174] br[174] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_175 bl[175] br[175] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_176 bl[176] br[176] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_177 bl[177] br[177] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_178 bl[178] br[178] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_179 bl[179] br[179] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_180 bl[180] br[180] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_181 bl[181] br[181] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_182 bl[182] br[182] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_183 bl[183] br[183] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_184 bl[184] br[184] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_185 bl[185] br[185] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_186 bl[186] br[186] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_187 bl[187] br[187] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_188 bl[188] br[188] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_189 bl[189] br[189] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_190 bl[190] br[190] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_191 bl[191] br[191] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_192 bl[192] br[192] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_193 bl[193] br[193] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_194 bl[194] br[194] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_195 bl[195] br[195] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_196 bl[196] br[196] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_197 bl[197] br[197] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_198 bl[198] br[198] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_199 bl[199] br[199] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_200 bl[200] br[200] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_201 bl[201] br[201] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_202 bl[202] br[202] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_203 bl[203] br[203] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_204 bl[204] br[204] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_205 bl[205] br[205] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_206 bl[206] br[206] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_207 bl[207] br[207] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_208 bl[208] br[208] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_209 bl[209] br[209] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_210 bl[210] br[210] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_211 bl[211] br[211] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_212 bl[212] br[212] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_213 bl[213] br[213] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_214 bl[214] br[214] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_215 bl[215] br[215] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_216 bl[216] br[216] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_217 bl[217] br[217] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_218 bl[218] br[218] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_219 bl[219] br[219] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_220 bl[220] br[220] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_221 bl[221] br[221] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_222 bl[222] br[222] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_223 bl[223] br[223] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_224 bl[224] br[224] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_225 bl[225] br[225] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_226 bl[226] br[226] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_227 bl[227] br[227] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_228 bl[228] br[228] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_229 bl[229] br[229] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_230 bl[230] br[230] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_231 bl[231] br[231] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_232 bl[232] br[232] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_233 bl[233] br[233] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_234 bl[234] br[234] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_235 bl[235] br[235] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_236 bl[236] br[236] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_237 bl[237] br[237] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_238 bl[238] br[238] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_239 bl[239] br[239] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_240 bl[240] br[240] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_241 bl[241] br[241] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_242 bl[242] br[242] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_243 bl[243] br[243] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_244 bl[244] br[244] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_245 bl[245] br[245] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_246 bl[246] br[246] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_247 bl[247] br[247] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_248 bl[248] br[248] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_249 bl[249] br[249] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_250 bl[250] br[250] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_251 bl[251] br[251] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_252 bl[252] br[252] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_253 bl[253] br[253] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_254 bl[254] br[254] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_255 bl[255] br[255] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_256 bl[256] br[256] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_257 bl[257] br[257] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_258 bl[258] br[258] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_259 bl[259] br[259] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_260 bl[260] br[260] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_261 bl[261] br[261] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_262 bl[262] br[262] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_263 bl[263] br[263] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_264 bl[264] br[264] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_265 bl[265] br[265] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_266 bl[266] br[266] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_267 bl[267] br[267] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_268 bl[268] br[268] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_269 bl[269] br[269] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_270 bl[270] br[270] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_271 bl[271] br[271] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_272 bl[272] br[272] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_273 bl[273] br[273] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_274 bl[274] br[274] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_275 bl[275] br[275] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_276 bl[276] br[276] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_277 bl[277] br[277] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_278 bl[278] br[278] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_279 bl[279] br[279] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_280 bl[280] br[280] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_281 bl[281] br[281] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_282 bl[282] br[282] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_283 bl[283] br[283] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_284 bl[284] br[284] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_285 bl[285] br[285] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_286 bl[286] br[286] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_287 bl[287] br[287] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_288 bl[288] br[288] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_289 bl[289] br[289] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_290 bl[290] br[290] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_291 bl[291] br[291] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_292 bl[292] br[292] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_293 bl[293] br[293] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_294 bl[294] br[294] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_295 bl[295] br[295] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_296 bl[296] br[296] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_297 bl[297] br[297] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_298 bl[298] br[298] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_299 bl[299] br[299] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_300 bl[300] br[300] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_301 bl[301] br[301] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_302 bl[302] br[302] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_303 bl[303] br[303] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_304 bl[304] br[304] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_305 bl[305] br[305] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_306 bl[306] br[306] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_307 bl[307] br[307] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_308 bl[308] br[308] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_309 bl[309] br[309] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_310 bl[310] br[310] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_311 bl[311] br[311] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_312 bl[312] br[312] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_313 bl[313] br[313] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_314 bl[314] br[314] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_315 bl[315] br[315] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_316 bl[316] br[316] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_317 bl[317] br[317] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_318 bl[318] br[318] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_319 bl[319] br[319] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_320 bl[320] br[320] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_321 bl[321] br[321] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_322 bl[322] br[322] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_323 bl[323] br[323] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_324 bl[324] br[324] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_325 bl[325] br[325] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_326 bl[326] br[326] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_327 bl[327] br[327] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_328 bl[328] br[328] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_329 bl[329] br[329] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_330 bl[330] br[330] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_331 bl[331] br[331] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_332 bl[332] br[332] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_333 bl[333] br[333] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_334 bl[334] br[334] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_335 bl[335] br[335] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_336 bl[336] br[336] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_337 bl[337] br[337] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_338 bl[338] br[338] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_339 bl[339] br[339] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_340 bl[340] br[340] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_341 bl[341] br[341] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_342 bl[342] br[342] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_343 bl[343] br[343] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_344 bl[344] br[344] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_345 bl[345] br[345] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_346 bl[346] br[346] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_347 bl[347] br[347] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_348 bl[348] br[348] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_349 bl[349] br[349] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_350 bl[350] br[350] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_351 bl[351] br[351] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_352 bl[352] br[352] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_353 bl[353] br[353] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_354 bl[354] br[354] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_355 bl[355] br[355] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_356 bl[356] br[356] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_357 bl[357] br[357] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_358 bl[358] br[358] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_359 bl[359] br[359] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_360 bl[360] br[360] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_361 bl[361] br[361] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_362 bl[362] br[362] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_363 bl[363] br[363] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_364 bl[364] br[364] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_365 bl[365] br[365] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_366 bl[366] br[366] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_367 bl[367] br[367] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_368 bl[368] br[368] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_369 bl[369] br[369] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_370 bl[370] br[370] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_371 bl[371] br[371] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_372 bl[372] br[372] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_373 bl[373] br[373] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_374 bl[374] br[374] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_375 bl[375] br[375] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_376 bl[376] br[376] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_377 bl[377] br[377] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_378 bl[378] br[378] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_379 bl[379] br[379] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_380 bl[380] br[380] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_381 bl[381] br[381] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_382 bl[382] br[382] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_383 bl[383] br[383] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_384 bl[384] br[384] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_385 bl[385] br[385] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_386 bl[386] br[386] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_387 bl[387] br[387] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_388 bl[388] br[388] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_389 bl[389] br[389] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_390 bl[390] br[390] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_391 bl[391] br[391] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_392 bl[392] br[392] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_393 bl[393] br[393] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_394 bl[394] br[394] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_395 bl[395] br[395] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_396 bl[396] br[396] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_397 bl[397] br[397] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_398 bl[398] br[398] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_399 bl[399] br[399] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_400 bl[400] br[400] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_401 bl[401] br[401] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_402 bl[402] br[402] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_403 bl[403] br[403] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_404 bl[404] br[404] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_405 bl[405] br[405] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_406 bl[406] br[406] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_407 bl[407] br[407] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_408 bl[408] br[408] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_409 bl[409] br[409] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_410 bl[410] br[410] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_411 bl[411] br[411] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_412 bl[412] br[412] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_413 bl[413] br[413] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_414 bl[414] br[414] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_415 bl[415] br[415] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_416 bl[416] br[416] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_417 bl[417] br[417] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_418 bl[418] br[418] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_419 bl[419] br[419] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_420 bl[420] br[420] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_421 bl[421] br[421] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_422 bl[422] br[422] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_423 bl[423] br[423] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_424 bl[424] br[424] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_425 bl[425] br[425] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_426 bl[426] br[426] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_427 bl[427] br[427] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_428 bl[428] br[428] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_429 bl[429] br[429] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_430 bl[430] br[430] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_431 bl[431] br[431] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_432 bl[432] br[432] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_433 bl[433] br[433] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_434 bl[434] br[434] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_435 bl[435] br[435] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_436 bl[436] br[436] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_437 bl[437] br[437] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_438 bl[438] br[438] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_439 bl[439] br[439] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_440 bl[440] br[440] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_441 bl[441] br[441] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_442 bl[442] br[442] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_443 bl[443] br[443] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_444 bl[444] br[444] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_445 bl[445] br[445] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_446 bl[446] br[446] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_447 bl[447] br[447] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_448 bl[448] br[448] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_449 bl[449] br[449] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_450 bl[450] br[450] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_451 bl[451] br[451] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_452 bl[452] br[452] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_453 bl[453] br[453] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_454 bl[454] br[454] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_455 bl[455] br[455] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_456 bl[456] br[456] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_457 bl[457] br[457] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_458 bl[458] br[458] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_459 bl[459] br[459] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_460 bl[460] br[460] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_461 bl[461] br[461] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_462 bl[462] br[462] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_463 bl[463] br[463] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_464 bl[464] br[464] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_465 bl[465] br[465] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_466 bl[466] br[466] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_467 bl[467] br[467] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_468 bl[468] br[468] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_469 bl[469] br[469] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_470 bl[470] br[470] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_471 bl[471] br[471] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_472 bl[472] br[472] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_473 bl[473] br[473] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_474 bl[474] br[474] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_475 bl[475] br[475] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_476 bl[476] br[476] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_477 bl[477] br[477] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_478 bl[478] br[478] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_479 bl[479] br[479] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_480 bl[480] br[480] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_481 bl[481] br[481] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_482 bl[482] br[482] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_483 bl[483] br[483] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_484 bl[484] br[484] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_485 bl[485] br[485] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_486 bl[486] br[486] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_487 bl[487] br[487] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_488 bl[488] br[488] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_489 bl[489] br[489] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_490 bl[490] br[490] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_491 bl[491] br[491] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_492 bl[492] br[492] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_493 bl[493] br[493] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_494 bl[494] br[494] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_495 bl[495] br[495] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_496 bl[496] br[496] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_497 bl[497] br[497] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_498 bl[498] br[498] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_499 bl[499] br[499] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_500 bl[500] br[500] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_501 bl[501] br[501] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_502 bl[502] br[502] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_503 bl[503] br[503] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_504 bl[504] br[504] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_505 bl[505] br[505] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_506 bl[506] br[506] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_507 bl[507] br[507] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_508 bl[508] br[508] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_509 bl[509] br[509] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_510 bl[510] br[510] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_27_511 bl[511] br[511] vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xcell_28_0 bl[0] br[0] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_1 bl[1] br[1] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_2 bl[2] br[2] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_3 bl[3] br[3] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_4 bl[4] br[4] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_5 bl[5] br[5] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_6 bl[6] br[6] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_7 bl[7] br[7] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_8 bl[8] br[8] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_9 bl[9] br[9] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_10 bl[10] br[10] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_11 bl[11] br[11] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_12 bl[12] br[12] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_13 bl[13] br[13] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_14 bl[14] br[14] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_15 bl[15] br[15] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_16 bl[16] br[16] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_17 bl[17] br[17] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_18 bl[18] br[18] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_19 bl[19] br[19] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_20 bl[20] br[20] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_21 bl[21] br[21] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_22 bl[22] br[22] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_23 bl[23] br[23] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_24 bl[24] br[24] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_25 bl[25] br[25] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_26 bl[26] br[26] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_27 bl[27] br[27] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_28 bl[28] br[28] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_29 bl[29] br[29] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_30 bl[30] br[30] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_31 bl[31] br[31] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_32 bl[32] br[32] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_33 bl[33] br[33] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_34 bl[34] br[34] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_35 bl[35] br[35] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_36 bl[36] br[36] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_37 bl[37] br[37] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_38 bl[38] br[38] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_39 bl[39] br[39] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_40 bl[40] br[40] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_41 bl[41] br[41] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_42 bl[42] br[42] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_43 bl[43] br[43] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_44 bl[44] br[44] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_45 bl[45] br[45] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_46 bl[46] br[46] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_47 bl[47] br[47] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_48 bl[48] br[48] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_49 bl[49] br[49] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_50 bl[50] br[50] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_51 bl[51] br[51] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_52 bl[52] br[52] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_53 bl[53] br[53] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_54 bl[54] br[54] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_55 bl[55] br[55] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_56 bl[56] br[56] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_57 bl[57] br[57] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_58 bl[58] br[58] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_59 bl[59] br[59] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_60 bl[60] br[60] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_61 bl[61] br[61] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_62 bl[62] br[62] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_63 bl[63] br[63] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_64 bl[64] br[64] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_65 bl[65] br[65] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_66 bl[66] br[66] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_67 bl[67] br[67] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_68 bl[68] br[68] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_69 bl[69] br[69] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_70 bl[70] br[70] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_71 bl[71] br[71] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_72 bl[72] br[72] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_73 bl[73] br[73] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_74 bl[74] br[74] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_75 bl[75] br[75] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_76 bl[76] br[76] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_77 bl[77] br[77] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_78 bl[78] br[78] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_79 bl[79] br[79] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_80 bl[80] br[80] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_81 bl[81] br[81] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_82 bl[82] br[82] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_83 bl[83] br[83] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_84 bl[84] br[84] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_85 bl[85] br[85] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_86 bl[86] br[86] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_87 bl[87] br[87] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_88 bl[88] br[88] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_89 bl[89] br[89] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_90 bl[90] br[90] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_91 bl[91] br[91] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_92 bl[92] br[92] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_93 bl[93] br[93] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_94 bl[94] br[94] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_95 bl[95] br[95] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_96 bl[96] br[96] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_97 bl[97] br[97] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_98 bl[98] br[98] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_99 bl[99] br[99] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_100 bl[100] br[100] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_101 bl[101] br[101] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_102 bl[102] br[102] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_103 bl[103] br[103] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_104 bl[104] br[104] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_105 bl[105] br[105] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_106 bl[106] br[106] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_107 bl[107] br[107] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_108 bl[108] br[108] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_109 bl[109] br[109] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_110 bl[110] br[110] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_111 bl[111] br[111] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_112 bl[112] br[112] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_113 bl[113] br[113] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_114 bl[114] br[114] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_115 bl[115] br[115] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_116 bl[116] br[116] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_117 bl[117] br[117] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_118 bl[118] br[118] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_119 bl[119] br[119] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_120 bl[120] br[120] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_121 bl[121] br[121] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_122 bl[122] br[122] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_123 bl[123] br[123] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_124 bl[124] br[124] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_125 bl[125] br[125] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_126 bl[126] br[126] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_127 bl[127] br[127] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_128 bl[128] br[128] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_129 bl[129] br[129] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_130 bl[130] br[130] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_131 bl[131] br[131] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_132 bl[132] br[132] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_133 bl[133] br[133] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_134 bl[134] br[134] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_135 bl[135] br[135] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_136 bl[136] br[136] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_137 bl[137] br[137] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_138 bl[138] br[138] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_139 bl[139] br[139] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_140 bl[140] br[140] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_141 bl[141] br[141] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_142 bl[142] br[142] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_143 bl[143] br[143] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_144 bl[144] br[144] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_145 bl[145] br[145] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_146 bl[146] br[146] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_147 bl[147] br[147] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_148 bl[148] br[148] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_149 bl[149] br[149] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_150 bl[150] br[150] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_151 bl[151] br[151] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_152 bl[152] br[152] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_153 bl[153] br[153] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_154 bl[154] br[154] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_155 bl[155] br[155] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_156 bl[156] br[156] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_157 bl[157] br[157] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_158 bl[158] br[158] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_159 bl[159] br[159] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_160 bl[160] br[160] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_161 bl[161] br[161] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_162 bl[162] br[162] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_163 bl[163] br[163] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_164 bl[164] br[164] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_165 bl[165] br[165] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_166 bl[166] br[166] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_167 bl[167] br[167] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_168 bl[168] br[168] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_169 bl[169] br[169] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_170 bl[170] br[170] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_171 bl[171] br[171] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_172 bl[172] br[172] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_173 bl[173] br[173] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_174 bl[174] br[174] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_175 bl[175] br[175] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_176 bl[176] br[176] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_177 bl[177] br[177] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_178 bl[178] br[178] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_179 bl[179] br[179] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_180 bl[180] br[180] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_181 bl[181] br[181] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_182 bl[182] br[182] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_183 bl[183] br[183] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_184 bl[184] br[184] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_185 bl[185] br[185] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_186 bl[186] br[186] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_187 bl[187] br[187] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_188 bl[188] br[188] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_189 bl[189] br[189] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_190 bl[190] br[190] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_191 bl[191] br[191] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_192 bl[192] br[192] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_193 bl[193] br[193] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_194 bl[194] br[194] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_195 bl[195] br[195] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_196 bl[196] br[196] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_197 bl[197] br[197] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_198 bl[198] br[198] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_199 bl[199] br[199] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_200 bl[200] br[200] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_201 bl[201] br[201] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_202 bl[202] br[202] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_203 bl[203] br[203] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_204 bl[204] br[204] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_205 bl[205] br[205] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_206 bl[206] br[206] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_207 bl[207] br[207] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_208 bl[208] br[208] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_209 bl[209] br[209] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_210 bl[210] br[210] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_211 bl[211] br[211] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_212 bl[212] br[212] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_213 bl[213] br[213] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_214 bl[214] br[214] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_215 bl[215] br[215] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_216 bl[216] br[216] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_217 bl[217] br[217] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_218 bl[218] br[218] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_219 bl[219] br[219] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_220 bl[220] br[220] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_221 bl[221] br[221] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_222 bl[222] br[222] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_223 bl[223] br[223] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_224 bl[224] br[224] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_225 bl[225] br[225] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_226 bl[226] br[226] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_227 bl[227] br[227] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_228 bl[228] br[228] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_229 bl[229] br[229] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_230 bl[230] br[230] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_231 bl[231] br[231] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_232 bl[232] br[232] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_233 bl[233] br[233] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_234 bl[234] br[234] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_235 bl[235] br[235] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_236 bl[236] br[236] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_237 bl[237] br[237] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_238 bl[238] br[238] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_239 bl[239] br[239] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_240 bl[240] br[240] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_241 bl[241] br[241] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_242 bl[242] br[242] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_243 bl[243] br[243] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_244 bl[244] br[244] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_245 bl[245] br[245] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_246 bl[246] br[246] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_247 bl[247] br[247] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_248 bl[248] br[248] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_249 bl[249] br[249] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_250 bl[250] br[250] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_251 bl[251] br[251] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_252 bl[252] br[252] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_253 bl[253] br[253] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_254 bl[254] br[254] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_255 bl[255] br[255] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_256 bl[256] br[256] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_257 bl[257] br[257] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_258 bl[258] br[258] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_259 bl[259] br[259] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_260 bl[260] br[260] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_261 bl[261] br[261] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_262 bl[262] br[262] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_263 bl[263] br[263] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_264 bl[264] br[264] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_265 bl[265] br[265] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_266 bl[266] br[266] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_267 bl[267] br[267] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_268 bl[268] br[268] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_269 bl[269] br[269] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_270 bl[270] br[270] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_271 bl[271] br[271] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_272 bl[272] br[272] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_273 bl[273] br[273] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_274 bl[274] br[274] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_275 bl[275] br[275] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_276 bl[276] br[276] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_277 bl[277] br[277] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_278 bl[278] br[278] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_279 bl[279] br[279] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_280 bl[280] br[280] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_281 bl[281] br[281] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_282 bl[282] br[282] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_283 bl[283] br[283] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_284 bl[284] br[284] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_285 bl[285] br[285] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_286 bl[286] br[286] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_287 bl[287] br[287] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_288 bl[288] br[288] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_289 bl[289] br[289] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_290 bl[290] br[290] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_291 bl[291] br[291] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_292 bl[292] br[292] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_293 bl[293] br[293] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_294 bl[294] br[294] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_295 bl[295] br[295] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_296 bl[296] br[296] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_297 bl[297] br[297] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_298 bl[298] br[298] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_299 bl[299] br[299] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_300 bl[300] br[300] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_301 bl[301] br[301] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_302 bl[302] br[302] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_303 bl[303] br[303] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_304 bl[304] br[304] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_305 bl[305] br[305] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_306 bl[306] br[306] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_307 bl[307] br[307] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_308 bl[308] br[308] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_309 bl[309] br[309] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_310 bl[310] br[310] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_311 bl[311] br[311] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_312 bl[312] br[312] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_313 bl[313] br[313] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_314 bl[314] br[314] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_315 bl[315] br[315] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_316 bl[316] br[316] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_317 bl[317] br[317] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_318 bl[318] br[318] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_319 bl[319] br[319] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_320 bl[320] br[320] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_321 bl[321] br[321] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_322 bl[322] br[322] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_323 bl[323] br[323] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_324 bl[324] br[324] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_325 bl[325] br[325] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_326 bl[326] br[326] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_327 bl[327] br[327] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_328 bl[328] br[328] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_329 bl[329] br[329] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_330 bl[330] br[330] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_331 bl[331] br[331] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_332 bl[332] br[332] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_333 bl[333] br[333] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_334 bl[334] br[334] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_335 bl[335] br[335] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_336 bl[336] br[336] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_337 bl[337] br[337] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_338 bl[338] br[338] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_339 bl[339] br[339] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_340 bl[340] br[340] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_341 bl[341] br[341] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_342 bl[342] br[342] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_343 bl[343] br[343] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_344 bl[344] br[344] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_345 bl[345] br[345] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_346 bl[346] br[346] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_347 bl[347] br[347] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_348 bl[348] br[348] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_349 bl[349] br[349] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_350 bl[350] br[350] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_351 bl[351] br[351] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_352 bl[352] br[352] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_353 bl[353] br[353] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_354 bl[354] br[354] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_355 bl[355] br[355] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_356 bl[356] br[356] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_357 bl[357] br[357] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_358 bl[358] br[358] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_359 bl[359] br[359] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_360 bl[360] br[360] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_361 bl[361] br[361] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_362 bl[362] br[362] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_363 bl[363] br[363] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_364 bl[364] br[364] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_365 bl[365] br[365] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_366 bl[366] br[366] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_367 bl[367] br[367] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_368 bl[368] br[368] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_369 bl[369] br[369] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_370 bl[370] br[370] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_371 bl[371] br[371] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_372 bl[372] br[372] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_373 bl[373] br[373] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_374 bl[374] br[374] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_375 bl[375] br[375] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_376 bl[376] br[376] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_377 bl[377] br[377] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_378 bl[378] br[378] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_379 bl[379] br[379] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_380 bl[380] br[380] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_381 bl[381] br[381] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_382 bl[382] br[382] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_383 bl[383] br[383] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_384 bl[384] br[384] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_385 bl[385] br[385] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_386 bl[386] br[386] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_387 bl[387] br[387] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_388 bl[388] br[388] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_389 bl[389] br[389] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_390 bl[390] br[390] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_391 bl[391] br[391] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_392 bl[392] br[392] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_393 bl[393] br[393] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_394 bl[394] br[394] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_395 bl[395] br[395] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_396 bl[396] br[396] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_397 bl[397] br[397] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_398 bl[398] br[398] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_399 bl[399] br[399] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_400 bl[400] br[400] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_401 bl[401] br[401] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_402 bl[402] br[402] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_403 bl[403] br[403] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_404 bl[404] br[404] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_405 bl[405] br[405] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_406 bl[406] br[406] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_407 bl[407] br[407] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_408 bl[408] br[408] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_409 bl[409] br[409] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_410 bl[410] br[410] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_411 bl[411] br[411] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_412 bl[412] br[412] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_413 bl[413] br[413] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_414 bl[414] br[414] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_415 bl[415] br[415] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_416 bl[416] br[416] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_417 bl[417] br[417] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_418 bl[418] br[418] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_419 bl[419] br[419] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_420 bl[420] br[420] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_421 bl[421] br[421] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_422 bl[422] br[422] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_423 bl[423] br[423] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_424 bl[424] br[424] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_425 bl[425] br[425] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_426 bl[426] br[426] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_427 bl[427] br[427] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_428 bl[428] br[428] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_429 bl[429] br[429] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_430 bl[430] br[430] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_431 bl[431] br[431] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_432 bl[432] br[432] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_433 bl[433] br[433] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_434 bl[434] br[434] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_435 bl[435] br[435] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_436 bl[436] br[436] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_437 bl[437] br[437] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_438 bl[438] br[438] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_439 bl[439] br[439] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_440 bl[440] br[440] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_441 bl[441] br[441] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_442 bl[442] br[442] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_443 bl[443] br[443] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_444 bl[444] br[444] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_445 bl[445] br[445] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_446 bl[446] br[446] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_447 bl[447] br[447] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_448 bl[448] br[448] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_449 bl[449] br[449] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_450 bl[450] br[450] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_451 bl[451] br[451] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_452 bl[452] br[452] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_453 bl[453] br[453] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_454 bl[454] br[454] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_455 bl[455] br[455] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_456 bl[456] br[456] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_457 bl[457] br[457] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_458 bl[458] br[458] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_459 bl[459] br[459] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_460 bl[460] br[460] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_461 bl[461] br[461] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_462 bl[462] br[462] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_463 bl[463] br[463] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_464 bl[464] br[464] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_465 bl[465] br[465] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_466 bl[466] br[466] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_467 bl[467] br[467] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_468 bl[468] br[468] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_469 bl[469] br[469] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_470 bl[470] br[470] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_471 bl[471] br[471] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_472 bl[472] br[472] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_473 bl[473] br[473] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_474 bl[474] br[474] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_475 bl[475] br[475] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_476 bl[476] br[476] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_477 bl[477] br[477] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_478 bl[478] br[478] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_479 bl[479] br[479] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_480 bl[480] br[480] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_481 bl[481] br[481] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_482 bl[482] br[482] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_483 bl[483] br[483] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_484 bl[484] br[484] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_485 bl[485] br[485] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_486 bl[486] br[486] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_487 bl[487] br[487] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_488 bl[488] br[488] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_489 bl[489] br[489] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_490 bl[490] br[490] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_491 bl[491] br[491] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_492 bl[492] br[492] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_493 bl[493] br[493] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_494 bl[494] br[494] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_495 bl[495] br[495] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_496 bl[496] br[496] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_497 bl[497] br[497] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_498 bl[498] br[498] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_499 bl[499] br[499] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_500 bl[500] br[500] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_501 bl[501] br[501] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_502 bl[502] br[502] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_503 bl[503] br[503] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_504 bl[504] br[504] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_505 bl[505] br[505] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_506 bl[506] br[506] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_507 bl[507] br[507] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_508 bl[508] br[508] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_509 bl[509] br[509] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_510 bl[510] br[510] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_28_511 bl[511] br[511] vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xcell_29_0 bl[0] br[0] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_1 bl[1] br[1] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_2 bl[2] br[2] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_3 bl[3] br[3] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_4 bl[4] br[4] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_5 bl[5] br[5] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_6 bl[6] br[6] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_7 bl[7] br[7] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_8 bl[8] br[8] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_9 bl[9] br[9] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_10 bl[10] br[10] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_11 bl[11] br[11] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_12 bl[12] br[12] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_13 bl[13] br[13] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_14 bl[14] br[14] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_15 bl[15] br[15] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_16 bl[16] br[16] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_17 bl[17] br[17] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_18 bl[18] br[18] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_19 bl[19] br[19] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_20 bl[20] br[20] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_21 bl[21] br[21] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_22 bl[22] br[22] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_23 bl[23] br[23] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_24 bl[24] br[24] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_25 bl[25] br[25] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_26 bl[26] br[26] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_27 bl[27] br[27] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_28 bl[28] br[28] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_29 bl[29] br[29] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_30 bl[30] br[30] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_31 bl[31] br[31] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_32 bl[32] br[32] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_33 bl[33] br[33] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_34 bl[34] br[34] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_35 bl[35] br[35] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_36 bl[36] br[36] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_37 bl[37] br[37] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_38 bl[38] br[38] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_39 bl[39] br[39] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_40 bl[40] br[40] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_41 bl[41] br[41] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_42 bl[42] br[42] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_43 bl[43] br[43] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_44 bl[44] br[44] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_45 bl[45] br[45] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_46 bl[46] br[46] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_47 bl[47] br[47] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_48 bl[48] br[48] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_49 bl[49] br[49] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_50 bl[50] br[50] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_51 bl[51] br[51] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_52 bl[52] br[52] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_53 bl[53] br[53] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_54 bl[54] br[54] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_55 bl[55] br[55] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_56 bl[56] br[56] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_57 bl[57] br[57] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_58 bl[58] br[58] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_59 bl[59] br[59] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_60 bl[60] br[60] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_61 bl[61] br[61] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_62 bl[62] br[62] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_63 bl[63] br[63] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_64 bl[64] br[64] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_65 bl[65] br[65] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_66 bl[66] br[66] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_67 bl[67] br[67] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_68 bl[68] br[68] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_69 bl[69] br[69] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_70 bl[70] br[70] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_71 bl[71] br[71] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_72 bl[72] br[72] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_73 bl[73] br[73] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_74 bl[74] br[74] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_75 bl[75] br[75] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_76 bl[76] br[76] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_77 bl[77] br[77] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_78 bl[78] br[78] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_79 bl[79] br[79] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_80 bl[80] br[80] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_81 bl[81] br[81] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_82 bl[82] br[82] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_83 bl[83] br[83] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_84 bl[84] br[84] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_85 bl[85] br[85] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_86 bl[86] br[86] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_87 bl[87] br[87] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_88 bl[88] br[88] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_89 bl[89] br[89] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_90 bl[90] br[90] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_91 bl[91] br[91] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_92 bl[92] br[92] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_93 bl[93] br[93] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_94 bl[94] br[94] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_95 bl[95] br[95] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_96 bl[96] br[96] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_97 bl[97] br[97] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_98 bl[98] br[98] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_99 bl[99] br[99] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_100 bl[100] br[100] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_101 bl[101] br[101] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_102 bl[102] br[102] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_103 bl[103] br[103] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_104 bl[104] br[104] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_105 bl[105] br[105] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_106 bl[106] br[106] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_107 bl[107] br[107] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_108 bl[108] br[108] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_109 bl[109] br[109] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_110 bl[110] br[110] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_111 bl[111] br[111] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_112 bl[112] br[112] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_113 bl[113] br[113] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_114 bl[114] br[114] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_115 bl[115] br[115] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_116 bl[116] br[116] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_117 bl[117] br[117] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_118 bl[118] br[118] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_119 bl[119] br[119] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_120 bl[120] br[120] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_121 bl[121] br[121] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_122 bl[122] br[122] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_123 bl[123] br[123] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_124 bl[124] br[124] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_125 bl[125] br[125] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_126 bl[126] br[126] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_127 bl[127] br[127] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_128 bl[128] br[128] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_129 bl[129] br[129] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_130 bl[130] br[130] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_131 bl[131] br[131] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_132 bl[132] br[132] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_133 bl[133] br[133] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_134 bl[134] br[134] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_135 bl[135] br[135] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_136 bl[136] br[136] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_137 bl[137] br[137] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_138 bl[138] br[138] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_139 bl[139] br[139] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_140 bl[140] br[140] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_141 bl[141] br[141] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_142 bl[142] br[142] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_143 bl[143] br[143] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_144 bl[144] br[144] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_145 bl[145] br[145] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_146 bl[146] br[146] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_147 bl[147] br[147] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_148 bl[148] br[148] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_149 bl[149] br[149] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_150 bl[150] br[150] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_151 bl[151] br[151] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_152 bl[152] br[152] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_153 bl[153] br[153] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_154 bl[154] br[154] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_155 bl[155] br[155] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_156 bl[156] br[156] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_157 bl[157] br[157] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_158 bl[158] br[158] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_159 bl[159] br[159] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_160 bl[160] br[160] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_161 bl[161] br[161] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_162 bl[162] br[162] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_163 bl[163] br[163] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_164 bl[164] br[164] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_165 bl[165] br[165] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_166 bl[166] br[166] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_167 bl[167] br[167] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_168 bl[168] br[168] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_169 bl[169] br[169] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_170 bl[170] br[170] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_171 bl[171] br[171] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_172 bl[172] br[172] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_173 bl[173] br[173] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_174 bl[174] br[174] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_175 bl[175] br[175] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_176 bl[176] br[176] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_177 bl[177] br[177] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_178 bl[178] br[178] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_179 bl[179] br[179] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_180 bl[180] br[180] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_181 bl[181] br[181] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_182 bl[182] br[182] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_183 bl[183] br[183] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_184 bl[184] br[184] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_185 bl[185] br[185] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_186 bl[186] br[186] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_187 bl[187] br[187] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_188 bl[188] br[188] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_189 bl[189] br[189] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_190 bl[190] br[190] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_191 bl[191] br[191] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_192 bl[192] br[192] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_193 bl[193] br[193] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_194 bl[194] br[194] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_195 bl[195] br[195] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_196 bl[196] br[196] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_197 bl[197] br[197] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_198 bl[198] br[198] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_199 bl[199] br[199] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_200 bl[200] br[200] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_201 bl[201] br[201] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_202 bl[202] br[202] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_203 bl[203] br[203] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_204 bl[204] br[204] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_205 bl[205] br[205] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_206 bl[206] br[206] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_207 bl[207] br[207] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_208 bl[208] br[208] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_209 bl[209] br[209] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_210 bl[210] br[210] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_211 bl[211] br[211] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_212 bl[212] br[212] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_213 bl[213] br[213] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_214 bl[214] br[214] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_215 bl[215] br[215] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_216 bl[216] br[216] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_217 bl[217] br[217] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_218 bl[218] br[218] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_219 bl[219] br[219] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_220 bl[220] br[220] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_221 bl[221] br[221] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_222 bl[222] br[222] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_223 bl[223] br[223] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_224 bl[224] br[224] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_225 bl[225] br[225] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_226 bl[226] br[226] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_227 bl[227] br[227] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_228 bl[228] br[228] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_229 bl[229] br[229] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_230 bl[230] br[230] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_231 bl[231] br[231] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_232 bl[232] br[232] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_233 bl[233] br[233] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_234 bl[234] br[234] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_235 bl[235] br[235] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_236 bl[236] br[236] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_237 bl[237] br[237] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_238 bl[238] br[238] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_239 bl[239] br[239] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_240 bl[240] br[240] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_241 bl[241] br[241] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_242 bl[242] br[242] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_243 bl[243] br[243] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_244 bl[244] br[244] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_245 bl[245] br[245] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_246 bl[246] br[246] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_247 bl[247] br[247] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_248 bl[248] br[248] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_249 bl[249] br[249] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_250 bl[250] br[250] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_251 bl[251] br[251] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_252 bl[252] br[252] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_253 bl[253] br[253] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_254 bl[254] br[254] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_255 bl[255] br[255] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_256 bl[256] br[256] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_257 bl[257] br[257] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_258 bl[258] br[258] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_259 bl[259] br[259] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_260 bl[260] br[260] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_261 bl[261] br[261] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_262 bl[262] br[262] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_263 bl[263] br[263] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_264 bl[264] br[264] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_265 bl[265] br[265] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_266 bl[266] br[266] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_267 bl[267] br[267] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_268 bl[268] br[268] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_269 bl[269] br[269] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_270 bl[270] br[270] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_271 bl[271] br[271] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_272 bl[272] br[272] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_273 bl[273] br[273] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_274 bl[274] br[274] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_275 bl[275] br[275] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_276 bl[276] br[276] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_277 bl[277] br[277] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_278 bl[278] br[278] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_279 bl[279] br[279] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_280 bl[280] br[280] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_281 bl[281] br[281] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_282 bl[282] br[282] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_283 bl[283] br[283] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_284 bl[284] br[284] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_285 bl[285] br[285] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_286 bl[286] br[286] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_287 bl[287] br[287] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_288 bl[288] br[288] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_289 bl[289] br[289] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_290 bl[290] br[290] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_291 bl[291] br[291] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_292 bl[292] br[292] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_293 bl[293] br[293] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_294 bl[294] br[294] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_295 bl[295] br[295] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_296 bl[296] br[296] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_297 bl[297] br[297] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_298 bl[298] br[298] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_299 bl[299] br[299] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_300 bl[300] br[300] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_301 bl[301] br[301] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_302 bl[302] br[302] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_303 bl[303] br[303] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_304 bl[304] br[304] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_305 bl[305] br[305] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_306 bl[306] br[306] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_307 bl[307] br[307] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_308 bl[308] br[308] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_309 bl[309] br[309] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_310 bl[310] br[310] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_311 bl[311] br[311] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_312 bl[312] br[312] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_313 bl[313] br[313] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_314 bl[314] br[314] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_315 bl[315] br[315] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_316 bl[316] br[316] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_317 bl[317] br[317] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_318 bl[318] br[318] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_319 bl[319] br[319] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_320 bl[320] br[320] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_321 bl[321] br[321] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_322 bl[322] br[322] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_323 bl[323] br[323] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_324 bl[324] br[324] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_325 bl[325] br[325] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_326 bl[326] br[326] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_327 bl[327] br[327] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_328 bl[328] br[328] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_329 bl[329] br[329] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_330 bl[330] br[330] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_331 bl[331] br[331] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_332 bl[332] br[332] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_333 bl[333] br[333] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_334 bl[334] br[334] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_335 bl[335] br[335] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_336 bl[336] br[336] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_337 bl[337] br[337] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_338 bl[338] br[338] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_339 bl[339] br[339] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_340 bl[340] br[340] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_341 bl[341] br[341] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_342 bl[342] br[342] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_343 bl[343] br[343] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_344 bl[344] br[344] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_345 bl[345] br[345] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_346 bl[346] br[346] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_347 bl[347] br[347] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_348 bl[348] br[348] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_349 bl[349] br[349] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_350 bl[350] br[350] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_351 bl[351] br[351] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_352 bl[352] br[352] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_353 bl[353] br[353] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_354 bl[354] br[354] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_355 bl[355] br[355] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_356 bl[356] br[356] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_357 bl[357] br[357] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_358 bl[358] br[358] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_359 bl[359] br[359] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_360 bl[360] br[360] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_361 bl[361] br[361] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_362 bl[362] br[362] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_363 bl[363] br[363] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_364 bl[364] br[364] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_365 bl[365] br[365] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_366 bl[366] br[366] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_367 bl[367] br[367] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_368 bl[368] br[368] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_369 bl[369] br[369] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_370 bl[370] br[370] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_371 bl[371] br[371] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_372 bl[372] br[372] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_373 bl[373] br[373] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_374 bl[374] br[374] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_375 bl[375] br[375] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_376 bl[376] br[376] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_377 bl[377] br[377] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_378 bl[378] br[378] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_379 bl[379] br[379] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_380 bl[380] br[380] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_381 bl[381] br[381] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_382 bl[382] br[382] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_383 bl[383] br[383] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_384 bl[384] br[384] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_385 bl[385] br[385] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_386 bl[386] br[386] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_387 bl[387] br[387] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_388 bl[388] br[388] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_389 bl[389] br[389] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_390 bl[390] br[390] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_391 bl[391] br[391] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_392 bl[392] br[392] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_393 bl[393] br[393] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_394 bl[394] br[394] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_395 bl[395] br[395] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_396 bl[396] br[396] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_397 bl[397] br[397] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_398 bl[398] br[398] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_399 bl[399] br[399] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_400 bl[400] br[400] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_401 bl[401] br[401] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_402 bl[402] br[402] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_403 bl[403] br[403] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_404 bl[404] br[404] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_405 bl[405] br[405] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_406 bl[406] br[406] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_407 bl[407] br[407] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_408 bl[408] br[408] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_409 bl[409] br[409] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_410 bl[410] br[410] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_411 bl[411] br[411] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_412 bl[412] br[412] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_413 bl[413] br[413] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_414 bl[414] br[414] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_415 bl[415] br[415] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_416 bl[416] br[416] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_417 bl[417] br[417] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_418 bl[418] br[418] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_419 bl[419] br[419] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_420 bl[420] br[420] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_421 bl[421] br[421] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_422 bl[422] br[422] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_423 bl[423] br[423] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_424 bl[424] br[424] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_425 bl[425] br[425] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_426 bl[426] br[426] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_427 bl[427] br[427] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_428 bl[428] br[428] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_429 bl[429] br[429] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_430 bl[430] br[430] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_431 bl[431] br[431] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_432 bl[432] br[432] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_433 bl[433] br[433] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_434 bl[434] br[434] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_435 bl[435] br[435] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_436 bl[436] br[436] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_437 bl[437] br[437] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_438 bl[438] br[438] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_439 bl[439] br[439] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_440 bl[440] br[440] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_441 bl[441] br[441] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_442 bl[442] br[442] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_443 bl[443] br[443] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_444 bl[444] br[444] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_445 bl[445] br[445] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_446 bl[446] br[446] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_447 bl[447] br[447] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_448 bl[448] br[448] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_449 bl[449] br[449] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_450 bl[450] br[450] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_451 bl[451] br[451] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_452 bl[452] br[452] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_453 bl[453] br[453] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_454 bl[454] br[454] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_455 bl[455] br[455] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_456 bl[456] br[456] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_457 bl[457] br[457] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_458 bl[458] br[458] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_459 bl[459] br[459] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_460 bl[460] br[460] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_461 bl[461] br[461] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_462 bl[462] br[462] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_463 bl[463] br[463] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_464 bl[464] br[464] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_465 bl[465] br[465] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_466 bl[466] br[466] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_467 bl[467] br[467] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_468 bl[468] br[468] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_469 bl[469] br[469] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_470 bl[470] br[470] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_471 bl[471] br[471] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_472 bl[472] br[472] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_473 bl[473] br[473] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_474 bl[474] br[474] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_475 bl[475] br[475] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_476 bl[476] br[476] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_477 bl[477] br[477] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_478 bl[478] br[478] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_479 bl[479] br[479] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_480 bl[480] br[480] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_481 bl[481] br[481] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_482 bl[482] br[482] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_483 bl[483] br[483] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_484 bl[484] br[484] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_485 bl[485] br[485] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_486 bl[486] br[486] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_487 bl[487] br[487] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_488 bl[488] br[488] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_489 bl[489] br[489] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_490 bl[490] br[490] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_491 bl[491] br[491] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_492 bl[492] br[492] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_493 bl[493] br[493] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_494 bl[494] br[494] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_495 bl[495] br[495] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_496 bl[496] br[496] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_497 bl[497] br[497] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_498 bl[498] br[498] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_499 bl[499] br[499] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_500 bl[500] br[500] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_501 bl[501] br[501] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_502 bl[502] br[502] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_503 bl[503] br[503] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_504 bl[504] br[504] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_505 bl[505] br[505] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_506 bl[506] br[506] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_507 bl[507] br[507] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_508 bl[508] br[508] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_509 bl[509] br[509] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_510 bl[510] br[510] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_29_511 bl[511] br[511] vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xcell_30_0 bl[0] br[0] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_1 bl[1] br[1] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_2 bl[2] br[2] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_3 bl[3] br[3] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_4 bl[4] br[4] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_5 bl[5] br[5] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_6 bl[6] br[6] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_7 bl[7] br[7] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_8 bl[8] br[8] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_9 bl[9] br[9] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_10 bl[10] br[10] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_11 bl[11] br[11] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_12 bl[12] br[12] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_13 bl[13] br[13] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_14 bl[14] br[14] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_15 bl[15] br[15] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_16 bl[16] br[16] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_17 bl[17] br[17] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_18 bl[18] br[18] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_19 bl[19] br[19] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_20 bl[20] br[20] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_21 bl[21] br[21] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_22 bl[22] br[22] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_23 bl[23] br[23] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_24 bl[24] br[24] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_25 bl[25] br[25] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_26 bl[26] br[26] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_27 bl[27] br[27] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_28 bl[28] br[28] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_29 bl[29] br[29] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_30 bl[30] br[30] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_31 bl[31] br[31] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_32 bl[32] br[32] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_33 bl[33] br[33] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_34 bl[34] br[34] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_35 bl[35] br[35] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_36 bl[36] br[36] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_37 bl[37] br[37] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_38 bl[38] br[38] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_39 bl[39] br[39] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_40 bl[40] br[40] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_41 bl[41] br[41] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_42 bl[42] br[42] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_43 bl[43] br[43] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_44 bl[44] br[44] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_45 bl[45] br[45] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_46 bl[46] br[46] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_47 bl[47] br[47] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_48 bl[48] br[48] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_49 bl[49] br[49] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_50 bl[50] br[50] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_51 bl[51] br[51] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_52 bl[52] br[52] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_53 bl[53] br[53] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_54 bl[54] br[54] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_55 bl[55] br[55] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_56 bl[56] br[56] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_57 bl[57] br[57] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_58 bl[58] br[58] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_59 bl[59] br[59] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_60 bl[60] br[60] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_61 bl[61] br[61] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_62 bl[62] br[62] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_63 bl[63] br[63] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_64 bl[64] br[64] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_65 bl[65] br[65] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_66 bl[66] br[66] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_67 bl[67] br[67] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_68 bl[68] br[68] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_69 bl[69] br[69] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_70 bl[70] br[70] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_71 bl[71] br[71] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_72 bl[72] br[72] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_73 bl[73] br[73] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_74 bl[74] br[74] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_75 bl[75] br[75] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_76 bl[76] br[76] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_77 bl[77] br[77] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_78 bl[78] br[78] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_79 bl[79] br[79] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_80 bl[80] br[80] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_81 bl[81] br[81] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_82 bl[82] br[82] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_83 bl[83] br[83] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_84 bl[84] br[84] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_85 bl[85] br[85] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_86 bl[86] br[86] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_87 bl[87] br[87] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_88 bl[88] br[88] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_89 bl[89] br[89] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_90 bl[90] br[90] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_91 bl[91] br[91] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_92 bl[92] br[92] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_93 bl[93] br[93] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_94 bl[94] br[94] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_95 bl[95] br[95] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_96 bl[96] br[96] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_97 bl[97] br[97] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_98 bl[98] br[98] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_99 bl[99] br[99] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_100 bl[100] br[100] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_101 bl[101] br[101] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_102 bl[102] br[102] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_103 bl[103] br[103] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_104 bl[104] br[104] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_105 bl[105] br[105] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_106 bl[106] br[106] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_107 bl[107] br[107] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_108 bl[108] br[108] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_109 bl[109] br[109] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_110 bl[110] br[110] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_111 bl[111] br[111] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_112 bl[112] br[112] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_113 bl[113] br[113] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_114 bl[114] br[114] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_115 bl[115] br[115] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_116 bl[116] br[116] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_117 bl[117] br[117] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_118 bl[118] br[118] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_119 bl[119] br[119] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_120 bl[120] br[120] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_121 bl[121] br[121] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_122 bl[122] br[122] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_123 bl[123] br[123] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_124 bl[124] br[124] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_125 bl[125] br[125] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_126 bl[126] br[126] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_127 bl[127] br[127] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_128 bl[128] br[128] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_129 bl[129] br[129] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_130 bl[130] br[130] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_131 bl[131] br[131] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_132 bl[132] br[132] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_133 bl[133] br[133] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_134 bl[134] br[134] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_135 bl[135] br[135] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_136 bl[136] br[136] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_137 bl[137] br[137] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_138 bl[138] br[138] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_139 bl[139] br[139] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_140 bl[140] br[140] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_141 bl[141] br[141] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_142 bl[142] br[142] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_143 bl[143] br[143] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_144 bl[144] br[144] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_145 bl[145] br[145] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_146 bl[146] br[146] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_147 bl[147] br[147] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_148 bl[148] br[148] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_149 bl[149] br[149] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_150 bl[150] br[150] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_151 bl[151] br[151] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_152 bl[152] br[152] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_153 bl[153] br[153] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_154 bl[154] br[154] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_155 bl[155] br[155] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_156 bl[156] br[156] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_157 bl[157] br[157] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_158 bl[158] br[158] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_159 bl[159] br[159] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_160 bl[160] br[160] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_161 bl[161] br[161] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_162 bl[162] br[162] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_163 bl[163] br[163] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_164 bl[164] br[164] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_165 bl[165] br[165] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_166 bl[166] br[166] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_167 bl[167] br[167] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_168 bl[168] br[168] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_169 bl[169] br[169] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_170 bl[170] br[170] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_171 bl[171] br[171] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_172 bl[172] br[172] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_173 bl[173] br[173] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_174 bl[174] br[174] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_175 bl[175] br[175] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_176 bl[176] br[176] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_177 bl[177] br[177] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_178 bl[178] br[178] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_179 bl[179] br[179] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_180 bl[180] br[180] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_181 bl[181] br[181] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_182 bl[182] br[182] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_183 bl[183] br[183] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_184 bl[184] br[184] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_185 bl[185] br[185] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_186 bl[186] br[186] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_187 bl[187] br[187] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_188 bl[188] br[188] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_189 bl[189] br[189] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_190 bl[190] br[190] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_191 bl[191] br[191] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_192 bl[192] br[192] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_193 bl[193] br[193] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_194 bl[194] br[194] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_195 bl[195] br[195] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_196 bl[196] br[196] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_197 bl[197] br[197] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_198 bl[198] br[198] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_199 bl[199] br[199] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_200 bl[200] br[200] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_201 bl[201] br[201] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_202 bl[202] br[202] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_203 bl[203] br[203] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_204 bl[204] br[204] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_205 bl[205] br[205] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_206 bl[206] br[206] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_207 bl[207] br[207] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_208 bl[208] br[208] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_209 bl[209] br[209] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_210 bl[210] br[210] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_211 bl[211] br[211] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_212 bl[212] br[212] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_213 bl[213] br[213] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_214 bl[214] br[214] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_215 bl[215] br[215] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_216 bl[216] br[216] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_217 bl[217] br[217] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_218 bl[218] br[218] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_219 bl[219] br[219] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_220 bl[220] br[220] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_221 bl[221] br[221] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_222 bl[222] br[222] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_223 bl[223] br[223] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_224 bl[224] br[224] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_225 bl[225] br[225] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_226 bl[226] br[226] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_227 bl[227] br[227] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_228 bl[228] br[228] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_229 bl[229] br[229] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_230 bl[230] br[230] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_231 bl[231] br[231] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_232 bl[232] br[232] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_233 bl[233] br[233] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_234 bl[234] br[234] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_235 bl[235] br[235] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_236 bl[236] br[236] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_237 bl[237] br[237] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_238 bl[238] br[238] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_239 bl[239] br[239] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_240 bl[240] br[240] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_241 bl[241] br[241] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_242 bl[242] br[242] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_243 bl[243] br[243] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_244 bl[244] br[244] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_245 bl[245] br[245] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_246 bl[246] br[246] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_247 bl[247] br[247] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_248 bl[248] br[248] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_249 bl[249] br[249] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_250 bl[250] br[250] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_251 bl[251] br[251] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_252 bl[252] br[252] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_253 bl[253] br[253] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_254 bl[254] br[254] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_255 bl[255] br[255] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_256 bl[256] br[256] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_257 bl[257] br[257] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_258 bl[258] br[258] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_259 bl[259] br[259] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_260 bl[260] br[260] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_261 bl[261] br[261] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_262 bl[262] br[262] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_263 bl[263] br[263] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_264 bl[264] br[264] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_265 bl[265] br[265] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_266 bl[266] br[266] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_267 bl[267] br[267] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_268 bl[268] br[268] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_269 bl[269] br[269] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_270 bl[270] br[270] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_271 bl[271] br[271] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_272 bl[272] br[272] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_273 bl[273] br[273] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_274 bl[274] br[274] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_275 bl[275] br[275] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_276 bl[276] br[276] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_277 bl[277] br[277] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_278 bl[278] br[278] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_279 bl[279] br[279] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_280 bl[280] br[280] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_281 bl[281] br[281] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_282 bl[282] br[282] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_283 bl[283] br[283] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_284 bl[284] br[284] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_285 bl[285] br[285] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_286 bl[286] br[286] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_287 bl[287] br[287] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_288 bl[288] br[288] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_289 bl[289] br[289] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_290 bl[290] br[290] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_291 bl[291] br[291] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_292 bl[292] br[292] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_293 bl[293] br[293] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_294 bl[294] br[294] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_295 bl[295] br[295] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_296 bl[296] br[296] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_297 bl[297] br[297] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_298 bl[298] br[298] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_299 bl[299] br[299] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_300 bl[300] br[300] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_301 bl[301] br[301] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_302 bl[302] br[302] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_303 bl[303] br[303] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_304 bl[304] br[304] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_305 bl[305] br[305] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_306 bl[306] br[306] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_307 bl[307] br[307] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_308 bl[308] br[308] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_309 bl[309] br[309] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_310 bl[310] br[310] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_311 bl[311] br[311] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_312 bl[312] br[312] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_313 bl[313] br[313] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_314 bl[314] br[314] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_315 bl[315] br[315] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_316 bl[316] br[316] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_317 bl[317] br[317] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_318 bl[318] br[318] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_319 bl[319] br[319] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_320 bl[320] br[320] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_321 bl[321] br[321] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_322 bl[322] br[322] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_323 bl[323] br[323] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_324 bl[324] br[324] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_325 bl[325] br[325] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_326 bl[326] br[326] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_327 bl[327] br[327] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_328 bl[328] br[328] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_329 bl[329] br[329] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_330 bl[330] br[330] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_331 bl[331] br[331] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_332 bl[332] br[332] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_333 bl[333] br[333] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_334 bl[334] br[334] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_335 bl[335] br[335] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_336 bl[336] br[336] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_337 bl[337] br[337] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_338 bl[338] br[338] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_339 bl[339] br[339] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_340 bl[340] br[340] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_341 bl[341] br[341] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_342 bl[342] br[342] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_343 bl[343] br[343] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_344 bl[344] br[344] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_345 bl[345] br[345] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_346 bl[346] br[346] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_347 bl[347] br[347] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_348 bl[348] br[348] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_349 bl[349] br[349] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_350 bl[350] br[350] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_351 bl[351] br[351] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_352 bl[352] br[352] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_353 bl[353] br[353] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_354 bl[354] br[354] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_355 bl[355] br[355] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_356 bl[356] br[356] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_357 bl[357] br[357] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_358 bl[358] br[358] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_359 bl[359] br[359] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_360 bl[360] br[360] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_361 bl[361] br[361] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_362 bl[362] br[362] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_363 bl[363] br[363] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_364 bl[364] br[364] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_365 bl[365] br[365] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_366 bl[366] br[366] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_367 bl[367] br[367] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_368 bl[368] br[368] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_369 bl[369] br[369] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_370 bl[370] br[370] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_371 bl[371] br[371] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_372 bl[372] br[372] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_373 bl[373] br[373] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_374 bl[374] br[374] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_375 bl[375] br[375] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_376 bl[376] br[376] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_377 bl[377] br[377] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_378 bl[378] br[378] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_379 bl[379] br[379] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_380 bl[380] br[380] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_381 bl[381] br[381] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_382 bl[382] br[382] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_383 bl[383] br[383] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_384 bl[384] br[384] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_385 bl[385] br[385] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_386 bl[386] br[386] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_387 bl[387] br[387] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_388 bl[388] br[388] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_389 bl[389] br[389] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_390 bl[390] br[390] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_391 bl[391] br[391] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_392 bl[392] br[392] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_393 bl[393] br[393] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_394 bl[394] br[394] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_395 bl[395] br[395] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_396 bl[396] br[396] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_397 bl[397] br[397] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_398 bl[398] br[398] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_399 bl[399] br[399] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_400 bl[400] br[400] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_401 bl[401] br[401] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_402 bl[402] br[402] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_403 bl[403] br[403] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_404 bl[404] br[404] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_405 bl[405] br[405] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_406 bl[406] br[406] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_407 bl[407] br[407] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_408 bl[408] br[408] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_409 bl[409] br[409] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_410 bl[410] br[410] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_411 bl[411] br[411] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_412 bl[412] br[412] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_413 bl[413] br[413] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_414 bl[414] br[414] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_415 bl[415] br[415] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_416 bl[416] br[416] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_417 bl[417] br[417] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_418 bl[418] br[418] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_419 bl[419] br[419] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_420 bl[420] br[420] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_421 bl[421] br[421] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_422 bl[422] br[422] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_423 bl[423] br[423] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_424 bl[424] br[424] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_425 bl[425] br[425] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_426 bl[426] br[426] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_427 bl[427] br[427] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_428 bl[428] br[428] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_429 bl[429] br[429] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_430 bl[430] br[430] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_431 bl[431] br[431] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_432 bl[432] br[432] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_433 bl[433] br[433] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_434 bl[434] br[434] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_435 bl[435] br[435] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_436 bl[436] br[436] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_437 bl[437] br[437] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_438 bl[438] br[438] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_439 bl[439] br[439] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_440 bl[440] br[440] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_441 bl[441] br[441] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_442 bl[442] br[442] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_443 bl[443] br[443] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_444 bl[444] br[444] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_445 bl[445] br[445] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_446 bl[446] br[446] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_447 bl[447] br[447] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_448 bl[448] br[448] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_449 bl[449] br[449] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_450 bl[450] br[450] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_451 bl[451] br[451] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_452 bl[452] br[452] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_453 bl[453] br[453] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_454 bl[454] br[454] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_455 bl[455] br[455] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_456 bl[456] br[456] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_457 bl[457] br[457] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_458 bl[458] br[458] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_459 bl[459] br[459] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_460 bl[460] br[460] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_461 bl[461] br[461] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_462 bl[462] br[462] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_463 bl[463] br[463] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_464 bl[464] br[464] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_465 bl[465] br[465] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_466 bl[466] br[466] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_467 bl[467] br[467] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_468 bl[468] br[468] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_469 bl[469] br[469] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_470 bl[470] br[470] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_471 bl[471] br[471] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_472 bl[472] br[472] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_473 bl[473] br[473] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_474 bl[474] br[474] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_475 bl[475] br[475] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_476 bl[476] br[476] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_477 bl[477] br[477] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_478 bl[478] br[478] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_479 bl[479] br[479] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_480 bl[480] br[480] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_481 bl[481] br[481] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_482 bl[482] br[482] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_483 bl[483] br[483] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_484 bl[484] br[484] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_485 bl[485] br[485] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_486 bl[486] br[486] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_487 bl[487] br[487] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_488 bl[488] br[488] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_489 bl[489] br[489] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_490 bl[490] br[490] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_491 bl[491] br[491] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_492 bl[492] br[492] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_493 bl[493] br[493] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_494 bl[494] br[494] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_495 bl[495] br[495] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_496 bl[496] br[496] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_497 bl[497] br[497] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_498 bl[498] br[498] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_499 bl[499] br[499] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_500 bl[500] br[500] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_501 bl[501] br[501] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_502 bl[502] br[502] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_503 bl[503] br[503] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_504 bl[504] br[504] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_505 bl[505] br[505] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_506 bl[506] br[506] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_507 bl[507] br[507] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_508 bl[508] br[508] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_509 bl[509] br[509] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_510 bl[510] br[510] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_30_511 bl[511] br[511] vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xcell_31_0 bl[0] br[0] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_1 bl[1] br[1] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_2 bl[2] br[2] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_3 bl[3] br[3] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_4 bl[4] br[4] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_5 bl[5] br[5] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_6 bl[6] br[6] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_7 bl[7] br[7] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_8 bl[8] br[8] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_9 bl[9] br[9] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_10 bl[10] br[10] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_11 bl[11] br[11] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_12 bl[12] br[12] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_13 bl[13] br[13] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_14 bl[14] br[14] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_15 bl[15] br[15] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_16 bl[16] br[16] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_17 bl[17] br[17] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_18 bl[18] br[18] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_19 bl[19] br[19] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_20 bl[20] br[20] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_21 bl[21] br[21] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_22 bl[22] br[22] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_23 bl[23] br[23] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_24 bl[24] br[24] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_25 bl[25] br[25] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_26 bl[26] br[26] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_27 bl[27] br[27] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_28 bl[28] br[28] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_29 bl[29] br[29] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_30 bl[30] br[30] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_31 bl[31] br[31] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_32 bl[32] br[32] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_33 bl[33] br[33] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_34 bl[34] br[34] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_35 bl[35] br[35] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_36 bl[36] br[36] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_37 bl[37] br[37] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_38 bl[38] br[38] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_39 bl[39] br[39] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_40 bl[40] br[40] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_41 bl[41] br[41] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_42 bl[42] br[42] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_43 bl[43] br[43] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_44 bl[44] br[44] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_45 bl[45] br[45] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_46 bl[46] br[46] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_47 bl[47] br[47] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_48 bl[48] br[48] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_49 bl[49] br[49] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_50 bl[50] br[50] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_51 bl[51] br[51] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_52 bl[52] br[52] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_53 bl[53] br[53] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_54 bl[54] br[54] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_55 bl[55] br[55] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_56 bl[56] br[56] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_57 bl[57] br[57] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_58 bl[58] br[58] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_59 bl[59] br[59] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_60 bl[60] br[60] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_61 bl[61] br[61] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_62 bl[62] br[62] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_63 bl[63] br[63] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_64 bl[64] br[64] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_65 bl[65] br[65] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_66 bl[66] br[66] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_67 bl[67] br[67] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_68 bl[68] br[68] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_69 bl[69] br[69] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_70 bl[70] br[70] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_71 bl[71] br[71] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_72 bl[72] br[72] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_73 bl[73] br[73] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_74 bl[74] br[74] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_75 bl[75] br[75] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_76 bl[76] br[76] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_77 bl[77] br[77] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_78 bl[78] br[78] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_79 bl[79] br[79] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_80 bl[80] br[80] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_81 bl[81] br[81] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_82 bl[82] br[82] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_83 bl[83] br[83] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_84 bl[84] br[84] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_85 bl[85] br[85] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_86 bl[86] br[86] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_87 bl[87] br[87] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_88 bl[88] br[88] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_89 bl[89] br[89] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_90 bl[90] br[90] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_91 bl[91] br[91] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_92 bl[92] br[92] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_93 bl[93] br[93] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_94 bl[94] br[94] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_95 bl[95] br[95] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_96 bl[96] br[96] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_97 bl[97] br[97] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_98 bl[98] br[98] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_99 bl[99] br[99] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_100 bl[100] br[100] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_101 bl[101] br[101] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_102 bl[102] br[102] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_103 bl[103] br[103] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_104 bl[104] br[104] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_105 bl[105] br[105] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_106 bl[106] br[106] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_107 bl[107] br[107] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_108 bl[108] br[108] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_109 bl[109] br[109] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_110 bl[110] br[110] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_111 bl[111] br[111] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_112 bl[112] br[112] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_113 bl[113] br[113] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_114 bl[114] br[114] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_115 bl[115] br[115] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_116 bl[116] br[116] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_117 bl[117] br[117] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_118 bl[118] br[118] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_119 bl[119] br[119] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_120 bl[120] br[120] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_121 bl[121] br[121] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_122 bl[122] br[122] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_123 bl[123] br[123] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_124 bl[124] br[124] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_125 bl[125] br[125] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_126 bl[126] br[126] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_127 bl[127] br[127] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_128 bl[128] br[128] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_129 bl[129] br[129] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_130 bl[130] br[130] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_131 bl[131] br[131] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_132 bl[132] br[132] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_133 bl[133] br[133] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_134 bl[134] br[134] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_135 bl[135] br[135] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_136 bl[136] br[136] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_137 bl[137] br[137] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_138 bl[138] br[138] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_139 bl[139] br[139] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_140 bl[140] br[140] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_141 bl[141] br[141] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_142 bl[142] br[142] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_143 bl[143] br[143] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_144 bl[144] br[144] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_145 bl[145] br[145] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_146 bl[146] br[146] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_147 bl[147] br[147] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_148 bl[148] br[148] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_149 bl[149] br[149] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_150 bl[150] br[150] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_151 bl[151] br[151] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_152 bl[152] br[152] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_153 bl[153] br[153] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_154 bl[154] br[154] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_155 bl[155] br[155] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_156 bl[156] br[156] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_157 bl[157] br[157] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_158 bl[158] br[158] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_159 bl[159] br[159] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_160 bl[160] br[160] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_161 bl[161] br[161] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_162 bl[162] br[162] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_163 bl[163] br[163] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_164 bl[164] br[164] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_165 bl[165] br[165] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_166 bl[166] br[166] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_167 bl[167] br[167] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_168 bl[168] br[168] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_169 bl[169] br[169] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_170 bl[170] br[170] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_171 bl[171] br[171] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_172 bl[172] br[172] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_173 bl[173] br[173] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_174 bl[174] br[174] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_175 bl[175] br[175] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_176 bl[176] br[176] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_177 bl[177] br[177] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_178 bl[178] br[178] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_179 bl[179] br[179] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_180 bl[180] br[180] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_181 bl[181] br[181] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_182 bl[182] br[182] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_183 bl[183] br[183] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_184 bl[184] br[184] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_185 bl[185] br[185] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_186 bl[186] br[186] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_187 bl[187] br[187] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_188 bl[188] br[188] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_189 bl[189] br[189] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_190 bl[190] br[190] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_191 bl[191] br[191] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_192 bl[192] br[192] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_193 bl[193] br[193] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_194 bl[194] br[194] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_195 bl[195] br[195] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_196 bl[196] br[196] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_197 bl[197] br[197] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_198 bl[198] br[198] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_199 bl[199] br[199] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_200 bl[200] br[200] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_201 bl[201] br[201] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_202 bl[202] br[202] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_203 bl[203] br[203] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_204 bl[204] br[204] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_205 bl[205] br[205] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_206 bl[206] br[206] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_207 bl[207] br[207] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_208 bl[208] br[208] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_209 bl[209] br[209] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_210 bl[210] br[210] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_211 bl[211] br[211] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_212 bl[212] br[212] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_213 bl[213] br[213] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_214 bl[214] br[214] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_215 bl[215] br[215] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_216 bl[216] br[216] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_217 bl[217] br[217] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_218 bl[218] br[218] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_219 bl[219] br[219] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_220 bl[220] br[220] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_221 bl[221] br[221] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_222 bl[222] br[222] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_223 bl[223] br[223] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_224 bl[224] br[224] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_225 bl[225] br[225] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_226 bl[226] br[226] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_227 bl[227] br[227] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_228 bl[228] br[228] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_229 bl[229] br[229] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_230 bl[230] br[230] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_231 bl[231] br[231] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_232 bl[232] br[232] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_233 bl[233] br[233] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_234 bl[234] br[234] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_235 bl[235] br[235] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_236 bl[236] br[236] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_237 bl[237] br[237] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_238 bl[238] br[238] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_239 bl[239] br[239] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_240 bl[240] br[240] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_241 bl[241] br[241] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_242 bl[242] br[242] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_243 bl[243] br[243] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_244 bl[244] br[244] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_245 bl[245] br[245] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_246 bl[246] br[246] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_247 bl[247] br[247] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_248 bl[248] br[248] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_249 bl[249] br[249] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_250 bl[250] br[250] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_251 bl[251] br[251] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_252 bl[252] br[252] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_253 bl[253] br[253] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_254 bl[254] br[254] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_255 bl[255] br[255] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_256 bl[256] br[256] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_257 bl[257] br[257] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_258 bl[258] br[258] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_259 bl[259] br[259] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_260 bl[260] br[260] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_261 bl[261] br[261] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_262 bl[262] br[262] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_263 bl[263] br[263] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_264 bl[264] br[264] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_265 bl[265] br[265] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_266 bl[266] br[266] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_267 bl[267] br[267] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_268 bl[268] br[268] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_269 bl[269] br[269] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_270 bl[270] br[270] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_271 bl[271] br[271] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_272 bl[272] br[272] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_273 bl[273] br[273] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_274 bl[274] br[274] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_275 bl[275] br[275] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_276 bl[276] br[276] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_277 bl[277] br[277] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_278 bl[278] br[278] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_279 bl[279] br[279] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_280 bl[280] br[280] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_281 bl[281] br[281] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_282 bl[282] br[282] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_283 bl[283] br[283] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_284 bl[284] br[284] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_285 bl[285] br[285] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_286 bl[286] br[286] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_287 bl[287] br[287] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_288 bl[288] br[288] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_289 bl[289] br[289] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_290 bl[290] br[290] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_291 bl[291] br[291] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_292 bl[292] br[292] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_293 bl[293] br[293] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_294 bl[294] br[294] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_295 bl[295] br[295] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_296 bl[296] br[296] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_297 bl[297] br[297] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_298 bl[298] br[298] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_299 bl[299] br[299] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_300 bl[300] br[300] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_301 bl[301] br[301] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_302 bl[302] br[302] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_303 bl[303] br[303] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_304 bl[304] br[304] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_305 bl[305] br[305] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_306 bl[306] br[306] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_307 bl[307] br[307] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_308 bl[308] br[308] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_309 bl[309] br[309] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_310 bl[310] br[310] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_311 bl[311] br[311] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_312 bl[312] br[312] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_313 bl[313] br[313] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_314 bl[314] br[314] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_315 bl[315] br[315] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_316 bl[316] br[316] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_317 bl[317] br[317] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_318 bl[318] br[318] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_319 bl[319] br[319] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_320 bl[320] br[320] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_321 bl[321] br[321] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_322 bl[322] br[322] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_323 bl[323] br[323] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_324 bl[324] br[324] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_325 bl[325] br[325] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_326 bl[326] br[326] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_327 bl[327] br[327] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_328 bl[328] br[328] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_329 bl[329] br[329] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_330 bl[330] br[330] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_331 bl[331] br[331] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_332 bl[332] br[332] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_333 bl[333] br[333] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_334 bl[334] br[334] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_335 bl[335] br[335] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_336 bl[336] br[336] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_337 bl[337] br[337] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_338 bl[338] br[338] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_339 bl[339] br[339] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_340 bl[340] br[340] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_341 bl[341] br[341] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_342 bl[342] br[342] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_343 bl[343] br[343] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_344 bl[344] br[344] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_345 bl[345] br[345] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_346 bl[346] br[346] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_347 bl[347] br[347] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_348 bl[348] br[348] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_349 bl[349] br[349] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_350 bl[350] br[350] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_351 bl[351] br[351] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_352 bl[352] br[352] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_353 bl[353] br[353] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_354 bl[354] br[354] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_355 bl[355] br[355] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_356 bl[356] br[356] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_357 bl[357] br[357] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_358 bl[358] br[358] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_359 bl[359] br[359] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_360 bl[360] br[360] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_361 bl[361] br[361] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_362 bl[362] br[362] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_363 bl[363] br[363] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_364 bl[364] br[364] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_365 bl[365] br[365] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_366 bl[366] br[366] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_367 bl[367] br[367] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_368 bl[368] br[368] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_369 bl[369] br[369] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_370 bl[370] br[370] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_371 bl[371] br[371] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_372 bl[372] br[372] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_373 bl[373] br[373] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_374 bl[374] br[374] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_375 bl[375] br[375] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_376 bl[376] br[376] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_377 bl[377] br[377] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_378 bl[378] br[378] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_379 bl[379] br[379] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_380 bl[380] br[380] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_381 bl[381] br[381] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_382 bl[382] br[382] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_383 bl[383] br[383] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_384 bl[384] br[384] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_385 bl[385] br[385] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_386 bl[386] br[386] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_387 bl[387] br[387] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_388 bl[388] br[388] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_389 bl[389] br[389] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_390 bl[390] br[390] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_391 bl[391] br[391] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_392 bl[392] br[392] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_393 bl[393] br[393] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_394 bl[394] br[394] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_395 bl[395] br[395] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_396 bl[396] br[396] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_397 bl[397] br[397] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_398 bl[398] br[398] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_399 bl[399] br[399] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_400 bl[400] br[400] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_401 bl[401] br[401] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_402 bl[402] br[402] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_403 bl[403] br[403] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_404 bl[404] br[404] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_405 bl[405] br[405] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_406 bl[406] br[406] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_407 bl[407] br[407] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_408 bl[408] br[408] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_409 bl[409] br[409] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_410 bl[410] br[410] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_411 bl[411] br[411] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_412 bl[412] br[412] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_413 bl[413] br[413] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_414 bl[414] br[414] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_415 bl[415] br[415] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_416 bl[416] br[416] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_417 bl[417] br[417] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_418 bl[418] br[418] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_419 bl[419] br[419] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_420 bl[420] br[420] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_421 bl[421] br[421] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_422 bl[422] br[422] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_423 bl[423] br[423] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_424 bl[424] br[424] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_425 bl[425] br[425] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_426 bl[426] br[426] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_427 bl[427] br[427] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_428 bl[428] br[428] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_429 bl[429] br[429] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_430 bl[430] br[430] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_431 bl[431] br[431] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_432 bl[432] br[432] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_433 bl[433] br[433] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_434 bl[434] br[434] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_435 bl[435] br[435] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_436 bl[436] br[436] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_437 bl[437] br[437] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_438 bl[438] br[438] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_439 bl[439] br[439] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_440 bl[440] br[440] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_441 bl[441] br[441] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_442 bl[442] br[442] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_443 bl[443] br[443] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_444 bl[444] br[444] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_445 bl[445] br[445] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_446 bl[446] br[446] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_447 bl[447] br[447] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_448 bl[448] br[448] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_449 bl[449] br[449] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_450 bl[450] br[450] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_451 bl[451] br[451] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_452 bl[452] br[452] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_453 bl[453] br[453] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_454 bl[454] br[454] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_455 bl[455] br[455] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_456 bl[456] br[456] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_457 bl[457] br[457] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_458 bl[458] br[458] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_459 bl[459] br[459] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_460 bl[460] br[460] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_461 bl[461] br[461] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_462 bl[462] br[462] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_463 bl[463] br[463] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_464 bl[464] br[464] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_465 bl[465] br[465] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_466 bl[466] br[466] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_467 bl[467] br[467] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_468 bl[468] br[468] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_469 bl[469] br[469] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_470 bl[470] br[470] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_471 bl[471] br[471] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_472 bl[472] br[472] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_473 bl[473] br[473] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_474 bl[474] br[474] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_475 bl[475] br[475] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_476 bl[476] br[476] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_477 bl[477] br[477] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_478 bl[478] br[478] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_479 bl[479] br[479] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_480 bl[480] br[480] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_481 bl[481] br[481] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_482 bl[482] br[482] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_483 bl[483] br[483] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_484 bl[484] br[484] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_485 bl[485] br[485] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_486 bl[486] br[486] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_487 bl[487] br[487] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_488 bl[488] br[488] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_489 bl[489] br[489] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_490 bl[490] br[490] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_491 bl[491] br[491] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_492 bl[492] br[492] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_493 bl[493] br[493] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_494 bl[494] br[494] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_495 bl[495] br[495] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_496 bl[496] br[496] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_497 bl[497] br[497] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_498 bl[498] br[498] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_499 bl[499] br[499] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_500 bl[500] br[500] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_501 bl[501] br[501] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_502 bl[502] br[502] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_503 bl[503] br[503] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_504 bl[504] br[504] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_505 bl[505] br[505] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_506 bl[506] br[506] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_507 bl[507] br[507] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_508 bl[508] br[508] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_509 bl[509] br[509] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_510 bl[510] br[510] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_31_511 bl[511] br[511] vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xcell_32_0 bl[0] br[0] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_1 bl[1] br[1] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_2 bl[2] br[2] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_3 bl[3] br[3] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_4 bl[4] br[4] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_5 bl[5] br[5] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_6 bl[6] br[6] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_7 bl[7] br[7] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_8 bl[8] br[8] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_9 bl[9] br[9] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_10 bl[10] br[10] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_11 bl[11] br[11] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_12 bl[12] br[12] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_13 bl[13] br[13] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_14 bl[14] br[14] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_15 bl[15] br[15] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_16 bl[16] br[16] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_17 bl[17] br[17] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_18 bl[18] br[18] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_19 bl[19] br[19] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_20 bl[20] br[20] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_21 bl[21] br[21] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_22 bl[22] br[22] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_23 bl[23] br[23] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_24 bl[24] br[24] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_25 bl[25] br[25] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_26 bl[26] br[26] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_27 bl[27] br[27] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_28 bl[28] br[28] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_29 bl[29] br[29] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_30 bl[30] br[30] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_31 bl[31] br[31] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_32 bl[32] br[32] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_33 bl[33] br[33] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_34 bl[34] br[34] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_35 bl[35] br[35] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_36 bl[36] br[36] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_37 bl[37] br[37] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_38 bl[38] br[38] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_39 bl[39] br[39] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_40 bl[40] br[40] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_41 bl[41] br[41] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_42 bl[42] br[42] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_43 bl[43] br[43] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_44 bl[44] br[44] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_45 bl[45] br[45] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_46 bl[46] br[46] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_47 bl[47] br[47] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_48 bl[48] br[48] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_49 bl[49] br[49] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_50 bl[50] br[50] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_51 bl[51] br[51] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_52 bl[52] br[52] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_53 bl[53] br[53] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_54 bl[54] br[54] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_55 bl[55] br[55] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_56 bl[56] br[56] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_57 bl[57] br[57] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_58 bl[58] br[58] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_59 bl[59] br[59] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_60 bl[60] br[60] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_61 bl[61] br[61] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_62 bl[62] br[62] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_63 bl[63] br[63] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_64 bl[64] br[64] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_65 bl[65] br[65] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_66 bl[66] br[66] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_67 bl[67] br[67] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_68 bl[68] br[68] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_69 bl[69] br[69] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_70 bl[70] br[70] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_71 bl[71] br[71] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_72 bl[72] br[72] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_73 bl[73] br[73] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_74 bl[74] br[74] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_75 bl[75] br[75] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_76 bl[76] br[76] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_77 bl[77] br[77] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_78 bl[78] br[78] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_79 bl[79] br[79] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_80 bl[80] br[80] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_81 bl[81] br[81] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_82 bl[82] br[82] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_83 bl[83] br[83] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_84 bl[84] br[84] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_85 bl[85] br[85] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_86 bl[86] br[86] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_87 bl[87] br[87] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_88 bl[88] br[88] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_89 bl[89] br[89] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_90 bl[90] br[90] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_91 bl[91] br[91] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_92 bl[92] br[92] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_93 bl[93] br[93] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_94 bl[94] br[94] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_95 bl[95] br[95] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_96 bl[96] br[96] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_97 bl[97] br[97] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_98 bl[98] br[98] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_99 bl[99] br[99] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_100 bl[100] br[100] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_101 bl[101] br[101] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_102 bl[102] br[102] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_103 bl[103] br[103] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_104 bl[104] br[104] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_105 bl[105] br[105] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_106 bl[106] br[106] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_107 bl[107] br[107] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_108 bl[108] br[108] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_109 bl[109] br[109] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_110 bl[110] br[110] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_111 bl[111] br[111] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_112 bl[112] br[112] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_113 bl[113] br[113] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_114 bl[114] br[114] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_115 bl[115] br[115] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_116 bl[116] br[116] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_117 bl[117] br[117] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_118 bl[118] br[118] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_119 bl[119] br[119] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_120 bl[120] br[120] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_121 bl[121] br[121] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_122 bl[122] br[122] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_123 bl[123] br[123] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_124 bl[124] br[124] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_125 bl[125] br[125] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_126 bl[126] br[126] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_127 bl[127] br[127] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_128 bl[128] br[128] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_129 bl[129] br[129] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_130 bl[130] br[130] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_131 bl[131] br[131] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_132 bl[132] br[132] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_133 bl[133] br[133] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_134 bl[134] br[134] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_135 bl[135] br[135] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_136 bl[136] br[136] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_137 bl[137] br[137] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_138 bl[138] br[138] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_139 bl[139] br[139] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_140 bl[140] br[140] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_141 bl[141] br[141] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_142 bl[142] br[142] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_143 bl[143] br[143] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_144 bl[144] br[144] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_145 bl[145] br[145] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_146 bl[146] br[146] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_147 bl[147] br[147] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_148 bl[148] br[148] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_149 bl[149] br[149] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_150 bl[150] br[150] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_151 bl[151] br[151] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_152 bl[152] br[152] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_153 bl[153] br[153] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_154 bl[154] br[154] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_155 bl[155] br[155] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_156 bl[156] br[156] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_157 bl[157] br[157] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_158 bl[158] br[158] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_159 bl[159] br[159] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_160 bl[160] br[160] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_161 bl[161] br[161] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_162 bl[162] br[162] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_163 bl[163] br[163] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_164 bl[164] br[164] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_165 bl[165] br[165] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_166 bl[166] br[166] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_167 bl[167] br[167] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_168 bl[168] br[168] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_169 bl[169] br[169] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_170 bl[170] br[170] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_171 bl[171] br[171] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_172 bl[172] br[172] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_173 bl[173] br[173] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_174 bl[174] br[174] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_175 bl[175] br[175] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_176 bl[176] br[176] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_177 bl[177] br[177] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_178 bl[178] br[178] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_179 bl[179] br[179] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_180 bl[180] br[180] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_181 bl[181] br[181] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_182 bl[182] br[182] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_183 bl[183] br[183] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_184 bl[184] br[184] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_185 bl[185] br[185] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_186 bl[186] br[186] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_187 bl[187] br[187] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_188 bl[188] br[188] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_189 bl[189] br[189] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_190 bl[190] br[190] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_191 bl[191] br[191] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_192 bl[192] br[192] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_193 bl[193] br[193] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_194 bl[194] br[194] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_195 bl[195] br[195] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_196 bl[196] br[196] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_197 bl[197] br[197] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_198 bl[198] br[198] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_199 bl[199] br[199] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_200 bl[200] br[200] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_201 bl[201] br[201] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_202 bl[202] br[202] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_203 bl[203] br[203] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_204 bl[204] br[204] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_205 bl[205] br[205] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_206 bl[206] br[206] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_207 bl[207] br[207] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_208 bl[208] br[208] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_209 bl[209] br[209] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_210 bl[210] br[210] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_211 bl[211] br[211] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_212 bl[212] br[212] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_213 bl[213] br[213] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_214 bl[214] br[214] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_215 bl[215] br[215] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_216 bl[216] br[216] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_217 bl[217] br[217] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_218 bl[218] br[218] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_219 bl[219] br[219] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_220 bl[220] br[220] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_221 bl[221] br[221] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_222 bl[222] br[222] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_223 bl[223] br[223] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_224 bl[224] br[224] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_225 bl[225] br[225] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_226 bl[226] br[226] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_227 bl[227] br[227] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_228 bl[228] br[228] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_229 bl[229] br[229] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_230 bl[230] br[230] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_231 bl[231] br[231] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_232 bl[232] br[232] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_233 bl[233] br[233] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_234 bl[234] br[234] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_235 bl[235] br[235] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_236 bl[236] br[236] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_237 bl[237] br[237] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_238 bl[238] br[238] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_239 bl[239] br[239] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_240 bl[240] br[240] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_241 bl[241] br[241] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_242 bl[242] br[242] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_243 bl[243] br[243] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_244 bl[244] br[244] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_245 bl[245] br[245] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_246 bl[246] br[246] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_247 bl[247] br[247] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_248 bl[248] br[248] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_249 bl[249] br[249] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_250 bl[250] br[250] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_251 bl[251] br[251] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_252 bl[252] br[252] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_253 bl[253] br[253] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_254 bl[254] br[254] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_255 bl[255] br[255] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_256 bl[256] br[256] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_257 bl[257] br[257] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_258 bl[258] br[258] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_259 bl[259] br[259] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_260 bl[260] br[260] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_261 bl[261] br[261] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_262 bl[262] br[262] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_263 bl[263] br[263] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_264 bl[264] br[264] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_265 bl[265] br[265] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_266 bl[266] br[266] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_267 bl[267] br[267] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_268 bl[268] br[268] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_269 bl[269] br[269] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_270 bl[270] br[270] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_271 bl[271] br[271] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_272 bl[272] br[272] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_273 bl[273] br[273] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_274 bl[274] br[274] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_275 bl[275] br[275] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_276 bl[276] br[276] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_277 bl[277] br[277] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_278 bl[278] br[278] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_279 bl[279] br[279] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_280 bl[280] br[280] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_281 bl[281] br[281] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_282 bl[282] br[282] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_283 bl[283] br[283] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_284 bl[284] br[284] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_285 bl[285] br[285] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_286 bl[286] br[286] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_287 bl[287] br[287] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_288 bl[288] br[288] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_289 bl[289] br[289] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_290 bl[290] br[290] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_291 bl[291] br[291] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_292 bl[292] br[292] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_293 bl[293] br[293] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_294 bl[294] br[294] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_295 bl[295] br[295] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_296 bl[296] br[296] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_297 bl[297] br[297] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_298 bl[298] br[298] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_299 bl[299] br[299] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_300 bl[300] br[300] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_301 bl[301] br[301] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_302 bl[302] br[302] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_303 bl[303] br[303] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_304 bl[304] br[304] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_305 bl[305] br[305] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_306 bl[306] br[306] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_307 bl[307] br[307] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_308 bl[308] br[308] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_309 bl[309] br[309] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_310 bl[310] br[310] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_311 bl[311] br[311] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_312 bl[312] br[312] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_313 bl[313] br[313] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_314 bl[314] br[314] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_315 bl[315] br[315] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_316 bl[316] br[316] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_317 bl[317] br[317] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_318 bl[318] br[318] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_319 bl[319] br[319] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_320 bl[320] br[320] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_321 bl[321] br[321] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_322 bl[322] br[322] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_323 bl[323] br[323] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_324 bl[324] br[324] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_325 bl[325] br[325] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_326 bl[326] br[326] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_327 bl[327] br[327] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_328 bl[328] br[328] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_329 bl[329] br[329] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_330 bl[330] br[330] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_331 bl[331] br[331] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_332 bl[332] br[332] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_333 bl[333] br[333] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_334 bl[334] br[334] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_335 bl[335] br[335] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_336 bl[336] br[336] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_337 bl[337] br[337] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_338 bl[338] br[338] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_339 bl[339] br[339] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_340 bl[340] br[340] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_341 bl[341] br[341] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_342 bl[342] br[342] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_343 bl[343] br[343] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_344 bl[344] br[344] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_345 bl[345] br[345] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_346 bl[346] br[346] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_347 bl[347] br[347] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_348 bl[348] br[348] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_349 bl[349] br[349] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_350 bl[350] br[350] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_351 bl[351] br[351] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_352 bl[352] br[352] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_353 bl[353] br[353] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_354 bl[354] br[354] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_355 bl[355] br[355] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_356 bl[356] br[356] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_357 bl[357] br[357] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_358 bl[358] br[358] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_359 bl[359] br[359] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_360 bl[360] br[360] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_361 bl[361] br[361] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_362 bl[362] br[362] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_363 bl[363] br[363] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_364 bl[364] br[364] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_365 bl[365] br[365] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_366 bl[366] br[366] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_367 bl[367] br[367] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_368 bl[368] br[368] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_369 bl[369] br[369] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_370 bl[370] br[370] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_371 bl[371] br[371] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_372 bl[372] br[372] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_373 bl[373] br[373] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_374 bl[374] br[374] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_375 bl[375] br[375] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_376 bl[376] br[376] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_377 bl[377] br[377] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_378 bl[378] br[378] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_379 bl[379] br[379] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_380 bl[380] br[380] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_381 bl[381] br[381] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_382 bl[382] br[382] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_383 bl[383] br[383] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_384 bl[384] br[384] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_385 bl[385] br[385] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_386 bl[386] br[386] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_387 bl[387] br[387] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_388 bl[388] br[388] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_389 bl[389] br[389] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_390 bl[390] br[390] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_391 bl[391] br[391] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_392 bl[392] br[392] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_393 bl[393] br[393] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_394 bl[394] br[394] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_395 bl[395] br[395] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_396 bl[396] br[396] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_397 bl[397] br[397] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_398 bl[398] br[398] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_399 bl[399] br[399] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_400 bl[400] br[400] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_401 bl[401] br[401] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_402 bl[402] br[402] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_403 bl[403] br[403] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_404 bl[404] br[404] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_405 bl[405] br[405] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_406 bl[406] br[406] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_407 bl[407] br[407] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_408 bl[408] br[408] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_409 bl[409] br[409] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_410 bl[410] br[410] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_411 bl[411] br[411] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_412 bl[412] br[412] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_413 bl[413] br[413] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_414 bl[414] br[414] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_415 bl[415] br[415] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_416 bl[416] br[416] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_417 bl[417] br[417] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_418 bl[418] br[418] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_419 bl[419] br[419] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_420 bl[420] br[420] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_421 bl[421] br[421] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_422 bl[422] br[422] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_423 bl[423] br[423] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_424 bl[424] br[424] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_425 bl[425] br[425] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_426 bl[426] br[426] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_427 bl[427] br[427] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_428 bl[428] br[428] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_429 bl[429] br[429] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_430 bl[430] br[430] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_431 bl[431] br[431] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_432 bl[432] br[432] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_433 bl[433] br[433] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_434 bl[434] br[434] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_435 bl[435] br[435] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_436 bl[436] br[436] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_437 bl[437] br[437] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_438 bl[438] br[438] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_439 bl[439] br[439] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_440 bl[440] br[440] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_441 bl[441] br[441] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_442 bl[442] br[442] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_443 bl[443] br[443] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_444 bl[444] br[444] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_445 bl[445] br[445] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_446 bl[446] br[446] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_447 bl[447] br[447] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_448 bl[448] br[448] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_449 bl[449] br[449] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_450 bl[450] br[450] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_451 bl[451] br[451] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_452 bl[452] br[452] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_453 bl[453] br[453] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_454 bl[454] br[454] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_455 bl[455] br[455] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_456 bl[456] br[456] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_457 bl[457] br[457] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_458 bl[458] br[458] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_459 bl[459] br[459] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_460 bl[460] br[460] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_461 bl[461] br[461] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_462 bl[462] br[462] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_463 bl[463] br[463] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_464 bl[464] br[464] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_465 bl[465] br[465] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_466 bl[466] br[466] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_467 bl[467] br[467] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_468 bl[468] br[468] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_469 bl[469] br[469] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_470 bl[470] br[470] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_471 bl[471] br[471] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_472 bl[472] br[472] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_473 bl[473] br[473] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_474 bl[474] br[474] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_475 bl[475] br[475] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_476 bl[476] br[476] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_477 bl[477] br[477] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_478 bl[478] br[478] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_479 bl[479] br[479] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_480 bl[480] br[480] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_481 bl[481] br[481] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_482 bl[482] br[482] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_483 bl[483] br[483] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_484 bl[484] br[484] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_485 bl[485] br[485] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_486 bl[486] br[486] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_487 bl[487] br[487] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_488 bl[488] br[488] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_489 bl[489] br[489] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_490 bl[490] br[490] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_491 bl[491] br[491] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_492 bl[492] br[492] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_493 bl[493] br[493] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_494 bl[494] br[494] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_495 bl[495] br[495] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_496 bl[496] br[496] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_497 bl[497] br[497] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_498 bl[498] br[498] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_499 bl[499] br[499] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_500 bl[500] br[500] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_501 bl[501] br[501] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_502 bl[502] br[502] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_503 bl[503] br[503] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_504 bl[504] br[504] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_505 bl[505] br[505] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_506 bl[506] br[506] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_507 bl[507] br[507] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_508 bl[508] br[508] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_509 bl[509] br[509] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_510 bl[510] br[510] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_32_511 bl[511] br[511] vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xcell_33_0 bl[0] br[0] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_1 bl[1] br[1] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_2 bl[2] br[2] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_3 bl[3] br[3] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_4 bl[4] br[4] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_5 bl[5] br[5] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_6 bl[6] br[6] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_7 bl[7] br[7] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_8 bl[8] br[8] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_9 bl[9] br[9] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_10 bl[10] br[10] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_11 bl[11] br[11] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_12 bl[12] br[12] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_13 bl[13] br[13] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_14 bl[14] br[14] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_15 bl[15] br[15] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_16 bl[16] br[16] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_17 bl[17] br[17] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_18 bl[18] br[18] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_19 bl[19] br[19] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_20 bl[20] br[20] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_21 bl[21] br[21] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_22 bl[22] br[22] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_23 bl[23] br[23] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_24 bl[24] br[24] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_25 bl[25] br[25] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_26 bl[26] br[26] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_27 bl[27] br[27] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_28 bl[28] br[28] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_29 bl[29] br[29] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_30 bl[30] br[30] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_31 bl[31] br[31] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_32 bl[32] br[32] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_33 bl[33] br[33] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_34 bl[34] br[34] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_35 bl[35] br[35] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_36 bl[36] br[36] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_37 bl[37] br[37] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_38 bl[38] br[38] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_39 bl[39] br[39] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_40 bl[40] br[40] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_41 bl[41] br[41] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_42 bl[42] br[42] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_43 bl[43] br[43] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_44 bl[44] br[44] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_45 bl[45] br[45] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_46 bl[46] br[46] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_47 bl[47] br[47] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_48 bl[48] br[48] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_49 bl[49] br[49] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_50 bl[50] br[50] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_51 bl[51] br[51] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_52 bl[52] br[52] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_53 bl[53] br[53] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_54 bl[54] br[54] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_55 bl[55] br[55] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_56 bl[56] br[56] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_57 bl[57] br[57] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_58 bl[58] br[58] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_59 bl[59] br[59] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_60 bl[60] br[60] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_61 bl[61] br[61] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_62 bl[62] br[62] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_63 bl[63] br[63] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_64 bl[64] br[64] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_65 bl[65] br[65] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_66 bl[66] br[66] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_67 bl[67] br[67] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_68 bl[68] br[68] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_69 bl[69] br[69] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_70 bl[70] br[70] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_71 bl[71] br[71] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_72 bl[72] br[72] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_73 bl[73] br[73] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_74 bl[74] br[74] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_75 bl[75] br[75] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_76 bl[76] br[76] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_77 bl[77] br[77] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_78 bl[78] br[78] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_79 bl[79] br[79] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_80 bl[80] br[80] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_81 bl[81] br[81] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_82 bl[82] br[82] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_83 bl[83] br[83] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_84 bl[84] br[84] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_85 bl[85] br[85] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_86 bl[86] br[86] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_87 bl[87] br[87] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_88 bl[88] br[88] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_89 bl[89] br[89] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_90 bl[90] br[90] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_91 bl[91] br[91] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_92 bl[92] br[92] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_93 bl[93] br[93] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_94 bl[94] br[94] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_95 bl[95] br[95] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_96 bl[96] br[96] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_97 bl[97] br[97] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_98 bl[98] br[98] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_99 bl[99] br[99] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_100 bl[100] br[100] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_101 bl[101] br[101] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_102 bl[102] br[102] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_103 bl[103] br[103] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_104 bl[104] br[104] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_105 bl[105] br[105] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_106 bl[106] br[106] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_107 bl[107] br[107] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_108 bl[108] br[108] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_109 bl[109] br[109] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_110 bl[110] br[110] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_111 bl[111] br[111] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_112 bl[112] br[112] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_113 bl[113] br[113] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_114 bl[114] br[114] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_115 bl[115] br[115] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_116 bl[116] br[116] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_117 bl[117] br[117] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_118 bl[118] br[118] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_119 bl[119] br[119] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_120 bl[120] br[120] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_121 bl[121] br[121] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_122 bl[122] br[122] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_123 bl[123] br[123] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_124 bl[124] br[124] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_125 bl[125] br[125] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_126 bl[126] br[126] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_127 bl[127] br[127] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_128 bl[128] br[128] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_129 bl[129] br[129] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_130 bl[130] br[130] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_131 bl[131] br[131] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_132 bl[132] br[132] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_133 bl[133] br[133] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_134 bl[134] br[134] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_135 bl[135] br[135] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_136 bl[136] br[136] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_137 bl[137] br[137] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_138 bl[138] br[138] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_139 bl[139] br[139] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_140 bl[140] br[140] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_141 bl[141] br[141] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_142 bl[142] br[142] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_143 bl[143] br[143] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_144 bl[144] br[144] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_145 bl[145] br[145] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_146 bl[146] br[146] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_147 bl[147] br[147] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_148 bl[148] br[148] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_149 bl[149] br[149] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_150 bl[150] br[150] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_151 bl[151] br[151] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_152 bl[152] br[152] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_153 bl[153] br[153] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_154 bl[154] br[154] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_155 bl[155] br[155] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_156 bl[156] br[156] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_157 bl[157] br[157] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_158 bl[158] br[158] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_159 bl[159] br[159] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_160 bl[160] br[160] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_161 bl[161] br[161] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_162 bl[162] br[162] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_163 bl[163] br[163] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_164 bl[164] br[164] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_165 bl[165] br[165] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_166 bl[166] br[166] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_167 bl[167] br[167] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_168 bl[168] br[168] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_169 bl[169] br[169] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_170 bl[170] br[170] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_171 bl[171] br[171] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_172 bl[172] br[172] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_173 bl[173] br[173] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_174 bl[174] br[174] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_175 bl[175] br[175] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_176 bl[176] br[176] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_177 bl[177] br[177] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_178 bl[178] br[178] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_179 bl[179] br[179] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_180 bl[180] br[180] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_181 bl[181] br[181] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_182 bl[182] br[182] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_183 bl[183] br[183] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_184 bl[184] br[184] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_185 bl[185] br[185] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_186 bl[186] br[186] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_187 bl[187] br[187] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_188 bl[188] br[188] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_189 bl[189] br[189] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_190 bl[190] br[190] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_191 bl[191] br[191] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_192 bl[192] br[192] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_193 bl[193] br[193] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_194 bl[194] br[194] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_195 bl[195] br[195] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_196 bl[196] br[196] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_197 bl[197] br[197] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_198 bl[198] br[198] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_199 bl[199] br[199] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_200 bl[200] br[200] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_201 bl[201] br[201] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_202 bl[202] br[202] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_203 bl[203] br[203] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_204 bl[204] br[204] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_205 bl[205] br[205] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_206 bl[206] br[206] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_207 bl[207] br[207] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_208 bl[208] br[208] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_209 bl[209] br[209] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_210 bl[210] br[210] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_211 bl[211] br[211] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_212 bl[212] br[212] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_213 bl[213] br[213] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_214 bl[214] br[214] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_215 bl[215] br[215] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_216 bl[216] br[216] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_217 bl[217] br[217] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_218 bl[218] br[218] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_219 bl[219] br[219] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_220 bl[220] br[220] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_221 bl[221] br[221] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_222 bl[222] br[222] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_223 bl[223] br[223] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_224 bl[224] br[224] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_225 bl[225] br[225] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_226 bl[226] br[226] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_227 bl[227] br[227] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_228 bl[228] br[228] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_229 bl[229] br[229] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_230 bl[230] br[230] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_231 bl[231] br[231] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_232 bl[232] br[232] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_233 bl[233] br[233] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_234 bl[234] br[234] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_235 bl[235] br[235] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_236 bl[236] br[236] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_237 bl[237] br[237] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_238 bl[238] br[238] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_239 bl[239] br[239] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_240 bl[240] br[240] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_241 bl[241] br[241] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_242 bl[242] br[242] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_243 bl[243] br[243] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_244 bl[244] br[244] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_245 bl[245] br[245] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_246 bl[246] br[246] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_247 bl[247] br[247] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_248 bl[248] br[248] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_249 bl[249] br[249] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_250 bl[250] br[250] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_251 bl[251] br[251] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_252 bl[252] br[252] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_253 bl[253] br[253] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_254 bl[254] br[254] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_255 bl[255] br[255] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_256 bl[256] br[256] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_257 bl[257] br[257] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_258 bl[258] br[258] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_259 bl[259] br[259] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_260 bl[260] br[260] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_261 bl[261] br[261] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_262 bl[262] br[262] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_263 bl[263] br[263] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_264 bl[264] br[264] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_265 bl[265] br[265] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_266 bl[266] br[266] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_267 bl[267] br[267] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_268 bl[268] br[268] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_269 bl[269] br[269] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_270 bl[270] br[270] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_271 bl[271] br[271] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_272 bl[272] br[272] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_273 bl[273] br[273] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_274 bl[274] br[274] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_275 bl[275] br[275] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_276 bl[276] br[276] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_277 bl[277] br[277] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_278 bl[278] br[278] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_279 bl[279] br[279] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_280 bl[280] br[280] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_281 bl[281] br[281] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_282 bl[282] br[282] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_283 bl[283] br[283] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_284 bl[284] br[284] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_285 bl[285] br[285] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_286 bl[286] br[286] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_287 bl[287] br[287] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_288 bl[288] br[288] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_289 bl[289] br[289] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_290 bl[290] br[290] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_291 bl[291] br[291] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_292 bl[292] br[292] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_293 bl[293] br[293] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_294 bl[294] br[294] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_295 bl[295] br[295] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_296 bl[296] br[296] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_297 bl[297] br[297] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_298 bl[298] br[298] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_299 bl[299] br[299] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_300 bl[300] br[300] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_301 bl[301] br[301] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_302 bl[302] br[302] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_303 bl[303] br[303] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_304 bl[304] br[304] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_305 bl[305] br[305] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_306 bl[306] br[306] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_307 bl[307] br[307] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_308 bl[308] br[308] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_309 bl[309] br[309] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_310 bl[310] br[310] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_311 bl[311] br[311] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_312 bl[312] br[312] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_313 bl[313] br[313] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_314 bl[314] br[314] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_315 bl[315] br[315] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_316 bl[316] br[316] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_317 bl[317] br[317] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_318 bl[318] br[318] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_319 bl[319] br[319] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_320 bl[320] br[320] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_321 bl[321] br[321] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_322 bl[322] br[322] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_323 bl[323] br[323] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_324 bl[324] br[324] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_325 bl[325] br[325] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_326 bl[326] br[326] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_327 bl[327] br[327] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_328 bl[328] br[328] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_329 bl[329] br[329] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_330 bl[330] br[330] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_331 bl[331] br[331] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_332 bl[332] br[332] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_333 bl[333] br[333] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_334 bl[334] br[334] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_335 bl[335] br[335] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_336 bl[336] br[336] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_337 bl[337] br[337] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_338 bl[338] br[338] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_339 bl[339] br[339] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_340 bl[340] br[340] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_341 bl[341] br[341] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_342 bl[342] br[342] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_343 bl[343] br[343] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_344 bl[344] br[344] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_345 bl[345] br[345] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_346 bl[346] br[346] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_347 bl[347] br[347] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_348 bl[348] br[348] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_349 bl[349] br[349] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_350 bl[350] br[350] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_351 bl[351] br[351] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_352 bl[352] br[352] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_353 bl[353] br[353] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_354 bl[354] br[354] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_355 bl[355] br[355] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_356 bl[356] br[356] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_357 bl[357] br[357] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_358 bl[358] br[358] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_359 bl[359] br[359] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_360 bl[360] br[360] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_361 bl[361] br[361] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_362 bl[362] br[362] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_363 bl[363] br[363] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_364 bl[364] br[364] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_365 bl[365] br[365] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_366 bl[366] br[366] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_367 bl[367] br[367] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_368 bl[368] br[368] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_369 bl[369] br[369] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_370 bl[370] br[370] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_371 bl[371] br[371] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_372 bl[372] br[372] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_373 bl[373] br[373] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_374 bl[374] br[374] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_375 bl[375] br[375] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_376 bl[376] br[376] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_377 bl[377] br[377] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_378 bl[378] br[378] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_379 bl[379] br[379] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_380 bl[380] br[380] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_381 bl[381] br[381] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_382 bl[382] br[382] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_383 bl[383] br[383] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_384 bl[384] br[384] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_385 bl[385] br[385] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_386 bl[386] br[386] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_387 bl[387] br[387] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_388 bl[388] br[388] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_389 bl[389] br[389] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_390 bl[390] br[390] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_391 bl[391] br[391] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_392 bl[392] br[392] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_393 bl[393] br[393] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_394 bl[394] br[394] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_395 bl[395] br[395] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_396 bl[396] br[396] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_397 bl[397] br[397] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_398 bl[398] br[398] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_399 bl[399] br[399] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_400 bl[400] br[400] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_401 bl[401] br[401] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_402 bl[402] br[402] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_403 bl[403] br[403] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_404 bl[404] br[404] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_405 bl[405] br[405] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_406 bl[406] br[406] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_407 bl[407] br[407] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_408 bl[408] br[408] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_409 bl[409] br[409] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_410 bl[410] br[410] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_411 bl[411] br[411] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_412 bl[412] br[412] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_413 bl[413] br[413] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_414 bl[414] br[414] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_415 bl[415] br[415] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_416 bl[416] br[416] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_417 bl[417] br[417] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_418 bl[418] br[418] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_419 bl[419] br[419] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_420 bl[420] br[420] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_421 bl[421] br[421] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_422 bl[422] br[422] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_423 bl[423] br[423] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_424 bl[424] br[424] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_425 bl[425] br[425] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_426 bl[426] br[426] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_427 bl[427] br[427] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_428 bl[428] br[428] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_429 bl[429] br[429] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_430 bl[430] br[430] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_431 bl[431] br[431] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_432 bl[432] br[432] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_433 bl[433] br[433] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_434 bl[434] br[434] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_435 bl[435] br[435] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_436 bl[436] br[436] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_437 bl[437] br[437] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_438 bl[438] br[438] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_439 bl[439] br[439] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_440 bl[440] br[440] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_441 bl[441] br[441] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_442 bl[442] br[442] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_443 bl[443] br[443] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_444 bl[444] br[444] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_445 bl[445] br[445] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_446 bl[446] br[446] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_447 bl[447] br[447] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_448 bl[448] br[448] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_449 bl[449] br[449] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_450 bl[450] br[450] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_451 bl[451] br[451] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_452 bl[452] br[452] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_453 bl[453] br[453] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_454 bl[454] br[454] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_455 bl[455] br[455] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_456 bl[456] br[456] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_457 bl[457] br[457] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_458 bl[458] br[458] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_459 bl[459] br[459] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_460 bl[460] br[460] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_461 bl[461] br[461] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_462 bl[462] br[462] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_463 bl[463] br[463] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_464 bl[464] br[464] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_465 bl[465] br[465] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_466 bl[466] br[466] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_467 bl[467] br[467] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_468 bl[468] br[468] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_469 bl[469] br[469] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_470 bl[470] br[470] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_471 bl[471] br[471] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_472 bl[472] br[472] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_473 bl[473] br[473] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_474 bl[474] br[474] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_475 bl[475] br[475] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_476 bl[476] br[476] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_477 bl[477] br[477] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_478 bl[478] br[478] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_479 bl[479] br[479] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_480 bl[480] br[480] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_481 bl[481] br[481] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_482 bl[482] br[482] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_483 bl[483] br[483] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_484 bl[484] br[484] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_485 bl[485] br[485] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_486 bl[486] br[486] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_487 bl[487] br[487] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_488 bl[488] br[488] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_489 bl[489] br[489] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_490 bl[490] br[490] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_491 bl[491] br[491] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_492 bl[492] br[492] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_493 bl[493] br[493] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_494 bl[494] br[494] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_495 bl[495] br[495] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_496 bl[496] br[496] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_497 bl[497] br[497] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_498 bl[498] br[498] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_499 bl[499] br[499] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_500 bl[500] br[500] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_501 bl[501] br[501] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_502 bl[502] br[502] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_503 bl[503] br[503] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_504 bl[504] br[504] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_505 bl[505] br[505] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_506 bl[506] br[506] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_507 bl[507] br[507] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_508 bl[508] br[508] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_509 bl[509] br[509] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_510 bl[510] br[510] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_33_511 bl[511] br[511] vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xcell_34_0 bl[0] br[0] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_1 bl[1] br[1] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_2 bl[2] br[2] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_3 bl[3] br[3] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_4 bl[4] br[4] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_5 bl[5] br[5] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_6 bl[6] br[6] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_7 bl[7] br[7] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_8 bl[8] br[8] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_9 bl[9] br[9] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_10 bl[10] br[10] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_11 bl[11] br[11] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_12 bl[12] br[12] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_13 bl[13] br[13] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_14 bl[14] br[14] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_15 bl[15] br[15] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_16 bl[16] br[16] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_17 bl[17] br[17] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_18 bl[18] br[18] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_19 bl[19] br[19] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_20 bl[20] br[20] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_21 bl[21] br[21] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_22 bl[22] br[22] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_23 bl[23] br[23] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_24 bl[24] br[24] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_25 bl[25] br[25] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_26 bl[26] br[26] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_27 bl[27] br[27] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_28 bl[28] br[28] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_29 bl[29] br[29] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_30 bl[30] br[30] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_31 bl[31] br[31] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_32 bl[32] br[32] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_33 bl[33] br[33] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_34 bl[34] br[34] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_35 bl[35] br[35] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_36 bl[36] br[36] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_37 bl[37] br[37] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_38 bl[38] br[38] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_39 bl[39] br[39] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_40 bl[40] br[40] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_41 bl[41] br[41] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_42 bl[42] br[42] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_43 bl[43] br[43] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_44 bl[44] br[44] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_45 bl[45] br[45] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_46 bl[46] br[46] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_47 bl[47] br[47] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_48 bl[48] br[48] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_49 bl[49] br[49] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_50 bl[50] br[50] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_51 bl[51] br[51] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_52 bl[52] br[52] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_53 bl[53] br[53] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_54 bl[54] br[54] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_55 bl[55] br[55] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_56 bl[56] br[56] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_57 bl[57] br[57] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_58 bl[58] br[58] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_59 bl[59] br[59] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_60 bl[60] br[60] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_61 bl[61] br[61] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_62 bl[62] br[62] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_63 bl[63] br[63] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_64 bl[64] br[64] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_65 bl[65] br[65] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_66 bl[66] br[66] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_67 bl[67] br[67] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_68 bl[68] br[68] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_69 bl[69] br[69] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_70 bl[70] br[70] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_71 bl[71] br[71] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_72 bl[72] br[72] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_73 bl[73] br[73] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_74 bl[74] br[74] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_75 bl[75] br[75] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_76 bl[76] br[76] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_77 bl[77] br[77] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_78 bl[78] br[78] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_79 bl[79] br[79] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_80 bl[80] br[80] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_81 bl[81] br[81] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_82 bl[82] br[82] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_83 bl[83] br[83] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_84 bl[84] br[84] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_85 bl[85] br[85] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_86 bl[86] br[86] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_87 bl[87] br[87] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_88 bl[88] br[88] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_89 bl[89] br[89] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_90 bl[90] br[90] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_91 bl[91] br[91] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_92 bl[92] br[92] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_93 bl[93] br[93] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_94 bl[94] br[94] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_95 bl[95] br[95] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_96 bl[96] br[96] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_97 bl[97] br[97] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_98 bl[98] br[98] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_99 bl[99] br[99] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_100 bl[100] br[100] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_101 bl[101] br[101] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_102 bl[102] br[102] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_103 bl[103] br[103] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_104 bl[104] br[104] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_105 bl[105] br[105] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_106 bl[106] br[106] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_107 bl[107] br[107] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_108 bl[108] br[108] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_109 bl[109] br[109] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_110 bl[110] br[110] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_111 bl[111] br[111] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_112 bl[112] br[112] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_113 bl[113] br[113] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_114 bl[114] br[114] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_115 bl[115] br[115] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_116 bl[116] br[116] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_117 bl[117] br[117] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_118 bl[118] br[118] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_119 bl[119] br[119] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_120 bl[120] br[120] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_121 bl[121] br[121] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_122 bl[122] br[122] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_123 bl[123] br[123] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_124 bl[124] br[124] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_125 bl[125] br[125] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_126 bl[126] br[126] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_127 bl[127] br[127] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_128 bl[128] br[128] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_129 bl[129] br[129] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_130 bl[130] br[130] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_131 bl[131] br[131] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_132 bl[132] br[132] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_133 bl[133] br[133] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_134 bl[134] br[134] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_135 bl[135] br[135] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_136 bl[136] br[136] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_137 bl[137] br[137] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_138 bl[138] br[138] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_139 bl[139] br[139] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_140 bl[140] br[140] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_141 bl[141] br[141] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_142 bl[142] br[142] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_143 bl[143] br[143] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_144 bl[144] br[144] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_145 bl[145] br[145] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_146 bl[146] br[146] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_147 bl[147] br[147] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_148 bl[148] br[148] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_149 bl[149] br[149] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_150 bl[150] br[150] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_151 bl[151] br[151] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_152 bl[152] br[152] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_153 bl[153] br[153] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_154 bl[154] br[154] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_155 bl[155] br[155] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_156 bl[156] br[156] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_157 bl[157] br[157] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_158 bl[158] br[158] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_159 bl[159] br[159] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_160 bl[160] br[160] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_161 bl[161] br[161] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_162 bl[162] br[162] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_163 bl[163] br[163] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_164 bl[164] br[164] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_165 bl[165] br[165] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_166 bl[166] br[166] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_167 bl[167] br[167] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_168 bl[168] br[168] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_169 bl[169] br[169] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_170 bl[170] br[170] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_171 bl[171] br[171] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_172 bl[172] br[172] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_173 bl[173] br[173] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_174 bl[174] br[174] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_175 bl[175] br[175] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_176 bl[176] br[176] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_177 bl[177] br[177] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_178 bl[178] br[178] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_179 bl[179] br[179] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_180 bl[180] br[180] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_181 bl[181] br[181] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_182 bl[182] br[182] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_183 bl[183] br[183] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_184 bl[184] br[184] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_185 bl[185] br[185] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_186 bl[186] br[186] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_187 bl[187] br[187] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_188 bl[188] br[188] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_189 bl[189] br[189] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_190 bl[190] br[190] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_191 bl[191] br[191] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_192 bl[192] br[192] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_193 bl[193] br[193] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_194 bl[194] br[194] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_195 bl[195] br[195] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_196 bl[196] br[196] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_197 bl[197] br[197] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_198 bl[198] br[198] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_199 bl[199] br[199] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_200 bl[200] br[200] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_201 bl[201] br[201] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_202 bl[202] br[202] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_203 bl[203] br[203] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_204 bl[204] br[204] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_205 bl[205] br[205] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_206 bl[206] br[206] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_207 bl[207] br[207] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_208 bl[208] br[208] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_209 bl[209] br[209] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_210 bl[210] br[210] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_211 bl[211] br[211] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_212 bl[212] br[212] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_213 bl[213] br[213] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_214 bl[214] br[214] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_215 bl[215] br[215] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_216 bl[216] br[216] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_217 bl[217] br[217] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_218 bl[218] br[218] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_219 bl[219] br[219] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_220 bl[220] br[220] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_221 bl[221] br[221] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_222 bl[222] br[222] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_223 bl[223] br[223] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_224 bl[224] br[224] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_225 bl[225] br[225] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_226 bl[226] br[226] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_227 bl[227] br[227] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_228 bl[228] br[228] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_229 bl[229] br[229] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_230 bl[230] br[230] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_231 bl[231] br[231] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_232 bl[232] br[232] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_233 bl[233] br[233] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_234 bl[234] br[234] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_235 bl[235] br[235] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_236 bl[236] br[236] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_237 bl[237] br[237] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_238 bl[238] br[238] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_239 bl[239] br[239] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_240 bl[240] br[240] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_241 bl[241] br[241] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_242 bl[242] br[242] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_243 bl[243] br[243] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_244 bl[244] br[244] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_245 bl[245] br[245] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_246 bl[246] br[246] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_247 bl[247] br[247] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_248 bl[248] br[248] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_249 bl[249] br[249] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_250 bl[250] br[250] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_251 bl[251] br[251] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_252 bl[252] br[252] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_253 bl[253] br[253] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_254 bl[254] br[254] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_255 bl[255] br[255] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_256 bl[256] br[256] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_257 bl[257] br[257] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_258 bl[258] br[258] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_259 bl[259] br[259] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_260 bl[260] br[260] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_261 bl[261] br[261] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_262 bl[262] br[262] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_263 bl[263] br[263] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_264 bl[264] br[264] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_265 bl[265] br[265] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_266 bl[266] br[266] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_267 bl[267] br[267] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_268 bl[268] br[268] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_269 bl[269] br[269] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_270 bl[270] br[270] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_271 bl[271] br[271] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_272 bl[272] br[272] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_273 bl[273] br[273] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_274 bl[274] br[274] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_275 bl[275] br[275] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_276 bl[276] br[276] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_277 bl[277] br[277] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_278 bl[278] br[278] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_279 bl[279] br[279] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_280 bl[280] br[280] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_281 bl[281] br[281] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_282 bl[282] br[282] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_283 bl[283] br[283] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_284 bl[284] br[284] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_285 bl[285] br[285] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_286 bl[286] br[286] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_287 bl[287] br[287] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_288 bl[288] br[288] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_289 bl[289] br[289] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_290 bl[290] br[290] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_291 bl[291] br[291] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_292 bl[292] br[292] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_293 bl[293] br[293] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_294 bl[294] br[294] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_295 bl[295] br[295] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_296 bl[296] br[296] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_297 bl[297] br[297] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_298 bl[298] br[298] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_299 bl[299] br[299] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_300 bl[300] br[300] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_301 bl[301] br[301] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_302 bl[302] br[302] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_303 bl[303] br[303] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_304 bl[304] br[304] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_305 bl[305] br[305] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_306 bl[306] br[306] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_307 bl[307] br[307] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_308 bl[308] br[308] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_309 bl[309] br[309] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_310 bl[310] br[310] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_311 bl[311] br[311] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_312 bl[312] br[312] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_313 bl[313] br[313] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_314 bl[314] br[314] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_315 bl[315] br[315] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_316 bl[316] br[316] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_317 bl[317] br[317] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_318 bl[318] br[318] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_319 bl[319] br[319] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_320 bl[320] br[320] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_321 bl[321] br[321] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_322 bl[322] br[322] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_323 bl[323] br[323] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_324 bl[324] br[324] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_325 bl[325] br[325] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_326 bl[326] br[326] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_327 bl[327] br[327] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_328 bl[328] br[328] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_329 bl[329] br[329] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_330 bl[330] br[330] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_331 bl[331] br[331] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_332 bl[332] br[332] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_333 bl[333] br[333] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_334 bl[334] br[334] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_335 bl[335] br[335] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_336 bl[336] br[336] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_337 bl[337] br[337] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_338 bl[338] br[338] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_339 bl[339] br[339] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_340 bl[340] br[340] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_341 bl[341] br[341] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_342 bl[342] br[342] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_343 bl[343] br[343] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_344 bl[344] br[344] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_345 bl[345] br[345] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_346 bl[346] br[346] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_347 bl[347] br[347] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_348 bl[348] br[348] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_349 bl[349] br[349] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_350 bl[350] br[350] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_351 bl[351] br[351] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_352 bl[352] br[352] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_353 bl[353] br[353] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_354 bl[354] br[354] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_355 bl[355] br[355] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_356 bl[356] br[356] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_357 bl[357] br[357] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_358 bl[358] br[358] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_359 bl[359] br[359] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_360 bl[360] br[360] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_361 bl[361] br[361] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_362 bl[362] br[362] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_363 bl[363] br[363] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_364 bl[364] br[364] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_365 bl[365] br[365] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_366 bl[366] br[366] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_367 bl[367] br[367] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_368 bl[368] br[368] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_369 bl[369] br[369] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_370 bl[370] br[370] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_371 bl[371] br[371] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_372 bl[372] br[372] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_373 bl[373] br[373] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_374 bl[374] br[374] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_375 bl[375] br[375] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_376 bl[376] br[376] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_377 bl[377] br[377] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_378 bl[378] br[378] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_379 bl[379] br[379] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_380 bl[380] br[380] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_381 bl[381] br[381] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_382 bl[382] br[382] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_383 bl[383] br[383] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_384 bl[384] br[384] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_385 bl[385] br[385] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_386 bl[386] br[386] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_387 bl[387] br[387] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_388 bl[388] br[388] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_389 bl[389] br[389] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_390 bl[390] br[390] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_391 bl[391] br[391] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_392 bl[392] br[392] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_393 bl[393] br[393] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_394 bl[394] br[394] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_395 bl[395] br[395] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_396 bl[396] br[396] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_397 bl[397] br[397] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_398 bl[398] br[398] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_399 bl[399] br[399] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_400 bl[400] br[400] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_401 bl[401] br[401] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_402 bl[402] br[402] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_403 bl[403] br[403] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_404 bl[404] br[404] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_405 bl[405] br[405] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_406 bl[406] br[406] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_407 bl[407] br[407] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_408 bl[408] br[408] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_409 bl[409] br[409] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_410 bl[410] br[410] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_411 bl[411] br[411] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_412 bl[412] br[412] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_413 bl[413] br[413] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_414 bl[414] br[414] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_415 bl[415] br[415] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_416 bl[416] br[416] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_417 bl[417] br[417] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_418 bl[418] br[418] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_419 bl[419] br[419] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_420 bl[420] br[420] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_421 bl[421] br[421] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_422 bl[422] br[422] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_423 bl[423] br[423] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_424 bl[424] br[424] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_425 bl[425] br[425] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_426 bl[426] br[426] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_427 bl[427] br[427] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_428 bl[428] br[428] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_429 bl[429] br[429] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_430 bl[430] br[430] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_431 bl[431] br[431] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_432 bl[432] br[432] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_433 bl[433] br[433] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_434 bl[434] br[434] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_435 bl[435] br[435] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_436 bl[436] br[436] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_437 bl[437] br[437] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_438 bl[438] br[438] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_439 bl[439] br[439] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_440 bl[440] br[440] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_441 bl[441] br[441] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_442 bl[442] br[442] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_443 bl[443] br[443] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_444 bl[444] br[444] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_445 bl[445] br[445] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_446 bl[446] br[446] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_447 bl[447] br[447] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_448 bl[448] br[448] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_449 bl[449] br[449] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_450 bl[450] br[450] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_451 bl[451] br[451] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_452 bl[452] br[452] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_453 bl[453] br[453] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_454 bl[454] br[454] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_455 bl[455] br[455] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_456 bl[456] br[456] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_457 bl[457] br[457] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_458 bl[458] br[458] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_459 bl[459] br[459] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_460 bl[460] br[460] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_461 bl[461] br[461] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_462 bl[462] br[462] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_463 bl[463] br[463] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_464 bl[464] br[464] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_465 bl[465] br[465] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_466 bl[466] br[466] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_467 bl[467] br[467] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_468 bl[468] br[468] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_469 bl[469] br[469] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_470 bl[470] br[470] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_471 bl[471] br[471] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_472 bl[472] br[472] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_473 bl[473] br[473] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_474 bl[474] br[474] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_475 bl[475] br[475] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_476 bl[476] br[476] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_477 bl[477] br[477] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_478 bl[478] br[478] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_479 bl[479] br[479] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_480 bl[480] br[480] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_481 bl[481] br[481] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_482 bl[482] br[482] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_483 bl[483] br[483] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_484 bl[484] br[484] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_485 bl[485] br[485] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_486 bl[486] br[486] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_487 bl[487] br[487] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_488 bl[488] br[488] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_489 bl[489] br[489] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_490 bl[490] br[490] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_491 bl[491] br[491] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_492 bl[492] br[492] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_493 bl[493] br[493] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_494 bl[494] br[494] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_495 bl[495] br[495] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_496 bl[496] br[496] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_497 bl[497] br[497] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_498 bl[498] br[498] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_499 bl[499] br[499] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_500 bl[500] br[500] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_501 bl[501] br[501] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_502 bl[502] br[502] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_503 bl[503] br[503] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_504 bl[504] br[504] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_505 bl[505] br[505] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_506 bl[506] br[506] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_507 bl[507] br[507] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_508 bl[508] br[508] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_509 bl[509] br[509] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_510 bl[510] br[510] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_34_511 bl[511] br[511] vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xcell_35_0 bl[0] br[0] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_1 bl[1] br[1] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_2 bl[2] br[2] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_3 bl[3] br[3] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_4 bl[4] br[4] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_5 bl[5] br[5] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_6 bl[6] br[6] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_7 bl[7] br[7] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_8 bl[8] br[8] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_9 bl[9] br[9] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_10 bl[10] br[10] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_11 bl[11] br[11] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_12 bl[12] br[12] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_13 bl[13] br[13] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_14 bl[14] br[14] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_15 bl[15] br[15] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_16 bl[16] br[16] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_17 bl[17] br[17] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_18 bl[18] br[18] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_19 bl[19] br[19] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_20 bl[20] br[20] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_21 bl[21] br[21] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_22 bl[22] br[22] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_23 bl[23] br[23] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_24 bl[24] br[24] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_25 bl[25] br[25] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_26 bl[26] br[26] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_27 bl[27] br[27] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_28 bl[28] br[28] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_29 bl[29] br[29] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_30 bl[30] br[30] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_31 bl[31] br[31] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_32 bl[32] br[32] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_33 bl[33] br[33] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_34 bl[34] br[34] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_35 bl[35] br[35] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_36 bl[36] br[36] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_37 bl[37] br[37] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_38 bl[38] br[38] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_39 bl[39] br[39] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_40 bl[40] br[40] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_41 bl[41] br[41] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_42 bl[42] br[42] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_43 bl[43] br[43] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_44 bl[44] br[44] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_45 bl[45] br[45] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_46 bl[46] br[46] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_47 bl[47] br[47] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_48 bl[48] br[48] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_49 bl[49] br[49] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_50 bl[50] br[50] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_51 bl[51] br[51] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_52 bl[52] br[52] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_53 bl[53] br[53] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_54 bl[54] br[54] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_55 bl[55] br[55] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_56 bl[56] br[56] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_57 bl[57] br[57] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_58 bl[58] br[58] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_59 bl[59] br[59] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_60 bl[60] br[60] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_61 bl[61] br[61] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_62 bl[62] br[62] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_63 bl[63] br[63] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_64 bl[64] br[64] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_65 bl[65] br[65] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_66 bl[66] br[66] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_67 bl[67] br[67] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_68 bl[68] br[68] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_69 bl[69] br[69] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_70 bl[70] br[70] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_71 bl[71] br[71] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_72 bl[72] br[72] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_73 bl[73] br[73] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_74 bl[74] br[74] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_75 bl[75] br[75] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_76 bl[76] br[76] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_77 bl[77] br[77] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_78 bl[78] br[78] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_79 bl[79] br[79] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_80 bl[80] br[80] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_81 bl[81] br[81] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_82 bl[82] br[82] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_83 bl[83] br[83] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_84 bl[84] br[84] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_85 bl[85] br[85] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_86 bl[86] br[86] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_87 bl[87] br[87] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_88 bl[88] br[88] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_89 bl[89] br[89] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_90 bl[90] br[90] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_91 bl[91] br[91] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_92 bl[92] br[92] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_93 bl[93] br[93] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_94 bl[94] br[94] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_95 bl[95] br[95] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_96 bl[96] br[96] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_97 bl[97] br[97] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_98 bl[98] br[98] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_99 bl[99] br[99] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_100 bl[100] br[100] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_101 bl[101] br[101] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_102 bl[102] br[102] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_103 bl[103] br[103] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_104 bl[104] br[104] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_105 bl[105] br[105] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_106 bl[106] br[106] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_107 bl[107] br[107] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_108 bl[108] br[108] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_109 bl[109] br[109] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_110 bl[110] br[110] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_111 bl[111] br[111] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_112 bl[112] br[112] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_113 bl[113] br[113] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_114 bl[114] br[114] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_115 bl[115] br[115] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_116 bl[116] br[116] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_117 bl[117] br[117] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_118 bl[118] br[118] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_119 bl[119] br[119] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_120 bl[120] br[120] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_121 bl[121] br[121] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_122 bl[122] br[122] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_123 bl[123] br[123] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_124 bl[124] br[124] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_125 bl[125] br[125] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_126 bl[126] br[126] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_127 bl[127] br[127] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_128 bl[128] br[128] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_129 bl[129] br[129] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_130 bl[130] br[130] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_131 bl[131] br[131] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_132 bl[132] br[132] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_133 bl[133] br[133] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_134 bl[134] br[134] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_135 bl[135] br[135] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_136 bl[136] br[136] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_137 bl[137] br[137] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_138 bl[138] br[138] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_139 bl[139] br[139] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_140 bl[140] br[140] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_141 bl[141] br[141] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_142 bl[142] br[142] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_143 bl[143] br[143] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_144 bl[144] br[144] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_145 bl[145] br[145] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_146 bl[146] br[146] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_147 bl[147] br[147] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_148 bl[148] br[148] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_149 bl[149] br[149] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_150 bl[150] br[150] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_151 bl[151] br[151] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_152 bl[152] br[152] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_153 bl[153] br[153] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_154 bl[154] br[154] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_155 bl[155] br[155] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_156 bl[156] br[156] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_157 bl[157] br[157] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_158 bl[158] br[158] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_159 bl[159] br[159] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_160 bl[160] br[160] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_161 bl[161] br[161] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_162 bl[162] br[162] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_163 bl[163] br[163] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_164 bl[164] br[164] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_165 bl[165] br[165] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_166 bl[166] br[166] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_167 bl[167] br[167] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_168 bl[168] br[168] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_169 bl[169] br[169] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_170 bl[170] br[170] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_171 bl[171] br[171] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_172 bl[172] br[172] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_173 bl[173] br[173] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_174 bl[174] br[174] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_175 bl[175] br[175] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_176 bl[176] br[176] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_177 bl[177] br[177] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_178 bl[178] br[178] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_179 bl[179] br[179] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_180 bl[180] br[180] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_181 bl[181] br[181] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_182 bl[182] br[182] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_183 bl[183] br[183] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_184 bl[184] br[184] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_185 bl[185] br[185] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_186 bl[186] br[186] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_187 bl[187] br[187] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_188 bl[188] br[188] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_189 bl[189] br[189] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_190 bl[190] br[190] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_191 bl[191] br[191] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_192 bl[192] br[192] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_193 bl[193] br[193] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_194 bl[194] br[194] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_195 bl[195] br[195] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_196 bl[196] br[196] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_197 bl[197] br[197] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_198 bl[198] br[198] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_199 bl[199] br[199] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_200 bl[200] br[200] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_201 bl[201] br[201] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_202 bl[202] br[202] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_203 bl[203] br[203] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_204 bl[204] br[204] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_205 bl[205] br[205] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_206 bl[206] br[206] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_207 bl[207] br[207] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_208 bl[208] br[208] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_209 bl[209] br[209] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_210 bl[210] br[210] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_211 bl[211] br[211] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_212 bl[212] br[212] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_213 bl[213] br[213] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_214 bl[214] br[214] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_215 bl[215] br[215] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_216 bl[216] br[216] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_217 bl[217] br[217] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_218 bl[218] br[218] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_219 bl[219] br[219] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_220 bl[220] br[220] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_221 bl[221] br[221] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_222 bl[222] br[222] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_223 bl[223] br[223] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_224 bl[224] br[224] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_225 bl[225] br[225] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_226 bl[226] br[226] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_227 bl[227] br[227] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_228 bl[228] br[228] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_229 bl[229] br[229] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_230 bl[230] br[230] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_231 bl[231] br[231] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_232 bl[232] br[232] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_233 bl[233] br[233] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_234 bl[234] br[234] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_235 bl[235] br[235] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_236 bl[236] br[236] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_237 bl[237] br[237] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_238 bl[238] br[238] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_239 bl[239] br[239] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_240 bl[240] br[240] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_241 bl[241] br[241] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_242 bl[242] br[242] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_243 bl[243] br[243] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_244 bl[244] br[244] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_245 bl[245] br[245] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_246 bl[246] br[246] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_247 bl[247] br[247] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_248 bl[248] br[248] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_249 bl[249] br[249] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_250 bl[250] br[250] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_251 bl[251] br[251] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_252 bl[252] br[252] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_253 bl[253] br[253] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_254 bl[254] br[254] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_255 bl[255] br[255] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_256 bl[256] br[256] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_257 bl[257] br[257] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_258 bl[258] br[258] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_259 bl[259] br[259] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_260 bl[260] br[260] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_261 bl[261] br[261] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_262 bl[262] br[262] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_263 bl[263] br[263] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_264 bl[264] br[264] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_265 bl[265] br[265] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_266 bl[266] br[266] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_267 bl[267] br[267] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_268 bl[268] br[268] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_269 bl[269] br[269] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_270 bl[270] br[270] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_271 bl[271] br[271] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_272 bl[272] br[272] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_273 bl[273] br[273] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_274 bl[274] br[274] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_275 bl[275] br[275] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_276 bl[276] br[276] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_277 bl[277] br[277] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_278 bl[278] br[278] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_279 bl[279] br[279] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_280 bl[280] br[280] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_281 bl[281] br[281] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_282 bl[282] br[282] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_283 bl[283] br[283] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_284 bl[284] br[284] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_285 bl[285] br[285] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_286 bl[286] br[286] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_287 bl[287] br[287] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_288 bl[288] br[288] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_289 bl[289] br[289] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_290 bl[290] br[290] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_291 bl[291] br[291] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_292 bl[292] br[292] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_293 bl[293] br[293] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_294 bl[294] br[294] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_295 bl[295] br[295] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_296 bl[296] br[296] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_297 bl[297] br[297] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_298 bl[298] br[298] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_299 bl[299] br[299] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_300 bl[300] br[300] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_301 bl[301] br[301] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_302 bl[302] br[302] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_303 bl[303] br[303] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_304 bl[304] br[304] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_305 bl[305] br[305] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_306 bl[306] br[306] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_307 bl[307] br[307] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_308 bl[308] br[308] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_309 bl[309] br[309] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_310 bl[310] br[310] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_311 bl[311] br[311] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_312 bl[312] br[312] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_313 bl[313] br[313] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_314 bl[314] br[314] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_315 bl[315] br[315] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_316 bl[316] br[316] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_317 bl[317] br[317] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_318 bl[318] br[318] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_319 bl[319] br[319] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_320 bl[320] br[320] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_321 bl[321] br[321] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_322 bl[322] br[322] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_323 bl[323] br[323] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_324 bl[324] br[324] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_325 bl[325] br[325] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_326 bl[326] br[326] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_327 bl[327] br[327] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_328 bl[328] br[328] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_329 bl[329] br[329] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_330 bl[330] br[330] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_331 bl[331] br[331] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_332 bl[332] br[332] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_333 bl[333] br[333] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_334 bl[334] br[334] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_335 bl[335] br[335] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_336 bl[336] br[336] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_337 bl[337] br[337] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_338 bl[338] br[338] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_339 bl[339] br[339] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_340 bl[340] br[340] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_341 bl[341] br[341] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_342 bl[342] br[342] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_343 bl[343] br[343] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_344 bl[344] br[344] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_345 bl[345] br[345] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_346 bl[346] br[346] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_347 bl[347] br[347] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_348 bl[348] br[348] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_349 bl[349] br[349] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_350 bl[350] br[350] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_351 bl[351] br[351] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_352 bl[352] br[352] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_353 bl[353] br[353] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_354 bl[354] br[354] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_355 bl[355] br[355] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_356 bl[356] br[356] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_357 bl[357] br[357] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_358 bl[358] br[358] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_359 bl[359] br[359] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_360 bl[360] br[360] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_361 bl[361] br[361] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_362 bl[362] br[362] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_363 bl[363] br[363] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_364 bl[364] br[364] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_365 bl[365] br[365] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_366 bl[366] br[366] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_367 bl[367] br[367] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_368 bl[368] br[368] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_369 bl[369] br[369] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_370 bl[370] br[370] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_371 bl[371] br[371] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_372 bl[372] br[372] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_373 bl[373] br[373] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_374 bl[374] br[374] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_375 bl[375] br[375] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_376 bl[376] br[376] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_377 bl[377] br[377] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_378 bl[378] br[378] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_379 bl[379] br[379] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_380 bl[380] br[380] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_381 bl[381] br[381] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_382 bl[382] br[382] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_383 bl[383] br[383] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_384 bl[384] br[384] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_385 bl[385] br[385] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_386 bl[386] br[386] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_387 bl[387] br[387] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_388 bl[388] br[388] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_389 bl[389] br[389] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_390 bl[390] br[390] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_391 bl[391] br[391] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_392 bl[392] br[392] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_393 bl[393] br[393] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_394 bl[394] br[394] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_395 bl[395] br[395] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_396 bl[396] br[396] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_397 bl[397] br[397] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_398 bl[398] br[398] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_399 bl[399] br[399] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_400 bl[400] br[400] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_401 bl[401] br[401] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_402 bl[402] br[402] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_403 bl[403] br[403] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_404 bl[404] br[404] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_405 bl[405] br[405] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_406 bl[406] br[406] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_407 bl[407] br[407] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_408 bl[408] br[408] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_409 bl[409] br[409] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_410 bl[410] br[410] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_411 bl[411] br[411] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_412 bl[412] br[412] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_413 bl[413] br[413] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_414 bl[414] br[414] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_415 bl[415] br[415] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_416 bl[416] br[416] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_417 bl[417] br[417] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_418 bl[418] br[418] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_419 bl[419] br[419] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_420 bl[420] br[420] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_421 bl[421] br[421] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_422 bl[422] br[422] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_423 bl[423] br[423] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_424 bl[424] br[424] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_425 bl[425] br[425] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_426 bl[426] br[426] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_427 bl[427] br[427] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_428 bl[428] br[428] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_429 bl[429] br[429] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_430 bl[430] br[430] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_431 bl[431] br[431] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_432 bl[432] br[432] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_433 bl[433] br[433] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_434 bl[434] br[434] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_435 bl[435] br[435] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_436 bl[436] br[436] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_437 bl[437] br[437] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_438 bl[438] br[438] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_439 bl[439] br[439] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_440 bl[440] br[440] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_441 bl[441] br[441] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_442 bl[442] br[442] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_443 bl[443] br[443] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_444 bl[444] br[444] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_445 bl[445] br[445] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_446 bl[446] br[446] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_447 bl[447] br[447] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_448 bl[448] br[448] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_449 bl[449] br[449] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_450 bl[450] br[450] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_451 bl[451] br[451] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_452 bl[452] br[452] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_453 bl[453] br[453] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_454 bl[454] br[454] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_455 bl[455] br[455] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_456 bl[456] br[456] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_457 bl[457] br[457] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_458 bl[458] br[458] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_459 bl[459] br[459] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_460 bl[460] br[460] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_461 bl[461] br[461] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_462 bl[462] br[462] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_463 bl[463] br[463] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_464 bl[464] br[464] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_465 bl[465] br[465] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_466 bl[466] br[466] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_467 bl[467] br[467] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_468 bl[468] br[468] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_469 bl[469] br[469] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_470 bl[470] br[470] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_471 bl[471] br[471] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_472 bl[472] br[472] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_473 bl[473] br[473] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_474 bl[474] br[474] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_475 bl[475] br[475] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_476 bl[476] br[476] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_477 bl[477] br[477] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_478 bl[478] br[478] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_479 bl[479] br[479] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_480 bl[480] br[480] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_481 bl[481] br[481] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_482 bl[482] br[482] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_483 bl[483] br[483] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_484 bl[484] br[484] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_485 bl[485] br[485] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_486 bl[486] br[486] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_487 bl[487] br[487] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_488 bl[488] br[488] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_489 bl[489] br[489] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_490 bl[490] br[490] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_491 bl[491] br[491] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_492 bl[492] br[492] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_493 bl[493] br[493] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_494 bl[494] br[494] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_495 bl[495] br[495] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_496 bl[496] br[496] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_497 bl[497] br[497] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_498 bl[498] br[498] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_499 bl[499] br[499] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_500 bl[500] br[500] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_501 bl[501] br[501] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_502 bl[502] br[502] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_503 bl[503] br[503] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_504 bl[504] br[504] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_505 bl[505] br[505] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_506 bl[506] br[506] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_507 bl[507] br[507] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_508 bl[508] br[508] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_509 bl[509] br[509] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_510 bl[510] br[510] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_35_511 bl[511] br[511] vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xcell_36_0 bl[0] br[0] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_1 bl[1] br[1] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_2 bl[2] br[2] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_3 bl[3] br[3] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_4 bl[4] br[4] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_5 bl[5] br[5] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_6 bl[6] br[6] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_7 bl[7] br[7] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_8 bl[8] br[8] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_9 bl[9] br[9] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_10 bl[10] br[10] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_11 bl[11] br[11] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_12 bl[12] br[12] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_13 bl[13] br[13] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_14 bl[14] br[14] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_15 bl[15] br[15] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_16 bl[16] br[16] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_17 bl[17] br[17] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_18 bl[18] br[18] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_19 bl[19] br[19] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_20 bl[20] br[20] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_21 bl[21] br[21] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_22 bl[22] br[22] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_23 bl[23] br[23] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_24 bl[24] br[24] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_25 bl[25] br[25] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_26 bl[26] br[26] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_27 bl[27] br[27] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_28 bl[28] br[28] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_29 bl[29] br[29] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_30 bl[30] br[30] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_31 bl[31] br[31] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_32 bl[32] br[32] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_33 bl[33] br[33] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_34 bl[34] br[34] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_35 bl[35] br[35] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_36 bl[36] br[36] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_37 bl[37] br[37] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_38 bl[38] br[38] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_39 bl[39] br[39] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_40 bl[40] br[40] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_41 bl[41] br[41] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_42 bl[42] br[42] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_43 bl[43] br[43] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_44 bl[44] br[44] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_45 bl[45] br[45] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_46 bl[46] br[46] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_47 bl[47] br[47] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_48 bl[48] br[48] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_49 bl[49] br[49] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_50 bl[50] br[50] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_51 bl[51] br[51] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_52 bl[52] br[52] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_53 bl[53] br[53] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_54 bl[54] br[54] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_55 bl[55] br[55] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_56 bl[56] br[56] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_57 bl[57] br[57] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_58 bl[58] br[58] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_59 bl[59] br[59] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_60 bl[60] br[60] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_61 bl[61] br[61] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_62 bl[62] br[62] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_63 bl[63] br[63] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_64 bl[64] br[64] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_65 bl[65] br[65] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_66 bl[66] br[66] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_67 bl[67] br[67] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_68 bl[68] br[68] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_69 bl[69] br[69] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_70 bl[70] br[70] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_71 bl[71] br[71] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_72 bl[72] br[72] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_73 bl[73] br[73] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_74 bl[74] br[74] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_75 bl[75] br[75] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_76 bl[76] br[76] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_77 bl[77] br[77] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_78 bl[78] br[78] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_79 bl[79] br[79] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_80 bl[80] br[80] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_81 bl[81] br[81] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_82 bl[82] br[82] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_83 bl[83] br[83] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_84 bl[84] br[84] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_85 bl[85] br[85] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_86 bl[86] br[86] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_87 bl[87] br[87] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_88 bl[88] br[88] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_89 bl[89] br[89] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_90 bl[90] br[90] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_91 bl[91] br[91] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_92 bl[92] br[92] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_93 bl[93] br[93] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_94 bl[94] br[94] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_95 bl[95] br[95] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_96 bl[96] br[96] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_97 bl[97] br[97] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_98 bl[98] br[98] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_99 bl[99] br[99] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_100 bl[100] br[100] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_101 bl[101] br[101] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_102 bl[102] br[102] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_103 bl[103] br[103] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_104 bl[104] br[104] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_105 bl[105] br[105] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_106 bl[106] br[106] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_107 bl[107] br[107] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_108 bl[108] br[108] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_109 bl[109] br[109] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_110 bl[110] br[110] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_111 bl[111] br[111] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_112 bl[112] br[112] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_113 bl[113] br[113] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_114 bl[114] br[114] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_115 bl[115] br[115] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_116 bl[116] br[116] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_117 bl[117] br[117] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_118 bl[118] br[118] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_119 bl[119] br[119] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_120 bl[120] br[120] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_121 bl[121] br[121] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_122 bl[122] br[122] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_123 bl[123] br[123] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_124 bl[124] br[124] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_125 bl[125] br[125] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_126 bl[126] br[126] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_127 bl[127] br[127] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_128 bl[128] br[128] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_129 bl[129] br[129] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_130 bl[130] br[130] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_131 bl[131] br[131] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_132 bl[132] br[132] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_133 bl[133] br[133] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_134 bl[134] br[134] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_135 bl[135] br[135] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_136 bl[136] br[136] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_137 bl[137] br[137] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_138 bl[138] br[138] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_139 bl[139] br[139] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_140 bl[140] br[140] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_141 bl[141] br[141] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_142 bl[142] br[142] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_143 bl[143] br[143] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_144 bl[144] br[144] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_145 bl[145] br[145] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_146 bl[146] br[146] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_147 bl[147] br[147] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_148 bl[148] br[148] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_149 bl[149] br[149] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_150 bl[150] br[150] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_151 bl[151] br[151] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_152 bl[152] br[152] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_153 bl[153] br[153] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_154 bl[154] br[154] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_155 bl[155] br[155] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_156 bl[156] br[156] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_157 bl[157] br[157] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_158 bl[158] br[158] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_159 bl[159] br[159] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_160 bl[160] br[160] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_161 bl[161] br[161] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_162 bl[162] br[162] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_163 bl[163] br[163] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_164 bl[164] br[164] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_165 bl[165] br[165] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_166 bl[166] br[166] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_167 bl[167] br[167] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_168 bl[168] br[168] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_169 bl[169] br[169] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_170 bl[170] br[170] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_171 bl[171] br[171] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_172 bl[172] br[172] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_173 bl[173] br[173] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_174 bl[174] br[174] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_175 bl[175] br[175] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_176 bl[176] br[176] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_177 bl[177] br[177] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_178 bl[178] br[178] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_179 bl[179] br[179] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_180 bl[180] br[180] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_181 bl[181] br[181] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_182 bl[182] br[182] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_183 bl[183] br[183] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_184 bl[184] br[184] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_185 bl[185] br[185] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_186 bl[186] br[186] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_187 bl[187] br[187] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_188 bl[188] br[188] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_189 bl[189] br[189] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_190 bl[190] br[190] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_191 bl[191] br[191] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_192 bl[192] br[192] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_193 bl[193] br[193] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_194 bl[194] br[194] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_195 bl[195] br[195] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_196 bl[196] br[196] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_197 bl[197] br[197] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_198 bl[198] br[198] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_199 bl[199] br[199] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_200 bl[200] br[200] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_201 bl[201] br[201] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_202 bl[202] br[202] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_203 bl[203] br[203] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_204 bl[204] br[204] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_205 bl[205] br[205] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_206 bl[206] br[206] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_207 bl[207] br[207] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_208 bl[208] br[208] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_209 bl[209] br[209] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_210 bl[210] br[210] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_211 bl[211] br[211] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_212 bl[212] br[212] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_213 bl[213] br[213] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_214 bl[214] br[214] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_215 bl[215] br[215] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_216 bl[216] br[216] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_217 bl[217] br[217] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_218 bl[218] br[218] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_219 bl[219] br[219] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_220 bl[220] br[220] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_221 bl[221] br[221] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_222 bl[222] br[222] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_223 bl[223] br[223] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_224 bl[224] br[224] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_225 bl[225] br[225] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_226 bl[226] br[226] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_227 bl[227] br[227] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_228 bl[228] br[228] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_229 bl[229] br[229] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_230 bl[230] br[230] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_231 bl[231] br[231] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_232 bl[232] br[232] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_233 bl[233] br[233] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_234 bl[234] br[234] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_235 bl[235] br[235] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_236 bl[236] br[236] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_237 bl[237] br[237] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_238 bl[238] br[238] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_239 bl[239] br[239] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_240 bl[240] br[240] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_241 bl[241] br[241] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_242 bl[242] br[242] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_243 bl[243] br[243] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_244 bl[244] br[244] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_245 bl[245] br[245] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_246 bl[246] br[246] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_247 bl[247] br[247] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_248 bl[248] br[248] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_249 bl[249] br[249] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_250 bl[250] br[250] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_251 bl[251] br[251] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_252 bl[252] br[252] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_253 bl[253] br[253] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_254 bl[254] br[254] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_255 bl[255] br[255] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_256 bl[256] br[256] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_257 bl[257] br[257] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_258 bl[258] br[258] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_259 bl[259] br[259] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_260 bl[260] br[260] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_261 bl[261] br[261] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_262 bl[262] br[262] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_263 bl[263] br[263] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_264 bl[264] br[264] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_265 bl[265] br[265] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_266 bl[266] br[266] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_267 bl[267] br[267] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_268 bl[268] br[268] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_269 bl[269] br[269] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_270 bl[270] br[270] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_271 bl[271] br[271] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_272 bl[272] br[272] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_273 bl[273] br[273] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_274 bl[274] br[274] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_275 bl[275] br[275] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_276 bl[276] br[276] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_277 bl[277] br[277] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_278 bl[278] br[278] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_279 bl[279] br[279] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_280 bl[280] br[280] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_281 bl[281] br[281] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_282 bl[282] br[282] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_283 bl[283] br[283] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_284 bl[284] br[284] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_285 bl[285] br[285] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_286 bl[286] br[286] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_287 bl[287] br[287] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_288 bl[288] br[288] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_289 bl[289] br[289] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_290 bl[290] br[290] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_291 bl[291] br[291] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_292 bl[292] br[292] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_293 bl[293] br[293] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_294 bl[294] br[294] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_295 bl[295] br[295] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_296 bl[296] br[296] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_297 bl[297] br[297] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_298 bl[298] br[298] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_299 bl[299] br[299] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_300 bl[300] br[300] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_301 bl[301] br[301] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_302 bl[302] br[302] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_303 bl[303] br[303] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_304 bl[304] br[304] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_305 bl[305] br[305] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_306 bl[306] br[306] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_307 bl[307] br[307] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_308 bl[308] br[308] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_309 bl[309] br[309] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_310 bl[310] br[310] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_311 bl[311] br[311] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_312 bl[312] br[312] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_313 bl[313] br[313] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_314 bl[314] br[314] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_315 bl[315] br[315] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_316 bl[316] br[316] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_317 bl[317] br[317] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_318 bl[318] br[318] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_319 bl[319] br[319] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_320 bl[320] br[320] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_321 bl[321] br[321] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_322 bl[322] br[322] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_323 bl[323] br[323] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_324 bl[324] br[324] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_325 bl[325] br[325] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_326 bl[326] br[326] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_327 bl[327] br[327] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_328 bl[328] br[328] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_329 bl[329] br[329] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_330 bl[330] br[330] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_331 bl[331] br[331] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_332 bl[332] br[332] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_333 bl[333] br[333] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_334 bl[334] br[334] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_335 bl[335] br[335] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_336 bl[336] br[336] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_337 bl[337] br[337] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_338 bl[338] br[338] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_339 bl[339] br[339] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_340 bl[340] br[340] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_341 bl[341] br[341] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_342 bl[342] br[342] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_343 bl[343] br[343] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_344 bl[344] br[344] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_345 bl[345] br[345] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_346 bl[346] br[346] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_347 bl[347] br[347] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_348 bl[348] br[348] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_349 bl[349] br[349] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_350 bl[350] br[350] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_351 bl[351] br[351] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_352 bl[352] br[352] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_353 bl[353] br[353] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_354 bl[354] br[354] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_355 bl[355] br[355] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_356 bl[356] br[356] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_357 bl[357] br[357] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_358 bl[358] br[358] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_359 bl[359] br[359] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_360 bl[360] br[360] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_361 bl[361] br[361] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_362 bl[362] br[362] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_363 bl[363] br[363] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_364 bl[364] br[364] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_365 bl[365] br[365] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_366 bl[366] br[366] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_367 bl[367] br[367] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_368 bl[368] br[368] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_369 bl[369] br[369] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_370 bl[370] br[370] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_371 bl[371] br[371] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_372 bl[372] br[372] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_373 bl[373] br[373] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_374 bl[374] br[374] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_375 bl[375] br[375] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_376 bl[376] br[376] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_377 bl[377] br[377] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_378 bl[378] br[378] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_379 bl[379] br[379] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_380 bl[380] br[380] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_381 bl[381] br[381] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_382 bl[382] br[382] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_383 bl[383] br[383] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_384 bl[384] br[384] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_385 bl[385] br[385] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_386 bl[386] br[386] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_387 bl[387] br[387] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_388 bl[388] br[388] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_389 bl[389] br[389] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_390 bl[390] br[390] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_391 bl[391] br[391] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_392 bl[392] br[392] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_393 bl[393] br[393] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_394 bl[394] br[394] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_395 bl[395] br[395] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_396 bl[396] br[396] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_397 bl[397] br[397] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_398 bl[398] br[398] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_399 bl[399] br[399] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_400 bl[400] br[400] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_401 bl[401] br[401] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_402 bl[402] br[402] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_403 bl[403] br[403] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_404 bl[404] br[404] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_405 bl[405] br[405] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_406 bl[406] br[406] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_407 bl[407] br[407] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_408 bl[408] br[408] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_409 bl[409] br[409] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_410 bl[410] br[410] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_411 bl[411] br[411] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_412 bl[412] br[412] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_413 bl[413] br[413] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_414 bl[414] br[414] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_415 bl[415] br[415] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_416 bl[416] br[416] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_417 bl[417] br[417] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_418 bl[418] br[418] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_419 bl[419] br[419] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_420 bl[420] br[420] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_421 bl[421] br[421] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_422 bl[422] br[422] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_423 bl[423] br[423] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_424 bl[424] br[424] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_425 bl[425] br[425] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_426 bl[426] br[426] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_427 bl[427] br[427] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_428 bl[428] br[428] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_429 bl[429] br[429] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_430 bl[430] br[430] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_431 bl[431] br[431] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_432 bl[432] br[432] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_433 bl[433] br[433] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_434 bl[434] br[434] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_435 bl[435] br[435] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_436 bl[436] br[436] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_437 bl[437] br[437] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_438 bl[438] br[438] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_439 bl[439] br[439] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_440 bl[440] br[440] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_441 bl[441] br[441] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_442 bl[442] br[442] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_443 bl[443] br[443] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_444 bl[444] br[444] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_445 bl[445] br[445] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_446 bl[446] br[446] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_447 bl[447] br[447] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_448 bl[448] br[448] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_449 bl[449] br[449] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_450 bl[450] br[450] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_451 bl[451] br[451] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_452 bl[452] br[452] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_453 bl[453] br[453] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_454 bl[454] br[454] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_455 bl[455] br[455] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_456 bl[456] br[456] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_457 bl[457] br[457] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_458 bl[458] br[458] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_459 bl[459] br[459] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_460 bl[460] br[460] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_461 bl[461] br[461] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_462 bl[462] br[462] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_463 bl[463] br[463] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_464 bl[464] br[464] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_465 bl[465] br[465] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_466 bl[466] br[466] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_467 bl[467] br[467] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_468 bl[468] br[468] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_469 bl[469] br[469] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_470 bl[470] br[470] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_471 bl[471] br[471] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_472 bl[472] br[472] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_473 bl[473] br[473] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_474 bl[474] br[474] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_475 bl[475] br[475] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_476 bl[476] br[476] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_477 bl[477] br[477] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_478 bl[478] br[478] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_479 bl[479] br[479] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_480 bl[480] br[480] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_481 bl[481] br[481] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_482 bl[482] br[482] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_483 bl[483] br[483] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_484 bl[484] br[484] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_485 bl[485] br[485] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_486 bl[486] br[486] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_487 bl[487] br[487] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_488 bl[488] br[488] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_489 bl[489] br[489] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_490 bl[490] br[490] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_491 bl[491] br[491] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_492 bl[492] br[492] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_493 bl[493] br[493] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_494 bl[494] br[494] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_495 bl[495] br[495] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_496 bl[496] br[496] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_497 bl[497] br[497] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_498 bl[498] br[498] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_499 bl[499] br[499] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_500 bl[500] br[500] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_501 bl[501] br[501] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_502 bl[502] br[502] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_503 bl[503] br[503] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_504 bl[504] br[504] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_505 bl[505] br[505] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_506 bl[506] br[506] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_507 bl[507] br[507] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_508 bl[508] br[508] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_509 bl[509] br[509] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_510 bl[510] br[510] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_36_511 bl[511] br[511] vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xcell_37_0 bl[0] br[0] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_1 bl[1] br[1] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_2 bl[2] br[2] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_3 bl[3] br[3] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_4 bl[4] br[4] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_5 bl[5] br[5] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_6 bl[6] br[6] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_7 bl[7] br[7] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_8 bl[8] br[8] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_9 bl[9] br[9] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_10 bl[10] br[10] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_11 bl[11] br[11] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_12 bl[12] br[12] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_13 bl[13] br[13] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_14 bl[14] br[14] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_15 bl[15] br[15] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_16 bl[16] br[16] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_17 bl[17] br[17] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_18 bl[18] br[18] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_19 bl[19] br[19] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_20 bl[20] br[20] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_21 bl[21] br[21] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_22 bl[22] br[22] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_23 bl[23] br[23] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_24 bl[24] br[24] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_25 bl[25] br[25] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_26 bl[26] br[26] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_27 bl[27] br[27] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_28 bl[28] br[28] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_29 bl[29] br[29] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_30 bl[30] br[30] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_31 bl[31] br[31] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_32 bl[32] br[32] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_33 bl[33] br[33] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_34 bl[34] br[34] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_35 bl[35] br[35] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_36 bl[36] br[36] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_37 bl[37] br[37] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_38 bl[38] br[38] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_39 bl[39] br[39] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_40 bl[40] br[40] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_41 bl[41] br[41] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_42 bl[42] br[42] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_43 bl[43] br[43] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_44 bl[44] br[44] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_45 bl[45] br[45] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_46 bl[46] br[46] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_47 bl[47] br[47] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_48 bl[48] br[48] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_49 bl[49] br[49] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_50 bl[50] br[50] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_51 bl[51] br[51] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_52 bl[52] br[52] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_53 bl[53] br[53] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_54 bl[54] br[54] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_55 bl[55] br[55] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_56 bl[56] br[56] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_57 bl[57] br[57] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_58 bl[58] br[58] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_59 bl[59] br[59] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_60 bl[60] br[60] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_61 bl[61] br[61] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_62 bl[62] br[62] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_63 bl[63] br[63] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_64 bl[64] br[64] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_65 bl[65] br[65] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_66 bl[66] br[66] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_67 bl[67] br[67] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_68 bl[68] br[68] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_69 bl[69] br[69] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_70 bl[70] br[70] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_71 bl[71] br[71] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_72 bl[72] br[72] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_73 bl[73] br[73] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_74 bl[74] br[74] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_75 bl[75] br[75] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_76 bl[76] br[76] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_77 bl[77] br[77] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_78 bl[78] br[78] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_79 bl[79] br[79] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_80 bl[80] br[80] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_81 bl[81] br[81] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_82 bl[82] br[82] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_83 bl[83] br[83] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_84 bl[84] br[84] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_85 bl[85] br[85] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_86 bl[86] br[86] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_87 bl[87] br[87] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_88 bl[88] br[88] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_89 bl[89] br[89] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_90 bl[90] br[90] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_91 bl[91] br[91] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_92 bl[92] br[92] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_93 bl[93] br[93] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_94 bl[94] br[94] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_95 bl[95] br[95] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_96 bl[96] br[96] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_97 bl[97] br[97] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_98 bl[98] br[98] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_99 bl[99] br[99] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_100 bl[100] br[100] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_101 bl[101] br[101] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_102 bl[102] br[102] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_103 bl[103] br[103] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_104 bl[104] br[104] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_105 bl[105] br[105] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_106 bl[106] br[106] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_107 bl[107] br[107] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_108 bl[108] br[108] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_109 bl[109] br[109] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_110 bl[110] br[110] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_111 bl[111] br[111] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_112 bl[112] br[112] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_113 bl[113] br[113] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_114 bl[114] br[114] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_115 bl[115] br[115] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_116 bl[116] br[116] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_117 bl[117] br[117] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_118 bl[118] br[118] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_119 bl[119] br[119] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_120 bl[120] br[120] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_121 bl[121] br[121] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_122 bl[122] br[122] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_123 bl[123] br[123] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_124 bl[124] br[124] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_125 bl[125] br[125] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_126 bl[126] br[126] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_127 bl[127] br[127] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_128 bl[128] br[128] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_129 bl[129] br[129] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_130 bl[130] br[130] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_131 bl[131] br[131] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_132 bl[132] br[132] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_133 bl[133] br[133] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_134 bl[134] br[134] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_135 bl[135] br[135] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_136 bl[136] br[136] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_137 bl[137] br[137] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_138 bl[138] br[138] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_139 bl[139] br[139] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_140 bl[140] br[140] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_141 bl[141] br[141] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_142 bl[142] br[142] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_143 bl[143] br[143] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_144 bl[144] br[144] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_145 bl[145] br[145] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_146 bl[146] br[146] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_147 bl[147] br[147] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_148 bl[148] br[148] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_149 bl[149] br[149] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_150 bl[150] br[150] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_151 bl[151] br[151] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_152 bl[152] br[152] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_153 bl[153] br[153] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_154 bl[154] br[154] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_155 bl[155] br[155] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_156 bl[156] br[156] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_157 bl[157] br[157] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_158 bl[158] br[158] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_159 bl[159] br[159] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_160 bl[160] br[160] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_161 bl[161] br[161] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_162 bl[162] br[162] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_163 bl[163] br[163] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_164 bl[164] br[164] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_165 bl[165] br[165] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_166 bl[166] br[166] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_167 bl[167] br[167] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_168 bl[168] br[168] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_169 bl[169] br[169] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_170 bl[170] br[170] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_171 bl[171] br[171] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_172 bl[172] br[172] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_173 bl[173] br[173] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_174 bl[174] br[174] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_175 bl[175] br[175] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_176 bl[176] br[176] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_177 bl[177] br[177] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_178 bl[178] br[178] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_179 bl[179] br[179] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_180 bl[180] br[180] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_181 bl[181] br[181] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_182 bl[182] br[182] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_183 bl[183] br[183] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_184 bl[184] br[184] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_185 bl[185] br[185] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_186 bl[186] br[186] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_187 bl[187] br[187] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_188 bl[188] br[188] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_189 bl[189] br[189] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_190 bl[190] br[190] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_191 bl[191] br[191] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_192 bl[192] br[192] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_193 bl[193] br[193] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_194 bl[194] br[194] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_195 bl[195] br[195] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_196 bl[196] br[196] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_197 bl[197] br[197] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_198 bl[198] br[198] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_199 bl[199] br[199] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_200 bl[200] br[200] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_201 bl[201] br[201] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_202 bl[202] br[202] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_203 bl[203] br[203] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_204 bl[204] br[204] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_205 bl[205] br[205] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_206 bl[206] br[206] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_207 bl[207] br[207] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_208 bl[208] br[208] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_209 bl[209] br[209] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_210 bl[210] br[210] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_211 bl[211] br[211] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_212 bl[212] br[212] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_213 bl[213] br[213] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_214 bl[214] br[214] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_215 bl[215] br[215] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_216 bl[216] br[216] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_217 bl[217] br[217] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_218 bl[218] br[218] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_219 bl[219] br[219] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_220 bl[220] br[220] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_221 bl[221] br[221] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_222 bl[222] br[222] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_223 bl[223] br[223] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_224 bl[224] br[224] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_225 bl[225] br[225] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_226 bl[226] br[226] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_227 bl[227] br[227] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_228 bl[228] br[228] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_229 bl[229] br[229] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_230 bl[230] br[230] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_231 bl[231] br[231] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_232 bl[232] br[232] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_233 bl[233] br[233] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_234 bl[234] br[234] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_235 bl[235] br[235] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_236 bl[236] br[236] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_237 bl[237] br[237] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_238 bl[238] br[238] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_239 bl[239] br[239] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_240 bl[240] br[240] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_241 bl[241] br[241] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_242 bl[242] br[242] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_243 bl[243] br[243] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_244 bl[244] br[244] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_245 bl[245] br[245] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_246 bl[246] br[246] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_247 bl[247] br[247] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_248 bl[248] br[248] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_249 bl[249] br[249] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_250 bl[250] br[250] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_251 bl[251] br[251] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_252 bl[252] br[252] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_253 bl[253] br[253] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_254 bl[254] br[254] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_255 bl[255] br[255] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_256 bl[256] br[256] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_257 bl[257] br[257] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_258 bl[258] br[258] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_259 bl[259] br[259] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_260 bl[260] br[260] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_261 bl[261] br[261] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_262 bl[262] br[262] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_263 bl[263] br[263] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_264 bl[264] br[264] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_265 bl[265] br[265] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_266 bl[266] br[266] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_267 bl[267] br[267] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_268 bl[268] br[268] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_269 bl[269] br[269] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_270 bl[270] br[270] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_271 bl[271] br[271] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_272 bl[272] br[272] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_273 bl[273] br[273] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_274 bl[274] br[274] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_275 bl[275] br[275] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_276 bl[276] br[276] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_277 bl[277] br[277] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_278 bl[278] br[278] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_279 bl[279] br[279] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_280 bl[280] br[280] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_281 bl[281] br[281] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_282 bl[282] br[282] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_283 bl[283] br[283] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_284 bl[284] br[284] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_285 bl[285] br[285] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_286 bl[286] br[286] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_287 bl[287] br[287] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_288 bl[288] br[288] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_289 bl[289] br[289] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_290 bl[290] br[290] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_291 bl[291] br[291] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_292 bl[292] br[292] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_293 bl[293] br[293] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_294 bl[294] br[294] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_295 bl[295] br[295] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_296 bl[296] br[296] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_297 bl[297] br[297] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_298 bl[298] br[298] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_299 bl[299] br[299] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_300 bl[300] br[300] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_301 bl[301] br[301] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_302 bl[302] br[302] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_303 bl[303] br[303] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_304 bl[304] br[304] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_305 bl[305] br[305] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_306 bl[306] br[306] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_307 bl[307] br[307] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_308 bl[308] br[308] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_309 bl[309] br[309] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_310 bl[310] br[310] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_311 bl[311] br[311] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_312 bl[312] br[312] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_313 bl[313] br[313] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_314 bl[314] br[314] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_315 bl[315] br[315] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_316 bl[316] br[316] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_317 bl[317] br[317] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_318 bl[318] br[318] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_319 bl[319] br[319] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_320 bl[320] br[320] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_321 bl[321] br[321] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_322 bl[322] br[322] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_323 bl[323] br[323] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_324 bl[324] br[324] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_325 bl[325] br[325] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_326 bl[326] br[326] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_327 bl[327] br[327] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_328 bl[328] br[328] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_329 bl[329] br[329] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_330 bl[330] br[330] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_331 bl[331] br[331] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_332 bl[332] br[332] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_333 bl[333] br[333] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_334 bl[334] br[334] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_335 bl[335] br[335] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_336 bl[336] br[336] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_337 bl[337] br[337] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_338 bl[338] br[338] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_339 bl[339] br[339] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_340 bl[340] br[340] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_341 bl[341] br[341] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_342 bl[342] br[342] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_343 bl[343] br[343] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_344 bl[344] br[344] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_345 bl[345] br[345] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_346 bl[346] br[346] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_347 bl[347] br[347] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_348 bl[348] br[348] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_349 bl[349] br[349] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_350 bl[350] br[350] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_351 bl[351] br[351] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_352 bl[352] br[352] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_353 bl[353] br[353] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_354 bl[354] br[354] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_355 bl[355] br[355] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_356 bl[356] br[356] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_357 bl[357] br[357] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_358 bl[358] br[358] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_359 bl[359] br[359] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_360 bl[360] br[360] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_361 bl[361] br[361] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_362 bl[362] br[362] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_363 bl[363] br[363] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_364 bl[364] br[364] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_365 bl[365] br[365] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_366 bl[366] br[366] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_367 bl[367] br[367] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_368 bl[368] br[368] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_369 bl[369] br[369] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_370 bl[370] br[370] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_371 bl[371] br[371] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_372 bl[372] br[372] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_373 bl[373] br[373] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_374 bl[374] br[374] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_375 bl[375] br[375] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_376 bl[376] br[376] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_377 bl[377] br[377] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_378 bl[378] br[378] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_379 bl[379] br[379] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_380 bl[380] br[380] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_381 bl[381] br[381] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_382 bl[382] br[382] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_383 bl[383] br[383] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_384 bl[384] br[384] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_385 bl[385] br[385] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_386 bl[386] br[386] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_387 bl[387] br[387] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_388 bl[388] br[388] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_389 bl[389] br[389] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_390 bl[390] br[390] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_391 bl[391] br[391] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_392 bl[392] br[392] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_393 bl[393] br[393] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_394 bl[394] br[394] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_395 bl[395] br[395] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_396 bl[396] br[396] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_397 bl[397] br[397] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_398 bl[398] br[398] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_399 bl[399] br[399] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_400 bl[400] br[400] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_401 bl[401] br[401] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_402 bl[402] br[402] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_403 bl[403] br[403] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_404 bl[404] br[404] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_405 bl[405] br[405] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_406 bl[406] br[406] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_407 bl[407] br[407] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_408 bl[408] br[408] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_409 bl[409] br[409] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_410 bl[410] br[410] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_411 bl[411] br[411] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_412 bl[412] br[412] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_413 bl[413] br[413] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_414 bl[414] br[414] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_415 bl[415] br[415] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_416 bl[416] br[416] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_417 bl[417] br[417] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_418 bl[418] br[418] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_419 bl[419] br[419] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_420 bl[420] br[420] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_421 bl[421] br[421] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_422 bl[422] br[422] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_423 bl[423] br[423] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_424 bl[424] br[424] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_425 bl[425] br[425] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_426 bl[426] br[426] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_427 bl[427] br[427] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_428 bl[428] br[428] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_429 bl[429] br[429] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_430 bl[430] br[430] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_431 bl[431] br[431] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_432 bl[432] br[432] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_433 bl[433] br[433] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_434 bl[434] br[434] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_435 bl[435] br[435] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_436 bl[436] br[436] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_437 bl[437] br[437] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_438 bl[438] br[438] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_439 bl[439] br[439] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_440 bl[440] br[440] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_441 bl[441] br[441] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_442 bl[442] br[442] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_443 bl[443] br[443] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_444 bl[444] br[444] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_445 bl[445] br[445] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_446 bl[446] br[446] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_447 bl[447] br[447] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_448 bl[448] br[448] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_449 bl[449] br[449] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_450 bl[450] br[450] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_451 bl[451] br[451] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_452 bl[452] br[452] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_453 bl[453] br[453] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_454 bl[454] br[454] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_455 bl[455] br[455] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_456 bl[456] br[456] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_457 bl[457] br[457] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_458 bl[458] br[458] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_459 bl[459] br[459] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_460 bl[460] br[460] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_461 bl[461] br[461] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_462 bl[462] br[462] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_463 bl[463] br[463] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_464 bl[464] br[464] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_465 bl[465] br[465] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_466 bl[466] br[466] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_467 bl[467] br[467] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_468 bl[468] br[468] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_469 bl[469] br[469] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_470 bl[470] br[470] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_471 bl[471] br[471] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_472 bl[472] br[472] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_473 bl[473] br[473] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_474 bl[474] br[474] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_475 bl[475] br[475] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_476 bl[476] br[476] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_477 bl[477] br[477] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_478 bl[478] br[478] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_479 bl[479] br[479] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_480 bl[480] br[480] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_481 bl[481] br[481] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_482 bl[482] br[482] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_483 bl[483] br[483] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_484 bl[484] br[484] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_485 bl[485] br[485] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_486 bl[486] br[486] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_487 bl[487] br[487] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_488 bl[488] br[488] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_489 bl[489] br[489] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_490 bl[490] br[490] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_491 bl[491] br[491] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_492 bl[492] br[492] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_493 bl[493] br[493] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_494 bl[494] br[494] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_495 bl[495] br[495] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_496 bl[496] br[496] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_497 bl[497] br[497] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_498 bl[498] br[498] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_499 bl[499] br[499] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_500 bl[500] br[500] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_501 bl[501] br[501] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_502 bl[502] br[502] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_503 bl[503] br[503] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_504 bl[504] br[504] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_505 bl[505] br[505] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_506 bl[506] br[506] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_507 bl[507] br[507] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_508 bl[508] br[508] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_509 bl[509] br[509] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_510 bl[510] br[510] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_37_511 bl[511] br[511] vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xcell_38_0 bl[0] br[0] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_1 bl[1] br[1] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_2 bl[2] br[2] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_3 bl[3] br[3] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_4 bl[4] br[4] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_5 bl[5] br[5] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_6 bl[6] br[6] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_7 bl[7] br[7] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_8 bl[8] br[8] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_9 bl[9] br[9] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_10 bl[10] br[10] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_11 bl[11] br[11] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_12 bl[12] br[12] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_13 bl[13] br[13] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_14 bl[14] br[14] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_15 bl[15] br[15] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_16 bl[16] br[16] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_17 bl[17] br[17] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_18 bl[18] br[18] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_19 bl[19] br[19] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_20 bl[20] br[20] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_21 bl[21] br[21] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_22 bl[22] br[22] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_23 bl[23] br[23] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_24 bl[24] br[24] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_25 bl[25] br[25] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_26 bl[26] br[26] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_27 bl[27] br[27] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_28 bl[28] br[28] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_29 bl[29] br[29] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_30 bl[30] br[30] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_31 bl[31] br[31] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_32 bl[32] br[32] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_33 bl[33] br[33] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_34 bl[34] br[34] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_35 bl[35] br[35] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_36 bl[36] br[36] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_37 bl[37] br[37] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_38 bl[38] br[38] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_39 bl[39] br[39] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_40 bl[40] br[40] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_41 bl[41] br[41] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_42 bl[42] br[42] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_43 bl[43] br[43] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_44 bl[44] br[44] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_45 bl[45] br[45] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_46 bl[46] br[46] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_47 bl[47] br[47] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_48 bl[48] br[48] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_49 bl[49] br[49] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_50 bl[50] br[50] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_51 bl[51] br[51] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_52 bl[52] br[52] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_53 bl[53] br[53] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_54 bl[54] br[54] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_55 bl[55] br[55] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_56 bl[56] br[56] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_57 bl[57] br[57] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_58 bl[58] br[58] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_59 bl[59] br[59] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_60 bl[60] br[60] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_61 bl[61] br[61] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_62 bl[62] br[62] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_63 bl[63] br[63] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_64 bl[64] br[64] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_65 bl[65] br[65] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_66 bl[66] br[66] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_67 bl[67] br[67] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_68 bl[68] br[68] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_69 bl[69] br[69] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_70 bl[70] br[70] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_71 bl[71] br[71] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_72 bl[72] br[72] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_73 bl[73] br[73] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_74 bl[74] br[74] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_75 bl[75] br[75] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_76 bl[76] br[76] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_77 bl[77] br[77] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_78 bl[78] br[78] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_79 bl[79] br[79] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_80 bl[80] br[80] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_81 bl[81] br[81] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_82 bl[82] br[82] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_83 bl[83] br[83] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_84 bl[84] br[84] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_85 bl[85] br[85] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_86 bl[86] br[86] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_87 bl[87] br[87] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_88 bl[88] br[88] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_89 bl[89] br[89] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_90 bl[90] br[90] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_91 bl[91] br[91] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_92 bl[92] br[92] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_93 bl[93] br[93] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_94 bl[94] br[94] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_95 bl[95] br[95] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_96 bl[96] br[96] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_97 bl[97] br[97] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_98 bl[98] br[98] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_99 bl[99] br[99] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_100 bl[100] br[100] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_101 bl[101] br[101] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_102 bl[102] br[102] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_103 bl[103] br[103] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_104 bl[104] br[104] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_105 bl[105] br[105] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_106 bl[106] br[106] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_107 bl[107] br[107] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_108 bl[108] br[108] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_109 bl[109] br[109] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_110 bl[110] br[110] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_111 bl[111] br[111] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_112 bl[112] br[112] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_113 bl[113] br[113] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_114 bl[114] br[114] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_115 bl[115] br[115] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_116 bl[116] br[116] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_117 bl[117] br[117] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_118 bl[118] br[118] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_119 bl[119] br[119] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_120 bl[120] br[120] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_121 bl[121] br[121] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_122 bl[122] br[122] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_123 bl[123] br[123] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_124 bl[124] br[124] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_125 bl[125] br[125] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_126 bl[126] br[126] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_127 bl[127] br[127] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_128 bl[128] br[128] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_129 bl[129] br[129] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_130 bl[130] br[130] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_131 bl[131] br[131] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_132 bl[132] br[132] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_133 bl[133] br[133] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_134 bl[134] br[134] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_135 bl[135] br[135] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_136 bl[136] br[136] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_137 bl[137] br[137] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_138 bl[138] br[138] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_139 bl[139] br[139] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_140 bl[140] br[140] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_141 bl[141] br[141] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_142 bl[142] br[142] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_143 bl[143] br[143] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_144 bl[144] br[144] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_145 bl[145] br[145] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_146 bl[146] br[146] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_147 bl[147] br[147] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_148 bl[148] br[148] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_149 bl[149] br[149] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_150 bl[150] br[150] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_151 bl[151] br[151] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_152 bl[152] br[152] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_153 bl[153] br[153] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_154 bl[154] br[154] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_155 bl[155] br[155] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_156 bl[156] br[156] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_157 bl[157] br[157] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_158 bl[158] br[158] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_159 bl[159] br[159] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_160 bl[160] br[160] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_161 bl[161] br[161] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_162 bl[162] br[162] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_163 bl[163] br[163] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_164 bl[164] br[164] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_165 bl[165] br[165] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_166 bl[166] br[166] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_167 bl[167] br[167] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_168 bl[168] br[168] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_169 bl[169] br[169] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_170 bl[170] br[170] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_171 bl[171] br[171] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_172 bl[172] br[172] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_173 bl[173] br[173] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_174 bl[174] br[174] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_175 bl[175] br[175] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_176 bl[176] br[176] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_177 bl[177] br[177] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_178 bl[178] br[178] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_179 bl[179] br[179] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_180 bl[180] br[180] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_181 bl[181] br[181] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_182 bl[182] br[182] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_183 bl[183] br[183] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_184 bl[184] br[184] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_185 bl[185] br[185] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_186 bl[186] br[186] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_187 bl[187] br[187] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_188 bl[188] br[188] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_189 bl[189] br[189] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_190 bl[190] br[190] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_191 bl[191] br[191] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_192 bl[192] br[192] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_193 bl[193] br[193] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_194 bl[194] br[194] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_195 bl[195] br[195] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_196 bl[196] br[196] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_197 bl[197] br[197] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_198 bl[198] br[198] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_199 bl[199] br[199] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_200 bl[200] br[200] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_201 bl[201] br[201] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_202 bl[202] br[202] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_203 bl[203] br[203] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_204 bl[204] br[204] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_205 bl[205] br[205] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_206 bl[206] br[206] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_207 bl[207] br[207] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_208 bl[208] br[208] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_209 bl[209] br[209] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_210 bl[210] br[210] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_211 bl[211] br[211] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_212 bl[212] br[212] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_213 bl[213] br[213] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_214 bl[214] br[214] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_215 bl[215] br[215] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_216 bl[216] br[216] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_217 bl[217] br[217] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_218 bl[218] br[218] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_219 bl[219] br[219] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_220 bl[220] br[220] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_221 bl[221] br[221] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_222 bl[222] br[222] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_223 bl[223] br[223] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_224 bl[224] br[224] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_225 bl[225] br[225] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_226 bl[226] br[226] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_227 bl[227] br[227] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_228 bl[228] br[228] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_229 bl[229] br[229] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_230 bl[230] br[230] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_231 bl[231] br[231] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_232 bl[232] br[232] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_233 bl[233] br[233] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_234 bl[234] br[234] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_235 bl[235] br[235] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_236 bl[236] br[236] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_237 bl[237] br[237] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_238 bl[238] br[238] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_239 bl[239] br[239] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_240 bl[240] br[240] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_241 bl[241] br[241] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_242 bl[242] br[242] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_243 bl[243] br[243] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_244 bl[244] br[244] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_245 bl[245] br[245] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_246 bl[246] br[246] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_247 bl[247] br[247] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_248 bl[248] br[248] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_249 bl[249] br[249] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_250 bl[250] br[250] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_251 bl[251] br[251] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_252 bl[252] br[252] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_253 bl[253] br[253] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_254 bl[254] br[254] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_255 bl[255] br[255] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_256 bl[256] br[256] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_257 bl[257] br[257] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_258 bl[258] br[258] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_259 bl[259] br[259] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_260 bl[260] br[260] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_261 bl[261] br[261] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_262 bl[262] br[262] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_263 bl[263] br[263] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_264 bl[264] br[264] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_265 bl[265] br[265] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_266 bl[266] br[266] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_267 bl[267] br[267] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_268 bl[268] br[268] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_269 bl[269] br[269] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_270 bl[270] br[270] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_271 bl[271] br[271] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_272 bl[272] br[272] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_273 bl[273] br[273] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_274 bl[274] br[274] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_275 bl[275] br[275] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_276 bl[276] br[276] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_277 bl[277] br[277] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_278 bl[278] br[278] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_279 bl[279] br[279] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_280 bl[280] br[280] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_281 bl[281] br[281] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_282 bl[282] br[282] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_283 bl[283] br[283] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_284 bl[284] br[284] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_285 bl[285] br[285] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_286 bl[286] br[286] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_287 bl[287] br[287] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_288 bl[288] br[288] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_289 bl[289] br[289] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_290 bl[290] br[290] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_291 bl[291] br[291] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_292 bl[292] br[292] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_293 bl[293] br[293] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_294 bl[294] br[294] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_295 bl[295] br[295] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_296 bl[296] br[296] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_297 bl[297] br[297] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_298 bl[298] br[298] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_299 bl[299] br[299] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_300 bl[300] br[300] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_301 bl[301] br[301] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_302 bl[302] br[302] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_303 bl[303] br[303] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_304 bl[304] br[304] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_305 bl[305] br[305] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_306 bl[306] br[306] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_307 bl[307] br[307] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_308 bl[308] br[308] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_309 bl[309] br[309] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_310 bl[310] br[310] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_311 bl[311] br[311] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_312 bl[312] br[312] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_313 bl[313] br[313] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_314 bl[314] br[314] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_315 bl[315] br[315] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_316 bl[316] br[316] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_317 bl[317] br[317] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_318 bl[318] br[318] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_319 bl[319] br[319] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_320 bl[320] br[320] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_321 bl[321] br[321] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_322 bl[322] br[322] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_323 bl[323] br[323] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_324 bl[324] br[324] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_325 bl[325] br[325] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_326 bl[326] br[326] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_327 bl[327] br[327] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_328 bl[328] br[328] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_329 bl[329] br[329] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_330 bl[330] br[330] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_331 bl[331] br[331] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_332 bl[332] br[332] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_333 bl[333] br[333] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_334 bl[334] br[334] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_335 bl[335] br[335] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_336 bl[336] br[336] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_337 bl[337] br[337] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_338 bl[338] br[338] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_339 bl[339] br[339] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_340 bl[340] br[340] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_341 bl[341] br[341] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_342 bl[342] br[342] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_343 bl[343] br[343] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_344 bl[344] br[344] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_345 bl[345] br[345] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_346 bl[346] br[346] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_347 bl[347] br[347] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_348 bl[348] br[348] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_349 bl[349] br[349] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_350 bl[350] br[350] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_351 bl[351] br[351] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_352 bl[352] br[352] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_353 bl[353] br[353] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_354 bl[354] br[354] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_355 bl[355] br[355] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_356 bl[356] br[356] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_357 bl[357] br[357] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_358 bl[358] br[358] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_359 bl[359] br[359] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_360 bl[360] br[360] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_361 bl[361] br[361] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_362 bl[362] br[362] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_363 bl[363] br[363] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_364 bl[364] br[364] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_365 bl[365] br[365] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_366 bl[366] br[366] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_367 bl[367] br[367] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_368 bl[368] br[368] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_369 bl[369] br[369] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_370 bl[370] br[370] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_371 bl[371] br[371] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_372 bl[372] br[372] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_373 bl[373] br[373] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_374 bl[374] br[374] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_375 bl[375] br[375] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_376 bl[376] br[376] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_377 bl[377] br[377] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_378 bl[378] br[378] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_379 bl[379] br[379] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_380 bl[380] br[380] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_381 bl[381] br[381] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_382 bl[382] br[382] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_383 bl[383] br[383] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_384 bl[384] br[384] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_385 bl[385] br[385] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_386 bl[386] br[386] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_387 bl[387] br[387] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_388 bl[388] br[388] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_389 bl[389] br[389] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_390 bl[390] br[390] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_391 bl[391] br[391] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_392 bl[392] br[392] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_393 bl[393] br[393] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_394 bl[394] br[394] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_395 bl[395] br[395] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_396 bl[396] br[396] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_397 bl[397] br[397] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_398 bl[398] br[398] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_399 bl[399] br[399] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_400 bl[400] br[400] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_401 bl[401] br[401] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_402 bl[402] br[402] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_403 bl[403] br[403] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_404 bl[404] br[404] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_405 bl[405] br[405] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_406 bl[406] br[406] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_407 bl[407] br[407] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_408 bl[408] br[408] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_409 bl[409] br[409] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_410 bl[410] br[410] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_411 bl[411] br[411] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_412 bl[412] br[412] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_413 bl[413] br[413] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_414 bl[414] br[414] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_415 bl[415] br[415] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_416 bl[416] br[416] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_417 bl[417] br[417] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_418 bl[418] br[418] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_419 bl[419] br[419] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_420 bl[420] br[420] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_421 bl[421] br[421] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_422 bl[422] br[422] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_423 bl[423] br[423] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_424 bl[424] br[424] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_425 bl[425] br[425] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_426 bl[426] br[426] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_427 bl[427] br[427] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_428 bl[428] br[428] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_429 bl[429] br[429] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_430 bl[430] br[430] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_431 bl[431] br[431] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_432 bl[432] br[432] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_433 bl[433] br[433] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_434 bl[434] br[434] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_435 bl[435] br[435] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_436 bl[436] br[436] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_437 bl[437] br[437] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_438 bl[438] br[438] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_439 bl[439] br[439] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_440 bl[440] br[440] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_441 bl[441] br[441] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_442 bl[442] br[442] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_443 bl[443] br[443] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_444 bl[444] br[444] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_445 bl[445] br[445] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_446 bl[446] br[446] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_447 bl[447] br[447] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_448 bl[448] br[448] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_449 bl[449] br[449] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_450 bl[450] br[450] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_451 bl[451] br[451] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_452 bl[452] br[452] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_453 bl[453] br[453] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_454 bl[454] br[454] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_455 bl[455] br[455] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_456 bl[456] br[456] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_457 bl[457] br[457] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_458 bl[458] br[458] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_459 bl[459] br[459] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_460 bl[460] br[460] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_461 bl[461] br[461] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_462 bl[462] br[462] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_463 bl[463] br[463] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_464 bl[464] br[464] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_465 bl[465] br[465] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_466 bl[466] br[466] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_467 bl[467] br[467] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_468 bl[468] br[468] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_469 bl[469] br[469] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_470 bl[470] br[470] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_471 bl[471] br[471] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_472 bl[472] br[472] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_473 bl[473] br[473] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_474 bl[474] br[474] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_475 bl[475] br[475] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_476 bl[476] br[476] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_477 bl[477] br[477] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_478 bl[478] br[478] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_479 bl[479] br[479] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_480 bl[480] br[480] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_481 bl[481] br[481] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_482 bl[482] br[482] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_483 bl[483] br[483] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_484 bl[484] br[484] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_485 bl[485] br[485] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_486 bl[486] br[486] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_487 bl[487] br[487] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_488 bl[488] br[488] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_489 bl[489] br[489] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_490 bl[490] br[490] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_491 bl[491] br[491] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_492 bl[492] br[492] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_493 bl[493] br[493] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_494 bl[494] br[494] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_495 bl[495] br[495] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_496 bl[496] br[496] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_497 bl[497] br[497] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_498 bl[498] br[498] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_499 bl[499] br[499] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_500 bl[500] br[500] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_501 bl[501] br[501] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_502 bl[502] br[502] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_503 bl[503] br[503] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_504 bl[504] br[504] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_505 bl[505] br[505] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_506 bl[506] br[506] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_507 bl[507] br[507] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_508 bl[508] br[508] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_509 bl[509] br[509] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_510 bl[510] br[510] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_38_511 bl[511] br[511] vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xcell_39_0 bl[0] br[0] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_1 bl[1] br[1] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_2 bl[2] br[2] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_3 bl[3] br[3] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_4 bl[4] br[4] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_5 bl[5] br[5] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_6 bl[6] br[6] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_7 bl[7] br[7] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_8 bl[8] br[8] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_9 bl[9] br[9] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_10 bl[10] br[10] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_11 bl[11] br[11] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_12 bl[12] br[12] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_13 bl[13] br[13] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_14 bl[14] br[14] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_15 bl[15] br[15] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_16 bl[16] br[16] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_17 bl[17] br[17] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_18 bl[18] br[18] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_19 bl[19] br[19] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_20 bl[20] br[20] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_21 bl[21] br[21] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_22 bl[22] br[22] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_23 bl[23] br[23] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_24 bl[24] br[24] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_25 bl[25] br[25] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_26 bl[26] br[26] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_27 bl[27] br[27] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_28 bl[28] br[28] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_29 bl[29] br[29] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_30 bl[30] br[30] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_31 bl[31] br[31] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_32 bl[32] br[32] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_33 bl[33] br[33] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_34 bl[34] br[34] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_35 bl[35] br[35] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_36 bl[36] br[36] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_37 bl[37] br[37] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_38 bl[38] br[38] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_39 bl[39] br[39] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_40 bl[40] br[40] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_41 bl[41] br[41] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_42 bl[42] br[42] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_43 bl[43] br[43] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_44 bl[44] br[44] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_45 bl[45] br[45] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_46 bl[46] br[46] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_47 bl[47] br[47] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_48 bl[48] br[48] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_49 bl[49] br[49] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_50 bl[50] br[50] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_51 bl[51] br[51] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_52 bl[52] br[52] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_53 bl[53] br[53] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_54 bl[54] br[54] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_55 bl[55] br[55] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_56 bl[56] br[56] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_57 bl[57] br[57] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_58 bl[58] br[58] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_59 bl[59] br[59] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_60 bl[60] br[60] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_61 bl[61] br[61] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_62 bl[62] br[62] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_63 bl[63] br[63] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_64 bl[64] br[64] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_65 bl[65] br[65] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_66 bl[66] br[66] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_67 bl[67] br[67] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_68 bl[68] br[68] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_69 bl[69] br[69] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_70 bl[70] br[70] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_71 bl[71] br[71] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_72 bl[72] br[72] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_73 bl[73] br[73] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_74 bl[74] br[74] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_75 bl[75] br[75] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_76 bl[76] br[76] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_77 bl[77] br[77] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_78 bl[78] br[78] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_79 bl[79] br[79] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_80 bl[80] br[80] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_81 bl[81] br[81] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_82 bl[82] br[82] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_83 bl[83] br[83] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_84 bl[84] br[84] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_85 bl[85] br[85] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_86 bl[86] br[86] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_87 bl[87] br[87] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_88 bl[88] br[88] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_89 bl[89] br[89] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_90 bl[90] br[90] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_91 bl[91] br[91] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_92 bl[92] br[92] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_93 bl[93] br[93] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_94 bl[94] br[94] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_95 bl[95] br[95] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_96 bl[96] br[96] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_97 bl[97] br[97] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_98 bl[98] br[98] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_99 bl[99] br[99] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_100 bl[100] br[100] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_101 bl[101] br[101] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_102 bl[102] br[102] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_103 bl[103] br[103] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_104 bl[104] br[104] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_105 bl[105] br[105] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_106 bl[106] br[106] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_107 bl[107] br[107] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_108 bl[108] br[108] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_109 bl[109] br[109] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_110 bl[110] br[110] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_111 bl[111] br[111] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_112 bl[112] br[112] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_113 bl[113] br[113] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_114 bl[114] br[114] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_115 bl[115] br[115] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_116 bl[116] br[116] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_117 bl[117] br[117] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_118 bl[118] br[118] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_119 bl[119] br[119] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_120 bl[120] br[120] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_121 bl[121] br[121] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_122 bl[122] br[122] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_123 bl[123] br[123] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_124 bl[124] br[124] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_125 bl[125] br[125] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_126 bl[126] br[126] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_127 bl[127] br[127] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_128 bl[128] br[128] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_129 bl[129] br[129] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_130 bl[130] br[130] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_131 bl[131] br[131] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_132 bl[132] br[132] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_133 bl[133] br[133] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_134 bl[134] br[134] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_135 bl[135] br[135] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_136 bl[136] br[136] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_137 bl[137] br[137] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_138 bl[138] br[138] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_139 bl[139] br[139] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_140 bl[140] br[140] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_141 bl[141] br[141] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_142 bl[142] br[142] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_143 bl[143] br[143] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_144 bl[144] br[144] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_145 bl[145] br[145] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_146 bl[146] br[146] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_147 bl[147] br[147] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_148 bl[148] br[148] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_149 bl[149] br[149] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_150 bl[150] br[150] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_151 bl[151] br[151] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_152 bl[152] br[152] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_153 bl[153] br[153] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_154 bl[154] br[154] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_155 bl[155] br[155] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_156 bl[156] br[156] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_157 bl[157] br[157] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_158 bl[158] br[158] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_159 bl[159] br[159] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_160 bl[160] br[160] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_161 bl[161] br[161] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_162 bl[162] br[162] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_163 bl[163] br[163] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_164 bl[164] br[164] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_165 bl[165] br[165] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_166 bl[166] br[166] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_167 bl[167] br[167] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_168 bl[168] br[168] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_169 bl[169] br[169] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_170 bl[170] br[170] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_171 bl[171] br[171] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_172 bl[172] br[172] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_173 bl[173] br[173] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_174 bl[174] br[174] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_175 bl[175] br[175] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_176 bl[176] br[176] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_177 bl[177] br[177] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_178 bl[178] br[178] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_179 bl[179] br[179] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_180 bl[180] br[180] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_181 bl[181] br[181] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_182 bl[182] br[182] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_183 bl[183] br[183] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_184 bl[184] br[184] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_185 bl[185] br[185] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_186 bl[186] br[186] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_187 bl[187] br[187] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_188 bl[188] br[188] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_189 bl[189] br[189] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_190 bl[190] br[190] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_191 bl[191] br[191] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_192 bl[192] br[192] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_193 bl[193] br[193] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_194 bl[194] br[194] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_195 bl[195] br[195] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_196 bl[196] br[196] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_197 bl[197] br[197] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_198 bl[198] br[198] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_199 bl[199] br[199] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_200 bl[200] br[200] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_201 bl[201] br[201] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_202 bl[202] br[202] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_203 bl[203] br[203] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_204 bl[204] br[204] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_205 bl[205] br[205] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_206 bl[206] br[206] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_207 bl[207] br[207] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_208 bl[208] br[208] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_209 bl[209] br[209] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_210 bl[210] br[210] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_211 bl[211] br[211] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_212 bl[212] br[212] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_213 bl[213] br[213] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_214 bl[214] br[214] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_215 bl[215] br[215] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_216 bl[216] br[216] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_217 bl[217] br[217] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_218 bl[218] br[218] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_219 bl[219] br[219] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_220 bl[220] br[220] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_221 bl[221] br[221] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_222 bl[222] br[222] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_223 bl[223] br[223] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_224 bl[224] br[224] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_225 bl[225] br[225] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_226 bl[226] br[226] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_227 bl[227] br[227] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_228 bl[228] br[228] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_229 bl[229] br[229] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_230 bl[230] br[230] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_231 bl[231] br[231] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_232 bl[232] br[232] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_233 bl[233] br[233] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_234 bl[234] br[234] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_235 bl[235] br[235] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_236 bl[236] br[236] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_237 bl[237] br[237] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_238 bl[238] br[238] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_239 bl[239] br[239] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_240 bl[240] br[240] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_241 bl[241] br[241] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_242 bl[242] br[242] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_243 bl[243] br[243] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_244 bl[244] br[244] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_245 bl[245] br[245] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_246 bl[246] br[246] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_247 bl[247] br[247] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_248 bl[248] br[248] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_249 bl[249] br[249] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_250 bl[250] br[250] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_251 bl[251] br[251] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_252 bl[252] br[252] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_253 bl[253] br[253] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_254 bl[254] br[254] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_255 bl[255] br[255] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_256 bl[256] br[256] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_257 bl[257] br[257] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_258 bl[258] br[258] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_259 bl[259] br[259] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_260 bl[260] br[260] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_261 bl[261] br[261] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_262 bl[262] br[262] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_263 bl[263] br[263] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_264 bl[264] br[264] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_265 bl[265] br[265] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_266 bl[266] br[266] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_267 bl[267] br[267] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_268 bl[268] br[268] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_269 bl[269] br[269] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_270 bl[270] br[270] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_271 bl[271] br[271] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_272 bl[272] br[272] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_273 bl[273] br[273] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_274 bl[274] br[274] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_275 bl[275] br[275] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_276 bl[276] br[276] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_277 bl[277] br[277] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_278 bl[278] br[278] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_279 bl[279] br[279] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_280 bl[280] br[280] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_281 bl[281] br[281] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_282 bl[282] br[282] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_283 bl[283] br[283] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_284 bl[284] br[284] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_285 bl[285] br[285] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_286 bl[286] br[286] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_287 bl[287] br[287] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_288 bl[288] br[288] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_289 bl[289] br[289] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_290 bl[290] br[290] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_291 bl[291] br[291] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_292 bl[292] br[292] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_293 bl[293] br[293] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_294 bl[294] br[294] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_295 bl[295] br[295] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_296 bl[296] br[296] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_297 bl[297] br[297] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_298 bl[298] br[298] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_299 bl[299] br[299] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_300 bl[300] br[300] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_301 bl[301] br[301] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_302 bl[302] br[302] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_303 bl[303] br[303] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_304 bl[304] br[304] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_305 bl[305] br[305] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_306 bl[306] br[306] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_307 bl[307] br[307] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_308 bl[308] br[308] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_309 bl[309] br[309] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_310 bl[310] br[310] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_311 bl[311] br[311] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_312 bl[312] br[312] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_313 bl[313] br[313] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_314 bl[314] br[314] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_315 bl[315] br[315] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_316 bl[316] br[316] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_317 bl[317] br[317] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_318 bl[318] br[318] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_319 bl[319] br[319] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_320 bl[320] br[320] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_321 bl[321] br[321] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_322 bl[322] br[322] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_323 bl[323] br[323] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_324 bl[324] br[324] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_325 bl[325] br[325] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_326 bl[326] br[326] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_327 bl[327] br[327] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_328 bl[328] br[328] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_329 bl[329] br[329] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_330 bl[330] br[330] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_331 bl[331] br[331] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_332 bl[332] br[332] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_333 bl[333] br[333] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_334 bl[334] br[334] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_335 bl[335] br[335] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_336 bl[336] br[336] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_337 bl[337] br[337] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_338 bl[338] br[338] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_339 bl[339] br[339] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_340 bl[340] br[340] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_341 bl[341] br[341] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_342 bl[342] br[342] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_343 bl[343] br[343] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_344 bl[344] br[344] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_345 bl[345] br[345] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_346 bl[346] br[346] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_347 bl[347] br[347] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_348 bl[348] br[348] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_349 bl[349] br[349] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_350 bl[350] br[350] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_351 bl[351] br[351] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_352 bl[352] br[352] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_353 bl[353] br[353] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_354 bl[354] br[354] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_355 bl[355] br[355] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_356 bl[356] br[356] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_357 bl[357] br[357] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_358 bl[358] br[358] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_359 bl[359] br[359] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_360 bl[360] br[360] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_361 bl[361] br[361] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_362 bl[362] br[362] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_363 bl[363] br[363] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_364 bl[364] br[364] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_365 bl[365] br[365] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_366 bl[366] br[366] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_367 bl[367] br[367] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_368 bl[368] br[368] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_369 bl[369] br[369] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_370 bl[370] br[370] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_371 bl[371] br[371] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_372 bl[372] br[372] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_373 bl[373] br[373] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_374 bl[374] br[374] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_375 bl[375] br[375] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_376 bl[376] br[376] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_377 bl[377] br[377] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_378 bl[378] br[378] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_379 bl[379] br[379] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_380 bl[380] br[380] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_381 bl[381] br[381] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_382 bl[382] br[382] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_383 bl[383] br[383] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_384 bl[384] br[384] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_385 bl[385] br[385] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_386 bl[386] br[386] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_387 bl[387] br[387] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_388 bl[388] br[388] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_389 bl[389] br[389] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_390 bl[390] br[390] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_391 bl[391] br[391] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_392 bl[392] br[392] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_393 bl[393] br[393] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_394 bl[394] br[394] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_395 bl[395] br[395] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_396 bl[396] br[396] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_397 bl[397] br[397] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_398 bl[398] br[398] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_399 bl[399] br[399] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_400 bl[400] br[400] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_401 bl[401] br[401] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_402 bl[402] br[402] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_403 bl[403] br[403] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_404 bl[404] br[404] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_405 bl[405] br[405] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_406 bl[406] br[406] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_407 bl[407] br[407] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_408 bl[408] br[408] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_409 bl[409] br[409] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_410 bl[410] br[410] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_411 bl[411] br[411] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_412 bl[412] br[412] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_413 bl[413] br[413] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_414 bl[414] br[414] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_415 bl[415] br[415] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_416 bl[416] br[416] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_417 bl[417] br[417] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_418 bl[418] br[418] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_419 bl[419] br[419] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_420 bl[420] br[420] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_421 bl[421] br[421] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_422 bl[422] br[422] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_423 bl[423] br[423] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_424 bl[424] br[424] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_425 bl[425] br[425] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_426 bl[426] br[426] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_427 bl[427] br[427] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_428 bl[428] br[428] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_429 bl[429] br[429] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_430 bl[430] br[430] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_431 bl[431] br[431] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_432 bl[432] br[432] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_433 bl[433] br[433] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_434 bl[434] br[434] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_435 bl[435] br[435] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_436 bl[436] br[436] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_437 bl[437] br[437] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_438 bl[438] br[438] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_439 bl[439] br[439] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_440 bl[440] br[440] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_441 bl[441] br[441] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_442 bl[442] br[442] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_443 bl[443] br[443] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_444 bl[444] br[444] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_445 bl[445] br[445] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_446 bl[446] br[446] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_447 bl[447] br[447] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_448 bl[448] br[448] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_449 bl[449] br[449] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_450 bl[450] br[450] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_451 bl[451] br[451] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_452 bl[452] br[452] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_453 bl[453] br[453] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_454 bl[454] br[454] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_455 bl[455] br[455] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_456 bl[456] br[456] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_457 bl[457] br[457] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_458 bl[458] br[458] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_459 bl[459] br[459] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_460 bl[460] br[460] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_461 bl[461] br[461] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_462 bl[462] br[462] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_463 bl[463] br[463] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_464 bl[464] br[464] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_465 bl[465] br[465] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_466 bl[466] br[466] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_467 bl[467] br[467] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_468 bl[468] br[468] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_469 bl[469] br[469] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_470 bl[470] br[470] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_471 bl[471] br[471] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_472 bl[472] br[472] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_473 bl[473] br[473] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_474 bl[474] br[474] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_475 bl[475] br[475] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_476 bl[476] br[476] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_477 bl[477] br[477] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_478 bl[478] br[478] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_479 bl[479] br[479] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_480 bl[480] br[480] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_481 bl[481] br[481] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_482 bl[482] br[482] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_483 bl[483] br[483] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_484 bl[484] br[484] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_485 bl[485] br[485] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_486 bl[486] br[486] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_487 bl[487] br[487] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_488 bl[488] br[488] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_489 bl[489] br[489] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_490 bl[490] br[490] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_491 bl[491] br[491] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_492 bl[492] br[492] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_493 bl[493] br[493] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_494 bl[494] br[494] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_495 bl[495] br[495] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_496 bl[496] br[496] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_497 bl[497] br[497] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_498 bl[498] br[498] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_499 bl[499] br[499] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_500 bl[500] br[500] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_501 bl[501] br[501] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_502 bl[502] br[502] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_503 bl[503] br[503] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_504 bl[504] br[504] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_505 bl[505] br[505] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_506 bl[506] br[506] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_507 bl[507] br[507] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_508 bl[508] br[508] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_509 bl[509] br[509] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_510 bl[510] br[510] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_39_511 bl[511] br[511] vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xcell_40_0 bl[0] br[0] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_1 bl[1] br[1] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_2 bl[2] br[2] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_3 bl[3] br[3] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_4 bl[4] br[4] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_5 bl[5] br[5] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_6 bl[6] br[6] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_7 bl[7] br[7] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_8 bl[8] br[8] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_9 bl[9] br[9] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_10 bl[10] br[10] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_11 bl[11] br[11] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_12 bl[12] br[12] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_13 bl[13] br[13] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_14 bl[14] br[14] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_15 bl[15] br[15] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_16 bl[16] br[16] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_17 bl[17] br[17] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_18 bl[18] br[18] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_19 bl[19] br[19] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_20 bl[20] br[20] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_21 bl[21] br[21] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_22 bl[22] br[22] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_23 bl[23] br[23] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_24 bl[24] br[24] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_25 bl[25] br[25] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_26 bl[26] br[26] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_27 bl[27] br[27] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_28 bl[28] br[28] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_29 bl[29] br[29] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_30 bl[30] br[30] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_31 bl[31] br[31] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_32 bl[32] br[32] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_33 bl[33] br[33] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_34 bl[34] br[34] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_35 bl[35] br[35] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_36 bl[36] br[36] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_37 bl[37] br[37] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_38 bl[38] br[38] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_39 bl[39] br[39] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_40 bl[40] br[40] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_41 bl[41] br[41] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_42 bl[42] br[42] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_43 bl[43] br[43] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_44 bl[44] br[44] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_45 bl[45] br[45] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_46 bl[46] br[46] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_47 bl[47] br[47] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_48 bl[48] br[48] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_49 bl[49] br[49] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_50 bl[50] br[50] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_51 bl[51] br[51] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_52 bl[52] br[52] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_53 bl[53] br[53] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_54 bl[54] br[54] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_55 bl[55] br[55] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_56 bl[56] br[56] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_57 bl[57] br[57] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_58 bl[58] br[58] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_59 bl[59] br[59] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_60 bl[60] br[60] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_61 bl[61] br[61] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_62 bl[62] br[62] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_63 bl[63] br[63] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_64 bl[64] br[64] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_65 bl[65] br[65] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_66 bl[66] br[66] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_67 bl[67] br[67] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_68 bl[68] br[68] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_69 bl[69] br[69] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_70 bl[70] br[70] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_71 bl[71] br[71] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_72 bl[72] br[72] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_73 bl[73] br[73] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_74 bl[74] br[74] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_75 bl[75] br[75] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_76 bl[76] br[76] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_77 bl[77] br[77] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_78 bl[78] br[78] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_79 bl[79] br[79] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_80 bl[80] br[80] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_81 bl[81] br[81] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_82 bl[82] br[82] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_83 bl[83] br[83] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_84 bl[84] br[84] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_85 bl[85] br[85] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_86 bl[86] br[86] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_87 bl[87] br[87] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_88 bl[88] br[88] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_89 bl[89] br[89] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_90 bl[90] br[90] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_91 bl[91] br[91] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_92 bl[92] br[92] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_93 bl[93] br[93] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_94 bl[94] br[94] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_95 bl[95] br[95] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_96 bl[96] br[96] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_97 bl[97] br[97] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_98 bl[98] br[98] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_99 bl[99] br[99] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_100 bl[100] br[100] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_101 bl[101] br[101] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_102 bl[102] br[102] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_103 bl[103] br[103] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_104 bl[104] br[104] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_105 bl[105] br[105] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_106 bl[106] br[106] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_107 bl[107] br[107] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_108 bl[108] br[108] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_109 bl[109] br[109] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_110 bl[110] br[110] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_111 bl[111] br[111] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_112 bl[112] br[112] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_113 bl[113] br[113] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_114 bl[114] br[114] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_115 bl[115] br[115] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_116 bl[116] br[116] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_117 bl[117] br[117] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_118 bl[118] br[118] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_119 bl[119] br[119] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_120 bl[120] br[120] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_121 bl[121] br[121] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_122 bl[122] br[122] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_123 bl[123] br[123] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_124 bl[124] br[124] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_125 bl[125] br[125] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_126 bl[126] br[126] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_127 bl[127] br[127] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_128 bl[128] br[128] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_129 bl[129] br[129] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_130 bl[130] br[130] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_131 bl[131] br[131] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_132 bl[132] br[132] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_133 bl[133] br[133] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_134 bl[134] br[134] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_135 bl[135] br[135] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_136 bl[136] br[136] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_137 bl[137] br[137] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_138 bl[138] br[138] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_139 bl[139] br[139] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_140 bl[140] br[140] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_141 bl[141] br[141] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_142 bl[142] br[142] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_143 bl[143] br[143] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_144 bl[144] br[144] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_145 bl[145] br[145] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_146 bl[146] br[146] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_147 bl[147] br[147] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_148 bl[148] br[148] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_149 bl[149] br[149] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_150 bl[150] br[150] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_151 bl[151] br[151] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_152 bl[152] br[152] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_153 bl[153] br[153] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_154 bl[154] br[154] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_155 bl[155] br[155] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_156 bl[156] br[156] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_157 bl[157] br[157] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_158 bl[158] br[158] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_159 bl[159] br[159] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_160 bl[160] br[160] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_161 bl[161] br[161] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_162 bl[162] br[162] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_163 bl[163] br[163] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_164 bl[164] br[164] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_165 bl[165] br[165] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_166 bl[166] br[166] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_167 bl[167] br[167] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_168 bl[168] br[168] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_169 bl[169] br[169] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_170 bl[170] br[170] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_171 bl[171] br[171] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_172 bl[172] br[172] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_173 bl[173] br[173] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_174 bl[174] br[174] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_175 bl[175] br[175] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_176 bl[176] br[176] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_177 bl[177] br[177] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_178 bl[178] br[178] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_179 bl[179] br[179] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_180 bl[180] br[180] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_181 bl[181] br[181] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_182 bl[182] br[182] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_183 bl[183] br[183] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_184 bl[184] br[184] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_185 bl[185] br[185] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_186 bl[186] br[186] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_187 bl[187] br[187] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_188 bl[188] br[188] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_189 bl[189] br[189] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_190 bl[190] br[190] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_191 bl[191] br[191] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_192 bl[192] br[192] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_193 bl[193] br[193] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_194 bl[194] br[194] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_195 bl[195] br[195] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_196 bl[196] br[196] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_197 bl[197] br[197] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_198 bl[198] br[198] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_199 bl[199] br[199] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_200 bl[200] br[200] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_201 bl[201] br[201] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_202 bl[202] br[202] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_203 bl[203] br[203] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_204 bl[204] br[204] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_205 bl[205] br[205] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_206 bl[206] br[206] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_207 bl[207] br[207] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_208 bl[208] br[208] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_209 bl[209] br[209] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_210 bl[210] br[210] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_211 bl[211] br[211] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_212 bl[212] br[212] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_213 bl[213] br[213] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_214 bl[214] br[214] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_215 bl[215] br[215] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_216 bl[216] br[216] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_217 bl[217] br[217] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_218 bl[218] br[218] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_219 bl[219] br[219] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_220 bl[220] br[220] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_221 bl[221] br[221] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_222 bl[222] br[222] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_223 bl[223] br[223] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_224 bl[224] br[224] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_225 bl[225] br[225] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_226 bl[226] br[226] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_227 bl[227] br[227] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_228 bl[228] br[228] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_229 bl[229] br[229] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_230 bl[230] br[230] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_231 bl[231] br[231] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_232 bl[232] br[232] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_233 bl[233] br[233] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_234 bl[234] br[234] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_235 bl[235] br[235] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_236 bl[236] br[236] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_237 bl[237] br[237] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_238 bl[238] br[238] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_239 bl[239] br[239] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_240 bl[240] br[240] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_241 bl[241] br[241] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_242 bl[242] br[242] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_243 bl[243] br[243] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_244 bl[244] br[244] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_245 bl[245] br[245] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_246 bl[246] br[246] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_247 bl[247] br[247] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_248 bl[248] br[248] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_249 bl[249] br[249] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_250 bl[250] br[250] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_251 bl[251] br[251] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_252 bl[252] br[252] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_253 bl[253] br[253] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_254 bl[254] br[254] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_255 bl[255] br[255] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_256 bl[256] br[256] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_257 bl[257] br[257] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_258 bl[258] br[258] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_259 bl[259] br[259] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_260 bl[260] br[260] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_261 bl[261] br[261] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_262 bl[262] br[262] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_263 bl[263] br[263] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_264 bl[264] br[264] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_265 bl[265] br[265] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_266 bl[266] br[266] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_267 bl[267] br[267] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_268 bl[268] br[268] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_269 bl[269] br[269] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_270 bl[270] br[270] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_271 bl[271] br[271] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_272 bl[272] br[272] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_273 bl[273] br[273] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_274 bl[274] br[274] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_275 bl[275] br[275] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_276 bl[276] br[276] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_277 bl[277] br[277] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_278 bl[278] br[278] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_279 bl[279] br[279] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_280 bl[280] br[280] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_281 bl[281] br[281] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_282 bl[282] br[282] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_283 bl[283] br[283] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_284 bl[284] br[284] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_285 bl[285] br[285] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_286 bl[286] br[286] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_287 bl[287] br[287] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_288 bl[288] br[288] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_289 bl[289] br[289] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_290 bl[290] br[290] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_291 bl[291] br[291] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_292 bl[292] br[292] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_293 bl[293] br[293] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_294 bl[294] br[294] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_295 bl[295] br[295] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_296 bl[296] br[296] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_297 bl[297] br[297] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_298 bl[298] br[298] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_299 bl[299] br[299] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_300 bl[300] br[300] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_301 bl[301] br[301] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_302 bl[302] br[302] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_303 bl[303] br[303] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_304 bl[304] br[304] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_305 bl[305] br[305] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_306 bl[306] br[306] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_307 bl[307] br[307] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_308 bl[308] br[308] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_309 bl[309] br[309] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_310 bl[310] br[310] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_311 bl[311] br[311] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_312 bl[312] br[312] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_313 bl[313] br[313] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_314 bl[314] br[314] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_315 bl[315] br[315] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_316 bl[316] br[316] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_317 bl[317] br[317] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_318 bl[318] br[318] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_319 bl[319] br[319] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_320 bl[320] br[320] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_321 bl[321] br[321] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_322 bl[322] br[322] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_323 bl[323] br[323] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_324 bl[324] br[324] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_325 bl[325] br[325] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_326 bl[326] br[326] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_327 bl[327] br[327] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_328 bl[328] br[328] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_329 bl[329] br[329] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_330 bl[330] br[330] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_331 bl[331] br[331] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_332 bl[332] br[332] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_333 bl[333] br[333] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_334 bl[334] br[334] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_335 bl[335] br[335] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_336 bl[336] br[336] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_337 bl[337] br[337] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_338 bl[338] br[338] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_339 bl[339] br[339] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_340 bl[340] br[340] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_341 bl[341] br[341] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_342 bl[342] br[342] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_343 bl[343] br[343] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_344 bl[344] br[344] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_345 bl[345] br[345] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_346 bl[346] br[346] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_347 bl[347] br[347] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_348 bl[348] br[348] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_349 bl[349] br[349] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_350 bl[350] br[350] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_351 bl[351] br[351] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_352 bl[352] br[352] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_353 bl[353] br[353] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_354 bl[354] br[354] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_355 bl[355] br[355] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_356 bl[356] br[356] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_357 bl[357] br[357] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_358 bl[358] br[358] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_359 bl[359] br[359] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_360 bl[360] br[360] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_361 bl[361] br[361] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_362 bl[362] br[362] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_363 bl[363] br[363] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_364 bl[364] br[364] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_365 bl[365] br[365] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_366 bl[366] br[366] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_367 bl[367] br[367] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_368 bl[368] br[368] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_369 bl[369] br[369] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_370 bl[370] br[370] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_371 bl[371] br[371] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_372 bl[372] br[372] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_373 bl[373] br[373] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_374 bl[374] br[374] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_375 bl[375] br[375] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_376 bl[376] br[376] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_377 bl[377] br[377] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_378 bl[378] br[378] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_379 bl[379] br[379] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_380 bl[380] br[380] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_381 bl[381] br[381] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_382 bl[382] br[382] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_383 bl[383] br[383] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_384 bl[384] br[384] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_385 bl[385] br[385] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_386 bl[386] br[386] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_387 bl[387] br[387] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_388 bl[388] br[388] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_389 bl[389] br[389] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_390 bl[390] br[390] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_391 bl[391] br[391] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_392 bl[392] br[392] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_393 bl[393] br[393] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_394 bl[394] br[394] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_395 bl[395] br[395] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_396 bl[396] br[396] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_397 bl[397] br[397] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_398 bl[398] br[398] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_399 bl[399] br[399] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_400 bl[400] br[400] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_401 bl[401] br[401] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_402 bl[402] br[402] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_403 bl[403] br[403] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_404 bl[404] br[404] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_405 bl[405] br[405] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_406 bl[406] br[406] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_407 bl[407] br[407] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_408 bl[408] br[408] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_409 bl[409] br[409] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_410 bl[410] br[410] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_411 bl[411] br[411] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_412 bl[412] br[412] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_413 bl[413] br[413] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_414 bl[414] br[414] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_415 bl[415] br[415] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_416 bl[416] br[416] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_417 bl[417] br[417] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_418 bl[418] br[418] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_419 bl[419] br[419] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_420 bl[420] br[420] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_421 bl[421] br[421] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_422 bl[422] br[422] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_423 bl[423] br[423] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_424 bl[424] br[424] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_425 bl[425] br[425] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_426 bl[426] br[426] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_427 bl[427] br[427] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_428 bl[428] br[428] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_429 bl[429] br[429] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_430 bl[430] br[430] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_431 bl[431] br[431] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_432 bl[432] br[432] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_433 bl[433] br[433] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_434 bl[434] br[434] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_435 bl[435] br[435] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_436 bl[436] br[436] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_437 bl[437] br[437] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_438 bl[438] br[438] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_439 bl[439] br[439] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_440 bl[440] br[440] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_441 bl[441] br[441] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_442 bl[442] br[442] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_443 bl[443] br[443] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_444 bl[444] br[444] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_445 bl[445] br[445] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_446 bl[446] br[446] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_447 bl[447] br[447] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_448 bl[448] br[448] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_449 bl[449] br[449] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_450 bl[450] br[450] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_451 bl[451] br[451] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_452 bl[452] br[452] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_453 bl[453] br[453] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_454 bl[454] br[454] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_455 bl[455] br[455] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_456 bl[456] br[456] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_457 bl[457] br[457] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_458 bl[458] br[458] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_459 bl[459] br[459] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_460 bl[460] br[460] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_461 bl[461] br[461] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_462 bl[462] br[462] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_463 bl[463] br[463] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_464 bl[464] br[464] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_465 bl[465] br[465] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_466 bl[466] br[466] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_467 bl[467] br[467] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_468 bl[468] br[468] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_469 bl[469] br[469] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_470 bl[470] br[470] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_471 bl[471] br[471] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_472 bl[472] br[472] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_473 bl[473] br[473] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_474 bl[474] br[474] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_475 bl[475] br[475] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_476 bl[476] br[476] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_477 bl[477] br[477] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_478 bl[478] br[478] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_479 bl[479] br[479] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_480 bl[480] br[480] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_481 bl[481] br[481] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_482 bl[482] br[482] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_483 bl[483] br[483] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_484 bl[484] br[484] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_485 bl[485] br[485] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_486 bl[486] br[486] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_487 bl[487] br[487] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_488 bl[488] br[488] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_489 bl[489] br[489] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_490 bl[490] br[490] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_491 bl[491] br[491] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_492 bl[492] br[492] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_493 bl[493] br[493] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_494 bl[494] br[494] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_495 bl[495] br[495] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_496 bl[496] br[496] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_497 bl[497] br[497] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_498 bl[498] br[498] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_499 bl[499] br[499] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_500 bl[500] br[500] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_501 bl[501] br[501] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_502 bl[502] br[502] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_503 bl[503] br[503] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_504 bl[504] br[504] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_505 bl[505] br[505] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_506 bl[506] br[506] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_507 bl[507] br[507] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_508 bl[508] br[508] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_509 bl[509] br[509] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_510 bl[510] br[510] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_40_511 bl[511] br[511] vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xcell_41_0 bl[0] br[0] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_1 bl[1] br[1] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_2 bl[2] br[2] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_3 bl[3] br[3] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_4 bl[4] br[4] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_5 bl[5] br[5] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_6 bl[6] br[6] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_7 bl[7] br[7] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_8 bl[8] br[8] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_9 bl[9] br[9] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_10 bl[10] br[10] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_11 bl[11] br[11] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_12 bl[12] br[12] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_13 bl[13] br[13] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_14 bl[14] br[14] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_15 bl[15] br[15] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_16 bl[16] br[16] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_17 bl[17] br[17] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_18 bl[18] br[18] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_19 bl[19] br[19] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_20 bl[20] br[20] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_21 bl[21] br[21] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_22 bl[22] br[22] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_23 bl[23] br[23] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_24 bl[24] br[24] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_25 bl[25] br[25] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_26 bl[26] br[26] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_27 bl[27] br[27] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_28 bl[28] br[28] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_29 bl[29] br[29] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_30 bl[30] br[30] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_31 bl[31] br[31] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_32 bl[32] br[32] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_33 bl[33] br[33] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_34 bl[34] br[34] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_35 bl[35] br[35] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_36 bl[36] br[36] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_37 bl[37] br[37] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_38 bl[38] br[38] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_39 bl[39] br[39] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_40 bl[40] br[40] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_41 bl[41] br[41] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_42 bl[42] br[42] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_43 bl[43] br[43] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_44 bl[44] br[44] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_45 bl[45] br[45] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_46 bl[46] br[46] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_47 bl[47] br[47] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_48 bl[48] br[48] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_49 bl[49] br[49] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_50 bl[50] br[50] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_51 bl[51] br[51] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_52 bl[52] br[52] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_53 bl[53] br[53] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_54 bl[54] br[54] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_55 bl[55] br[55] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_56 bl[56] br[56] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_57 bl[57] br[57] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_58 bl[58] br[58] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_59 bl[59] br[59] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_60 bl[60] br[60] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_61 bl[61] br[61] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_62 bl[62] br[62] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_63 bl[63] br[63] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_64 bl[64] br[64] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_65 bl[65] br[65] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_66 bl[66] br[66] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_67 bl[67] br[67] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_68 bl[68] br[68] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_69 bl[69] br[69] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_70 bl[70] br[70] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_71 bl[71] br[71] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_72 bl[72] br[72] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_73 bl[73] br[73] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_74 bl[74] br[74] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_75 bl[75] br[75] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_76 bl[76] br[76] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_77 bl[77] br[77] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_78 bl[78] br[78] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_79 bl[79] br[79] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_80 bl[80] br[80] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_81 bl[81] br[81] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_82 bl[82] br[82] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_83 bl[83] br[83] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_84 bl[84] br[84] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_85 bl[85] br[85] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_86 bl[86] br[86] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_87 bl[87] br[87] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_88 bl[88] br[88] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_89 bl[89] br[89] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_90 bl[90] br[90] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_91 bl[91] br[91] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_92 bl[92] br[92] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_93 bl[93] br[93] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_94 bl[94] br[94] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_95 bl[95] br[95] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_96 bl[96] br[96] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_97 bl[97] br[97] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_98 bl[98] br[98] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_99 bl[99] br[99] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_100 bl[100] br[100] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_101 bl[101] br[101] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_102 bl[102] br[102] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_103 bl[103] br[103] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_104 bl[104] br[104] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_105 bl[105] br[105] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_106 bl[106] br[106] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_107 bl[107] br[107] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_108 bl[108] br[108] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_109 bl[109] br[109] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_110 bl[110] br[110] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_111 bl[111] br[111] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_112 bl[112] br[112] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_113 bl[113] br[113] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_114 bl[114] br[114] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_115 bl[115] br[115] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_116 bl[116] br[116] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_117 bl[117] br[117] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_118 bl[118] br[118] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_119 bl[119] br[119] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_120 bl[120] br[120] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_121 bl[121] br[121] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_122 bl[122] br[122] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_123 bl[123] br[123] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_124 bl[124] br[124] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_125 bl[125] br[125] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_126 bl[126] br[126] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_127 bl[127] br[127] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_128 bl[128] br[128] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_129 bl[129] br[129] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_130 bl[130] br[130] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_131 bl[131] br[131] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_132 bl[132] br[132] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_133 bl[133] br[133] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_134 bl[134] br[134] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_135 bl[135] br[135] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_136 bl[136] br[136] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_137 bl[137] br[137] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_138 bl[138] br[138] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_139 bl[139] br[139] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_140 bl[140] br[140] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_141 bl[141] br[141] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_142 bl[142] br[142] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_143 bl[143] br[143] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_144 bl[144] br[144] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_145 bl[145] br[145] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_146 bl[146] br[146] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_147 bl[147] br[147] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_148 bl[148] br[148] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_149 bl[149] br[149] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_150 bl[150] br[150] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_151 bl[151] br[151] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_152 bl[152] br[152] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_153 bl[153] br[153] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_154 bl[154] br[154] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_155 bl[155] br[155] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_156 bl[156] br[156] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_157 bl[157] br[157] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_158 bl[158] br[158] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_159 bl[159] br[159] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_160 bl[160] br[160] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_161 bl[161] br[161] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_162 bl[162] br[162] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_163 bl[163] br[163] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_164 bl[164] br[164] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_165 bl[165] br[165] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_166 bl[166] br[166] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_167 bl[167] br[167] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_168 bl[168] br[168] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_169 bl[169] br[169] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_170 bl[170] br[170] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_171 bl[171] br[171] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_172 bl[172] br[172] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_173 bl[173] br[173] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_174 bl[174] br[174] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_175 bl[175] br[175] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_176 bl[176] br[176] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_177 bl[177] br[177] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_178 bl[178] br[178] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_179 bl[179] br[179] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_180 bl[180] br[180] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_181 bl[181] br[181] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_182 bl[182] br[182] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_183 bl[183] br[183] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_184 bl[184] br[184] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_185 bl[185] br[185] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_186 bl[186] br[186] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_187 bl[187] br[187] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_188 bl[188] br[188] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_189 bl[189] br[189] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_190 bl[190] br[190] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_191 bl[191] br[191] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_192 bl[192] br[192] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_193 bl[193] br[193] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_194 bl[194] br[194] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_195 bl[195] br[195] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_196 bl[196] br[196] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_197 bl[197] br[197] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_198 bl[198] br[198] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_199 bl[199] br[199] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_200 bl[200] br[200] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_201 bl[201] br[201] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_202 bl[202] br[202] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_203 bl[203] br[203] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_204 bl[204] br[204] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_205 bl[205] br[205] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_206 bl[206] br[206] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_207 bl[207] br[207] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_208 bl[208] br[208] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_209 bl[209] br[209] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_210 bl[210] br[210] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_211 bl[211] br[211] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_212 bl[212] br[212] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_213 bl[213] br[213] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_214 bl[214] br[214] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_215 bl[215] br[215] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_216 bl[216] br[216] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_217 bl[217] br[217] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_218 bl[218] br[218] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_219 bl[219] br[219] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_220 bl[220] br[220] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_221 bl[221] br[221] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_222 bl[222] br[222] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_223 bl[223] br[223] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_224 bl[224] br[224] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_225 bl[225] br[225] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_226 bl[226] br[226] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_227 bl[227] br[227] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_228 bl[228] br[228] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_229 bl[229] br[229] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_230 bl[230] br[230] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_231 bl[231] br[231] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_232 bl[232] br[232] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_233 bl[233] br[233] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_234 bl[234] br[234] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_235 bl[235] br[235] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_236 bl[236] br[236] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_237 bl[237] br[237] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_238 bl[238] br[238] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_239 bl[239] br[239] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_240 bl[240] br[240] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_241 bl[241] br[241] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_242 bl[242] br[242] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_243 bl[243] br[243] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_244 bl[244] br[244] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_245 bl[245] br[245] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_246 bl[246] br[246] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_247 bl[247] br[247] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_248 bl[248] br[248] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_249 bl[249] br[249] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_250 bl[250] br[250] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_251 bl[251] br[251] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_252 bl[252] br[252] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_253 bl[253] br[253] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_254 bl[254] br[254] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_255 bl[255] br[255] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_256 bl[256] br[256] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_257 bl[257] br[257] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_258 bl[258] br[258] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_259 bl[259] br[259] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_260 bl[260] br[260] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_261 bl[261] br[261] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_262 bl[262] br[262] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_263 bl[263] br[263] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_264 bl[264] br[264] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_265 bl[265] br[265] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_266 bl[266] br[266] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_267 bl[267] br[267] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_268 bl[268] br[268] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_269 bl[269] br[269] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_270 bl[270] br[270] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_271 bl[271] br[271] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_272 bl[272] br[272] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_273 bl[273] br[273] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_274 bl[274] br[274] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_275 bl[275] br[275] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_276 bl[276] br[276] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_277 bl[277] br[277] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_278 bl[278] br[278] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_279 bl[279] br[279] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_280 bl[280] br[280] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_281 bl[281] br[281] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_282 bl[282] br[282] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_283 bl[283] br[283] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_284 bl[284] br[284] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_285 bl[285] br[285] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_286 bl[286] br[286] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_287 bl[287] br[287] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_288 bl[288] br[288] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_289 bl[289] br[289] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_290 bl[290] br[290] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_291 bl[291] br[291] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_292 bl[292] br[292] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_293 bl[293] br[293] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_294 bl[294] br[294] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_295 bl[295] br[295] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_296 bl[296] br[296] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_297 bl[297] br[297] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_298 bl[298] br[298] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_299 bl[299] br[299] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_300 bl[300] br[300] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_301 bl[301] br[301] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_302 bl[302] br[302] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_303 bl[303] br[303] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_304 bl[304] br[304] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_305 bl[305] br[305] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_306 bl[306] br[306] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_307 bl[307] br[307] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_308 bl[308] br[308] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_309 bl[309] br[309] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_310 bl[310] br[310] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_311 bl[311] br[311] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_312 bl[312] br[312] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_313 bl[313] br[313] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_314 bl[314] br[314] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_315 bl[315] br[315] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_316 bl[316] br[316] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_317 bl[317] br[317] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_318 bl[318] br[318] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_319 bl[319] br[319] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_320 bl[320] br[320] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_321 bl[321] br[321] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_322 bl[322] br[322] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_323 bl[323] br[323] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_324 bl[324] br[324] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_325 bl[325] br[325] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_326 bl[326] br[326] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_327 bl[327] br[327] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_328 bl[328] br[328] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_329 bl[329] br[329] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_330 bl[330] br[330] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_331 bl[331] br[331] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_332 bl[332] br[332] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_333 bl[333] br[333] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_334 bl[334] br[334] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_335 bl[335] br[335] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_336 bl[336] br[336] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_337 bl[337] br[337] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_338 bl[338] br[338] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_339 bl[339] br[339] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_340 bl[340] br[340] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_341 bl[341] br[341] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_342 bl[342] br[342] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_343 bl[343] br[343] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_344 bl[344] br[344] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_345 bl[345] br[345] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_346 bl[346] br[346] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_347 bl[347] br[347] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_348 bl[348] br[348] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_349 bl[349] br[349] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_350 bl[350] br[350] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_351 bl[351] br[351] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_352 bl[352] br[352] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_353 bl[353] br[353] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_354 bl[354] br[354] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_355 bl[355] br[355] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_356 bl[356] br[356] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_357 bl[357] br[357] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_358 bl[358] br[358] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_359 bl[359] br[359] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_360 bl[360] br[360] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_361 bl[361] br[361] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_362 bl[362] br[362] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_363 bl[363] br[363] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_364 bl[364] br[364] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_365 bl[365] br[365] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_366 bl[366] br[366] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_367 bl[367] br[367] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_368 bl[368] br[368] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_369 bl[369] br[369] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_370 bl[370] br[370] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_371 bl[371] br[371] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_372 bl[372] br[372] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_373 bl[373] br[373] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_374 bl[374] br[374] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_375 bl[375] br[375] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_376 bl[376] br[376] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_377 bl[377] br[377] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_378 bl[378] br[378] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_379 bl[379] br[379] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_380 bl[380] br[380] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_381 bl[381] br[381] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_382 bl[382] br[382] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_383 bl[383] br[383] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_384 bl[384] br[384] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_385 bl[385] br[385] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_386 bl[386] br[386] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_387 bl[387] br[387] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_388 bl[388] br[388] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_389 bl[389] br[389] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_390 bl[390] br[390] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_391 bl[391] br[391] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_392 bl[392] br[392] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_393 bl[393] br[393] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_394 bl[394] br[394] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_395 bl[395] br[395] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_396 bl[396] br[396] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_397 bl[397] br[397] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_398 bl[398] br[398] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_399 bl[399] br[399] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_400 bl[400] br[400] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_401 bl[401] br[401] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_402 bl[402] br[402] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_403 bl[403] br[403] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_404 bl[404] br[404] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_405 bl[405] br[405] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_406 bl[406] br[406] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_407 bl[407] br[407] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_408 bl[408] br[408] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_409 bl[409] br[409] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_410 bl[410] br[410] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_411 bl[411] br[411] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_412 bl[412] br[412] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_413 bl[413] br[413] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_414 bl[414] br[414] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_415 bl[415] br[415] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_416 bl[416] br[416] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_417 bl[417] br[417] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_418 bl[418] br[418] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_419 bl[419] br[419] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_420 bl[420] br[420] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_421 bl[421] br[421] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_422 bl[422] br[422] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_423 bl[423] br[423] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_424 bl[424] br[424] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_425 bl[425] br[425] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_426 bl[426] br[426] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_427 bl[427] br[427] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_428 bl[428] br[428] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_429 bl[429] br[429] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_430 bl[430] br[430] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_431 bl[431] br[431] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_432 bl[432] br[432] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_433 bl[433] br[433] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_434 bl[434] br[434] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_435 bl[435] br[435] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_436 bl[436] br[436] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_437 bl[437] br[437] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_438 bl[438] br[438] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_439 bl[439] br[439] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_440 bl[440] br[440] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_441 bl[441] br[441] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_442 bl[442] br[442] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_443 bl[443] br[443] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_444 bl[444] br[444] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_445 bl[445] br[445] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_446 bl[446] br[446] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_447 bl[447] br[447] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_448 bl[448] br[448] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_449 bl[449] br[449] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_450 bl[450] br[450] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_451 bl[451] br[451] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_452 bl[452] br[452] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_453 bl[453] br[453] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_454 bl[454] br[454] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_455 bl[455] br[455] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_456 bl[456] br[456] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_457 bl[457] br[457] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_458 bl[458] br[458] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_459 bl[459] br[459] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_460 bl[460] br[460] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_461 bl[461] br[461] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_462 bl[462] br[462] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_463 bl[463] br[463] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_464 bl[464] br[464] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_465 bl[465] br[465] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_466 bl[466] br[466] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_467 bl[467] br[467] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_468 bl[468] br[468] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_469 bl[469] br[469] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_470 bl[470] br[470] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_471 bl[471] br[471] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_472 bl[472] br[472] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_473 bl[473] br[473] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_474 bl[474] br[474] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_475 bl[475] br[475] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_476 bl[476] br[476] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_477 bl[477] br[477] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_478 bl[478] br[478] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_479 bl[479] br[479] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_480 bl[480] br[480] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_481 bl[481] br[481] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_482 bl[482] br[482] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_483 bl[483] br[483] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_484 bl[484] br[484] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_485 bl[485] br[485] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_486 bl[486] br[486] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_487 bl[487] br[487] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_488 bl[488] br[488] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_489 bl[489] br[489] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_490 bl[490] br[490] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_491 bl[491] br[491] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_492 bl[492] br[492] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_493 bl[493] br[493] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_494 bl[494] br[494] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_495 bl[495] br[495] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_496 bl[496] br[496] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_497 bl[497] br[497] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_498 bl[498] br[498] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_499 bl[499] br[499] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_500 bl[500] br[500] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_501 bl[501] br[501] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_502 bl[502] br[502] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_503 bl[503] br[503] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_504 bl[504] br[504] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_505 bl[505] br[505] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_506 bl[506] br[506] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_507 bl[507] br[507] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_508 bl[508] br[508] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_509 bl[509] br[509] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_510 bl[510] br[510] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_41_511 bl[511] br[511] vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xcell_42_0 bl[0] br[0] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_1 bl[1] br[1] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_2 bl[2] br[2] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_3 bl[3] br[3] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_4 bl[4] br[4] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_5 bl[5] br[5] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_6 bl[6] br[6] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_7 bl[7] br[7] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_8 bl[8] br[8] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_9 bl[9] br[9] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_10 bl[10] br[10] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_11 bl[11] br[11] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_12 bl[12] br[12] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_13 bl[13] br[13] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_14 bl[14] br[14] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_15 bl[15] br[15] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_16 bl[16] br[16] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_17 bl[17] br[17] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_18 bl[18] br[18] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_19 bl[19] br[19] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_20 bl[20] br[20] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_21 bl[21] br[21] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_22 bl[22] br[22] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_23 bl[23] br[23] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_24 bl[24] br[24] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_25 bl[25] br[25] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_26 bl[26] br[26] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_27 bl[27] br[27] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_28 bl[28] br[28] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_29 bl[29] br[29] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_30 bl[30] br[30] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_31 bl[31] br[31] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_32 bl[32] br[32] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_33 bl[33] br[33] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_34 bl[34] br[34] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_35 bl[35] br[35] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_36 bl[36] br[36] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_37 bl[37] br[37] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_38 bl[38] br[38] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_39 bl[39] br[39] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_40 bl[40] br[40] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_41 bl[41] br[41] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_42 bl[42] br[42] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_43 bl[43] br[43] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_44 bl[44] br[44] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_45 bl[45] br[45] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_46 bl[46] br[46] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_47 bl[47] br[47] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_48 bl[48] br[48] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_49 bl[49] br[49] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_50 bl[50] br[50] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_51 bl[51] br[51] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_52 bl[52] br[52] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_53 bl[53] br[53] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_54 bl[54] br[54] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_55 bl[55] br[55] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_56 bl[56] br[56] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_57 bl[57] br[57] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_58 bl[58] br[58] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_59 bl[59] br[59] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_60 bl[60] br[60] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_61 bl[61] br[61] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_62 bl[62] br[62] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_63 bl[63] br[63] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_64 bl[64] br[64] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_65 bl[65] br[65] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_66 bl[66] br[66] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_67 bl[67] br[67] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_68 bl[68] br[68] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_69 bl[69] br[69] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_70 bl[70] br[70] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_71 bl[71] br[71] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_72 bl[72] br[72] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_73 bl[73] br[73] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_74 bl[74] br[74] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_75 bl[75] br[75] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_76 bl[76] br[76] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_77 bl[77] br[77] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_78 bl[78] br[78] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_79 bl[79] br[79] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_80 bl[80] br[80] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_81 bl[81] br[81] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_82 bl[82] br[82] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_83 bl[83] br[83] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_84 bl[84] br[84] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_85 bl[85] br[85] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_86 bl[86] br[86] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_87 bl[87] br[87] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_88 bl[88] br[88] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_89 bl[89] br[89] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_90 bl[90] br[90] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_91 bl[91] br[91] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_92 bl[92] br[92] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_93 bl[93] br[93] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_94 bl[94] br[94] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_95 bl[95] br[95] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_96 bl[96] br[96] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_97 bl[97] br[97] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_98 bl[98] br[98] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_99 bl[99] br[99] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_100 bl[100] br[100] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_101 bl[101] br[101] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_102 bl[102] br[102] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_103 bl[103] br[103] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_104 bl[104] br[104] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_105 bl[105] br[105] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_106 bl[106] br[106] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_107 bl[107] br[107] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_108 bl[108] br[108] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_109 bl[109] br[109] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_110 bl[110] br[110] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_111 bl[111] br[111] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_112 bl[112] br[112] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_113 bl[113] br[113] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_114 bl[114] br[114] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_115 bl[115] br[115] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_116 bl[116] br[116] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_117 bl[117] br[117] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_118 bl[118] br[118] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_119 bl[119] br[119] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_120 bl[120] br[120] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_121 bl[121] br[121] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_122 bl[122] br[122] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_123 bl[123] br[123] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_124 bl[124] br[124] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_125 bl[125] br[125] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_126 bl[126] br[126] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_127 bl[127] br[127] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_128 bl[128] br[128] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_129 bl[129] br[129] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_130 bl[130] br[130] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_131 bl[131] br[131] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_132 bl[132] br[132] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_133 bl[133] br[133] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_134 bl[134] br[134] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_135 bl[135] br[135] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_136 bl[136] br[136] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_137 bl[137] br[137] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_138 bl[138] br[138] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_139 bl[139] br[139] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_140 bl[140] br[140] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_141 bl[141] br[141] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_142 bl[142] br[142] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_143 bl[143] br[143] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_144 bl[144] br[144] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_145 bl[145] br[145] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_146 bl[146] br[146] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_147 bl[147] br[147] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_148 bl[148] br[148] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_149 bl[149] br[149] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_150 bl[150] br[150] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_151 bl[151] br[151] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_152 bl[152] br[152] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_153 bl[153] br[153] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_154 bl[154] br[154] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_155 bl[155] br[155] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_156 bl[156] br[156] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_157 bl[157] br[157] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_158 bl[158] br[158] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_159 bl[159] br[159] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_160 bl[160] br[160] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_161 bl[161] br[161] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_162 bl[162] br[162] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_163 bl[163] br[163] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_164 bl[164] br[164] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_165 bl[165] br[165] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_166 bl[166] br[166] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_167 bl[167] br[167] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_168 bl[168] br[168] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_169 bl[169] br[169] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_170 bl[170] br[170] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_171 bl[171] br[171] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_172 bl[172] br[172] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_173 bl[173] br[173] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_174 bl[174] br[174] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_175 bl[175] br[175] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_176 bl[176] br[176] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_177 bl[177] br[177] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_178 bl[178] br[178] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_179 bl[179] br[179] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_180 bl[180] br[180] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_181 bl[181] br[181] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_182 bl[182] br[182] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_183 bl[183] br[183] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_184 bl[184] br[184] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_185 bl[185] br[185] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_186 bl[186] br[186] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_187 bl[187] br[187] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_188 bl[188] br[188] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_189 bl[189] br[189] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_190 bl[190] br[190] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_191 bl[191] br[191] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_192 bl[192] br[192] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_193 bl[193] br[193] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_194 bl[194] br[194] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_195 bl[195] br[195] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_196 bl[196] br[196] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_197 bl[197] br[197] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_198 bl[198] br[198] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_199 bl[199] br[199] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_200 bl[200] br[200] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_201 bl[201] br[201] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_202 bl[202] br[202] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_203 bl[203] br[203] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_204 bl[204] br[204] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_205 bl[205] br[205] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_206 bl[206] br[206] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_207 bl[207] br[207] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_208 bl[208] br[208] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_209 bl[209] br[209] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_210 bl[210] br[210] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_211 bl[211] br[211] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_212 bl[212] br[212] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_213 bl[213] br[213] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_214 bl[214] br[214] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_215 bl[215] br[215] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_216 bl[216] br[216] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_217 bl[217] br[217] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_218 bl[218] br[218] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_219 bl[219] br[219] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_220 bl[220] br[220] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_221 bl[221] br[221] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_222 bl[222] br[222] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_223 bl[223] br[223] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_224 bl[224] br[224] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_225 bl[225] br[225] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_226 bl[226] br[226] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_227 bl[227] br[227] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_228 bl[228] br[228] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_229 bl[229] br[229] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_230 bl[230] br[230] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_231 bl[231] br[231] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_232 bl[232] br[232] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_233 bl[233] br[233] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_234 bl[234] br[234] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_235 bl[235] br[235] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_236 bl[236] br[236] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_237 bl[237] br[237] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_238 bl[238] br[238] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_239 bl[239] br[239] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_240 bl[240] br[240] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_241 bl[241] br[241] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_242 bl[242] br[242] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_243 bl[243] br[243] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_244 bl[244] br[244] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_245 bl[245] br[245] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_246 bl[246] br[246] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_247 bl[247] br[247] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_248 bl[248] br[248] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_249 bl[249] br[249] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_250 bl[250] br[250] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_251 bl[251] br[251] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_252 bl[252] br[252] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_253 bl[253] br[253] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_254 bl[254] br[254] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_255 bl[255] br[255] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_256 bl[256] br[256] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_257 bl[257] br[257] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_258 bl[258] br[258] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_259 bl[259] br[259] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_260 bl[260] br[260] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_261 bl[261] br[261] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_262 bl[262] br[262] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_263 bl[263] br[263] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_264 bl[264] br[264] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_265 bl[265] br[265] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_266 bl[266] br[266] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_267 bl[267] br[267] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_268 bl[268] br[268] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_269 bl[269] br[269] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_270 bl[270] br[270] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_271 bl[271] br[271] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_272 bl[272] br[272] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_273 bl[273] br[273] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_274 bl[274] br[274] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_275 bl[275] br[275] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_276 bl[276] br[276] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_277 bl[277] br[277] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_278 bl[278] br[278] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_279 bl[279] br[279] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_280 bl[280] br[280] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_281 bl[281] br[281] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_282 bl[282] br[282] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_283 bl[283] br[283] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_284 bl[284] br[284] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_285 bl[285] br[285] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_286 bl[286] br[286] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_287 bl[287] br[287] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_288 bl[288] br[288] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_289 bl[289] br[289] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_290 bl[290] br[290] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_291 bl[291] br[291] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_292 bl[292] br[292] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_293 bl[293] br[293] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_294 bl[294] br[294] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_295 bl[295] br[295] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_296 bl[296] br[296] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_297 bl[297] br[297] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_298 bl[298] br[298] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_299 bl[299] br[299] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_300 bl[300] br[300] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_301 bl[301] br[301] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_302 bl[302] br[302] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_303 bl[303] br[303] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_304 bl[304] br[304] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_305 bl[305] br[305] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_306 bl[306] br[306] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_307 bl[307] br[307] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_308 bl[308] br[308] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_309 bl[309] br[309] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_310 bl[310] br[310] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_311 bl[311] br[311] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_312 bl[312] br[312] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_313 bl[313] br[313] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_314 bl[314] br[314] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_315 bl[315] br[315] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_316 bl[316] br[316] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_317 bl[317] br[317] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_318 bl[318] br[318] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_319 bl[319] br[319] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_320 bl[320] br[320] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_321 bl[321] br[321] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_322 bl[322] br[322] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_323 bl[323] br[323] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_324 bl[324] br[324] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_325 bl[325] br[325] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_326 bl[326] br[326] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_327 bl[327] br[327] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_328 bl[328] br[328] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_329 bl[329] br[329] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_330 bl[330] br[330] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_331 bl[331] br[331] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_332 bl[332] br[332] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_333 bl[333] br[333] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_334 bl[334] br[334] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_335 bl[335] br[335] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_336 bl[336] br[336] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_337 bl[337] br[337] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_338 bl[338] br[338] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_339 bl[339] br[339] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_340 bl[340] br[340] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_341 bl[341] br[341] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_342 bl[342] br[342] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_343 bl[343] br[343] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_344 bl[344] br[344] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_345 bl[345] br[345] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_346 bl[346] br[346] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_347 bl[347] br[347] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_348 bl[348] br[348] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_349 bl[349] br[349] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_350 bl[350] br[350] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_351 bl[351] br[351] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_352 bl[352] br[352] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_353 bl[353] br[353] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_354 bl[354] br[354] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_355 bl[355] br[355] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_356 bl[356] br[356] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_357 bl[357] br[357] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_358 bl[358] br[358] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_359 bl[359] br[359] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_360 bl[360] br[360] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_361 bl[361] br[361] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_362 bl[362] br[362] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_363 bl[363] br[363] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_364 bl[364] br[364] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_365 bl[365] br[365] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_366 bl[366] br[366] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_367 bl[367] br[367] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_368 bl[368] br[368] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_369 bl[369] br[369] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_370 bl[370] br[370] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_371 bl[371] br[371] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_372 bl[372] br[372] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_373 bl[373] br[373] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_374 bl[374] br[374] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_375 bl[375] br[375] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_376 bl[376] br[376] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_377 bl[377] br[377] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_378 bl[378] br[378] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_379 bl[379] br[379] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_380 bl[380] br[380] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_381 bl[381] br[381] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_382 bl[382] br[382] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_383 bl[383] br[383] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_384 bl[384] br[384] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_385 bl[385] br[385] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_386 bl[386] br[386] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_387 bl[387] br[387] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_388 bl[388] br[388] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_389 bl[389] br[389] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_390 bl[390] br[390] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_391 bl[391] br[391] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_392 bl[392] br[392] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_393 bl[393] br[393] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_394 bl[394] br[394] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_395 bl[395] br[395] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_396 bl[396] br[396] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_397 bl[397] br[397] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_398 bl[398] br[398] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_399 bl[399] br[399] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_400 bl[400] br[400] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_401 bl[401] br[401] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_402 bl[402] br[402] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_403 bl[403] br[403] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_404 bl[404] br[404] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_405 bl[405] br[405] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_406 bl[406] br[406] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_407 bl[407] br[407] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_408 bl[408] br[408] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_409 bl[409] br[409] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_410 bl[410] br[410] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_411 bl[411] br[411] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_412 bl[412] br[412] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_413 bl[413] br[413] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_414 bl[414] br[414] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_415 bl[415] br[415] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_416 bl[416] br[416] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_417 bl[417] br[417] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_418 bl[418] br[418] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_419 bl[419] br[419] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_420 bl[420] br[420] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_421 bl[421] br[421] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_422 bl[422] br[422] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_423 bl[423] br[423] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_424 bl[424] br[424] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_425 bl[425] br[425] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_426 bl[426] br[426] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_427 bl[427] br[427] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_428 bl[428] br[428] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_429 bl[429] br[429] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_430 bl[430] br[430] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_431 bl[431] br[431] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_432 bl[432] br[432] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_433 bl[433] br[433] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_434 bl[434] br[434] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_435 bl[435] br[435] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_436 bl[436] br[436] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_437 bl[437] br[437] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_438 bl[438] br[438] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_439 bl[439] br[439] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_440 bl[440] br[440] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_441 bl[441] br[441] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_442 bl[442] br[442] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_443 bl[443] br[443] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_444 bl[444] br[444] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_445 bl[445] br[445] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_446 bl[446] br[446] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_447 bl[447] br[447] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_448 bl[448] br[448] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_449 bl[449] br[449] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_450 bl[450] br[450] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_451 bl[451] br[451] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_452 bl[452] br[452] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_453 bl[453] br[453] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_454 bl[454] br[454] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_455 bl[455] br[455] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_456 bl[456] br[456] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_457 bl[457] br[457] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_458 bl[458] br[458] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_459 bl[459] br[459] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_460 bl[460] br[460] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_461 bl[461] br[461] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_462 bl[462] br[462] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_463 bl[463] br[463] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_464 bl[464] br[464] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_465 bl[465] br[465] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_466 bl[466] br[466] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_467 bl[467] br[467] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_468 bl[468] br[468] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_469 bl[469] br[469] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_470 bl[470] br[470] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_471 bl[471] br[471] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_472 bl[472] br[472] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_473 bl[473] br[473] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_474 bl[474] br[474] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_475 bl[475] br[475] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_476 bl[476] br[476] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_477 bl[477] br[477] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_478 bl[478] br[478] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_479 bl[479] br[479] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_480 bl[480] br[480] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_481 bl[481] br[481] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_482 bl[482] br[482] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_483 bl[483] br[483] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_484 bl[484] br[484] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_485 bl[485] br[485] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_486 bl[486] br[486] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_487 bl[487] br[487] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_488 bl[488] br[488] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_489 bl[489] br[489] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_490 bl[490] br[490] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_491 bl[491] br[491] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_492 bl[492] br[492] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_493 bl[493] br[493] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_494 bl[494] br[494] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_495 bl[495] br[495] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_496 bl[496] br[496] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_497 bl[497] br[497] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_498 bl[498] br[498] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_499 bl[499] br[499] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_500 bl[500] br[500] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_501 bl[501] br[501] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_502 bl[502] br[502] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_503 bl[503] br[503] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_504 bl[504] br[504] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_505 bl[505] br[505] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_506 bl[506] br[506] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_507 bl[507] br[507] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_508 bl[508] br[508] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_509 bl[509] br[509] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_510 bl[510] br[510] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_42_511 bl[511] br[511] vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xcell_43_0 bl[0] br[0] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_1 bl[1] br[1] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_2 bl[2] br[2] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_3 bl[3] br[3] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_4 bl[4] br[4] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_5 bl[5] br[5] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_6 bl[6] br[6] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_7 bl[7] br[7] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_8 bl[8] br[8] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_9 bl[9] br[9] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_10 bl[10] br[10] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_11 bl[11] br[11] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_12 bl[12] br[12] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_13 bl[13] br[13] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_14 bl[14] br[14] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_15 bl[15] br[15] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_16 bl[16] br[16] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_17 bl[17] br[17] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_18 bl[18] br[18] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_19 bl[19] br[19] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_20 bl[20] br[20] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_21 bl[21] br[21] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_22 bl[22] br[22] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_23 bl[23] br[23] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_24 bl[24] br[24] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_25 bl[25] br[25] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_26 bl[26] br[26] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_27 bl[27] br[27] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_28 bl[28] br[28] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_29 bl[29] br[29] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_30 bl[30] br[30] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_31 bl[31] br[31] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_32 bl[32] br[32] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_33 bl[33] br[33] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_34 bl[34] br[34] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_35 bl[35] br[35] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_36 bl[36] br[36] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_37 bl[37] br[37] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_38 bl[38] br[38] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_39 bl[39] br[39] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_40 bl[40] br[40] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_41 bl[41] br[41] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_42 bl[42] br[42] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_43 bl[43] br[43] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_44 bl[44] br[44] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_45 bl[45] br[45] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_46 bl[46] br[46] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_47 bl[47] br[47] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_48 bl[48] br[48] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_49 bl[49] br[49] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_50 bl[50] br[50] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_51 bl[51] br[51] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_52 bl[52] br[52] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_53 bl[53] br[53] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_54 bl[54] br[54] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_55 bl[55] br[55] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_56 bl[56] br[56] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_57 bl[57] br[57] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_58 bl[58] br[58] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_59 bl[59] br[59] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_60 bl[60] br[60] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_61 bl[61] br[61] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_62 bl[62] br[62] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_63 bl[63] br[63] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_64 bl[64] br[64] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_65 bl[65] br[65] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_66 bl[66] br[66] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_67 bl[67] br[67] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_68 bl[68] br[68] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_69 bl[69] br[69] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_70 bl[70] br[70] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_71 bl[71] br[71] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_72 bl[72] br[72] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_73 bl[73] br[73] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_74 bl[74] br[74] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_75 bl[75] br[75] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_76 bl[76] br[76] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_77 bl[77] br[77] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_78 bl[78] br[78] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_79 bl[79] br[79] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_80 bl[80] br[80] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_81 bl[81] br[81] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_82 bl[82] br[82] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_83 bl[83] br[83] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_84 bl[84] br[84] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_85 bl[85] br[85] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_86 bl[86] br[86] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_87 bl[87] br[87] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_88 bl[88] br[88] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_89 bl[89] br[89] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_90 bl[90] br[90] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_91 bl[91] br[91] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_92 bl[92] br[92] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_93 bl[93] br[93] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_94 bl[94] br[94] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_95 bl[95] br[95] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_96 bl[96] br[96] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_97 bl[97] br[97] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_98 bl[98] br[98] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_99 bl[99] br[99] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_100 bl[100] br[100] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_101 bl[101] br[101] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_102 bl[102] br[102] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_103 bl[103] br[103] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_104 bl[104] br[104] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_105 bl[105] br[105] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_106 bl[106] br[106] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_107 bl[107] br[107] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_108 bl[108] br[108] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_109 bl[109] br[109] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_110 bl[110] br[110] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_111 bl[111] br[111] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_112 bl[112] br[112] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_113 bl[113] br[113] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_114 bl[114] br[114] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_115 bl[115] br[115] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_116 bl[116] br[116] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_117 bl[117] br[117] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_118 bl[118] br[118] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_119 bl[119] br[119] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_120 bl[120] br[120] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_121 bl[121] br[121] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_122 bl[122] br[122] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_123 bl[123] br[123] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_124 bl[124] br[124] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_125 bl[125] br[125] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_126 bl[126] br[126] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_127 bl[127] br[127] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_128 bl[128] br[128] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_129 bl[129] br[129] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_130 bl[130] br[130] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_131 bl[131] br[131] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_132 bl[132] br[132] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_133 bl[133] br[133] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_134 bl[134] br[134] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_135 bl[135] br[135] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_136 bl[136] br[136] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_137 bl[137] br[137] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_138 bl[138] br[138] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_139 bl[139] br[139] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_140 bl[140] br[140] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_141 bl[141] br[141] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_142 bl[142] br[142] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_143 bl[143] br[143] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_144 bl[144] br[144] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_145 bl[145] br[145] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_146 bl[146] br[146] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_147 bl[147] br[147] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_148 bl[148] br[148] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_149 bl[149] br[149] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_150 bl[150] br[150] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_151 bl[151] br[151] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_152 bl[152] br[152] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_153 bl[153] br[153] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_154 bl[154] br[154] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_155 bl[155] br[155] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_156 bl[156] br[156] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_157 bl[157] br[157] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_158 bl[158] br[158] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_159 bl[159] br[159] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_160 bl[160] br[160] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_161 bl[161] br[161] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_162 bl[162] br[162] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_163 bl[163] br[163] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_164 bl[164] br[164] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_165 bl[165] br[165] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_166 bl[166] br[166] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_167 bl[167] br[167] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_168 bl[168] br[168] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_169 bl[169] br[169] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_170 bl[170] br[170] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_171 bl[171] br[171] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_172 bl[172] br[172] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_173 bl[173] br[173] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_174 bl[174] br[174] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_175 bl[175] br[175] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_176 bl[176] br[176] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_177 bl[177] br[177] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_178 bl[178] br[178] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_179 bl[179] br[179] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_180 bl[180] br[180] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_181 bl[181] br[181] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_182 bl[182] br[182] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_183 bl[183] br[183] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_184 bl[184] br[184] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_185 bl[185] br[185] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_186 bl[186] br[186] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_187 bl[187] br[187] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_188 bl[188] br[188] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_189 bl[189] br[189] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_190 bl[190] br[190] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_191 bl[191] br[191] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_192 bl[192] br[192] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_193 bl[193] br[193] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_194 bl[194] br[194] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_195 bl[195] br[195] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_196 bl[196] br[196] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_197 bl[197] br[197] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_198 bl[198] br[198] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_199 bl[199] br[199] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_200 bl[200] br[200] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_201 bl[201] br[201] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_202 bl[202] br[202] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_203 bl[203] br[203] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_204 bl[204] br[204] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_205 bl[205] br[205] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_206 bl[206] br[206] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_207 bl[207] br[207] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_208 bl[208] br[208] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_209 bl[209] br[209] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_210 bl[210] br[210] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_211 bl[211] br[211] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_212 bl[212] br[212] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_213 bl[213] br[213] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_214 bl[214] br[214] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_215 bl[215] br[215] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_216 bl[216] br[216] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_217 bl[217] br[217] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_218 bl[218] br[218] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_219 bl[219] br[219] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_220 bl[220] br[220] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_221 bl[221] br[221] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_222 bl[222] br[222] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_223 bl[223] br[223] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_224 bl[224] br[224] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_225 bl[225] br[225] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_226 bl[226] br[226] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_227 bl[227] br[227] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_228 bl[228] br[228] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_229 bl[229] br[229] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_230 bl[230] br[230] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_231 bl[231] br[231] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_232 bl[232] br[232] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_233 bl[233] br[233] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_234 bl[234] br[234] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_235 bl[235] br[235] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_236 bl[236] br[236] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_237 bl[237] br[237] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_238 bl[238] br[238] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_239 bl[239] br[239] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_240 bl[240] br[240] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_241 bl[241] br[241] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_242 bl[242] br[242] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_243 bl[243] br[243] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_244 bl[244] br[244] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_245 bl[245] br[245] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_246 bl[246] br[246] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_247 bl[247] br[247] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_248 bl[248] br[248] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_249 bl[249] br[249] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_250 bl[250] br[250] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_251 bl[251] br[251] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_252 bl[252] br[252] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_253 bl[253] br[253] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_254 bl[254] br[254] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_255 bl[255] br[255] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_256 bl[256] br[256] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_257 bl[257] br[257] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_258 bl[258] br[258] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_259 bl[259] br[259] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_260 bl[260] br[260] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_261 bl[261] br[261] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_262 bl[262] br[262] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_263 bl[263] br[263] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_264 bl[264] br[264] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_265 bl[265] br[265] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_266 bl[266] br[266] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_267 bl[267] br[267] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_268 bl[268] br[268] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_269 bl[269] br[269] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_270 bl[270] br[270] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_271 bl[271] br[271] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_272 bl[272] br[272] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_273 bl[273] br[273] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_274 bl[274] br[274] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_275 bl[275] br[275] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_276 bl[276] br[276] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_277 bl[277] br[277] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_278 bl[278] br[278] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_279 bl[279] br[279] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_280 bl[280] br[280] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_281 bl[281] br[281] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_282 bl[282] br[282] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_283 bl[283] br[283] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_284 bl[284] br[284] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_285 bl[285] br[285] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_286 bl[286] br[286] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_287 bl[287] br[287] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_288 bl[288] br[288] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_289 bl[289] br[289] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_290 bl[290] br[290] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_291 bl[291] br[291] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_292 bl[292] br[292] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_293 bl[293] br[293] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_294 bl[294] br[294] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_295 bl[295] br[295] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_296 bl[296] br[296] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_297 bl[297] br[297] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_298 bl[298] br[298] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_299 bl[299] br[299] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_300 bl[300] br[300] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_301 bl[301] br[301] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_302 bl[302] br[302] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_303 bl[303] br[303] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_304 bl[304] br[304] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_305 bl[305] br[305] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_306 bl[306] br[306] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_307 bl[307] br[307] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_308 bl[308] br[308] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_309 bl[309] br[309] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_310 bl[310] br[310] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_311 bl[311] br[311] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_312 bl[312] br[312] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_313 bl[313] br[313] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_314 bl[314] br[314] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_315 bl[315] br[315] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_316 bl[316] br[316] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_317 bl[317] br[317] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_318 bl[318] br[318] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_319 bl[319] br[319] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_320 bl[320] br[320] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_321 bl[321] br[321] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_322 bl[322] br[322] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_323 bl[323] br[323] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_324 bl[324] br[324] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_325 bl[325] br[325] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_326 bl[326] br[326] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_327 bl[327] br[327] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_328 bl[328] br[328] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_329 bl[329] br[329] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_330 bl[330] br[330] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_331 bl[331] br[331] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_332 bl[332] br[332] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_333 bl[333] br[333] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_334 bl[334] br[334] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_335 bl[335] br[335] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_336 bl[336] br[336] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_337 bl[337] br[337] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_338 bl[338] br[338] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_339 bl[339] br[339] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_340 bl[340] br[340] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_341 bl[341] br[341] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_342 bl[342] br[342] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_343 bl[343] br[343] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_344 bl[344] br[344] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_345 bl[345] br[345] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_346 bl[346] br[346] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_347 bl[347] br[347] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_348 bl[348] br[348] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_349 bl[349] br[349] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_350 bl[350] br[350] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_351 bl[351] br[351] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_352 bl[352] br[352] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_353 bl[353] br[353] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_354 bl[354] br[354] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_355 bl[355] br[355] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_356 bl[356] br[356] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_357 bl[357] br[357] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_358 bl[358] br[358] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_359 bl[359] br[359] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_360 bl[360] br[360] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_361 bl[361] br[361] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_362 bl[362] br[362] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_363 bl[363] br[363] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_364 bl[364] br[364] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_365 bl[365] br[365] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_366 bl[366] br[366] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_367 bl[367] br[367] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_368 bl[368] br[368] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_369 bl[369] br[369] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_370 bl[370] br[370] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_371 bl[371] br[371] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_372 bl[372] br[372] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_373 bl[373] br[373] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_374 bl[374] br[374] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_375 bl[375] br[375] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_376 bl[376] br[376] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_377 bl[377] br[377] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_378 bl[378] br[378] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_379 bl[379] br[379] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_380 bl[380] br[380] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_381 bl[381] br[381] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_382 bl[382] br[382] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_383 bl[383] br[383] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_384 bl[384] br[384] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_385 bl[385] br[385] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_386 bl[386] br[386] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_387 bl[387] br[387] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_388 bl[388] br[388] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_389 bl[389] br[389] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_390 bl[390] br[390] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_391 bl[391] br[391] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_392 bl[392] br[392] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_393 bl[393] br[393] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_394 bl[394] br[394] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_395 bl[395] br[395] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_396 bl[396] br[396] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_397 bl[397] br[397] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_398 bl[398] br[398] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_399 bl[399] br[399] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_400 bl[400] br[400] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_401 bl[401] br[401] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_402 bl[402] br[402] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_403 bl[403] br[403] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_404 bl[404] br[404] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_405 bl[405] br[405] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_406 bl[406] br[406] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_407 bl[407] br[407] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_408 bl[408] br[408] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_409 bl[409] br[409] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_410 bl[410] br[410] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_411 bl[411] br[411] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_412 bl[412] br[412] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_413 bl[413] br[413] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_414 bl[414] br[414] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_415 bl[415] br[415] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_416 bl[416] br[416] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_417 bl[417] br[417] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_418 bl[418] br[418] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_419 bl[419] br[419] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_420 bl[420] br[420] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_421 bl[421] br[421] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_422 bl[422] br[422] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_423 bl[423] br[423] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_424 bl[424] br[424] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_425 bl[425] br[425] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_426 bl[426] br[426] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_427 bl[427] br[427] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_428 bl[428] br[428] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_429 bl[429] br[429] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_430 bl[430] br[430] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_431 bl[431] br[431] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_432 bl[432] br[432] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_433 bl[433] br[433] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_434 bl[434] br[434] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_435 bl[435] br[435] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_436 bl[436] br[436] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_437 bl[437] br[437] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_438 bl[438] br[438] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_439 bl[439] br[439] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_440 bl[440] br[440] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_441 bl[441] br[441] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_442 bl[442] br[442] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_443 bl[443] br[443] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_444 bl[444] br[444] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_445 bl[445] br[445] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_446 bl[446] br[446] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_447 bl[447] br[447] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_448 bl[448] br[448] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_449 bl[449] br[449] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_450 bl[450] br[450] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_451 bl[451] br[451] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_452 bl[452] br[452] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_453 bl[453] br[453] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_454 bl[454] br[454] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_455 bl[455] br[455] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_456 bl[456] br[456] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_457 bl[457] br[457] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_458 bl[458] br[458] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_459 bl[459] br[459] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_460 bl[460] br[460] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_461 bl[461] br[461] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_462 bl[462] br[462] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_463 bl[463] br[463] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_464 bl[464] br[464] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_465 bl[465] br[465] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_466 bl[466] br[466] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_467 bl[467] br[467] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_468 bl[468] br[468] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_469 bl[469] br[469] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_470 bl[470] br[470] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_471 bl[471] br[471] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_472 bl[472] br[472] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_473 bl[473] br[473] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_474 bl[474] br[474] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_475 bl[475] br[475] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_476 bl[476] br[476] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_477 bl[477] br[477] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_478 bl[478] br[478] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_479 bl[479] br[479] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_480 bl[480] br[480] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_481 bl[481] br[481] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_482 bl[482] br[482] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_483 bl[483] br[483] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_484 bl[484] br[484] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_485 bl[485] br[485] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_486 bl[486] br[486] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_487 bl[487] br[487] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_488 bl[488] br[488] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_489 bl[489] br[489] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_490 bl[490] br[490] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_491 bl[491] br[491] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_492 bl[492] br[492] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_493 bl[493] br[493] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_494 bl[494] br[494] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_495 bl[495] br[495] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_496 bl[496] br[496] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_497 bl[497] br[497] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_498 bl[498] br[498] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_499 bl[499] br[499] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_500 bl[500] br[500] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_501 bl[501] br[501] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_502 bl[502] br[502] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_503 bl[503] br[503] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_504 bl[504] br[504] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_505 bl[505] br[505] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_506 bl[506] br[506] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_507 bl[507] br[507] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_508 bl[508] br[508] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_509 bl[509] br[509] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_510 bl[510] br[510] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_43_511 bl[511] br[511] vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xcell_44_0 bl[0] br[0] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_1 bl[1] br[1] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_2 bl[2] br[2] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_3 bl[3] br[3] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_4 bl[4] br[4] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_5 bl[5] br[5] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_6 bl[6] br[6] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_7 bl[7] br[7] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_8 bl[8] br[8] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_9 bl[9] br[9] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_10 bl[10] br[10] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_11 bl[11] br[11] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_12 bl[12] br[12] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_13 bl[13] br[13] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_14 bl[14] br[14] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_15 bl[15] br[15] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_16 bl[16] br[16] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_17 bl[17] br[17] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_18 bl[18] br[18] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_19 bl[19] br[19] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_20 bl[20] br[20] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_21 bl[21] br[21] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_22 bl[22] br[22] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_23 bl[23] br[23] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_24 bl[24] br[24] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_25 bl[25] br[25] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_26 bl[26] br[26] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_27 bl[27] br[27] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_28 bl[28] br[28] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_29 bl[29] br[29] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_30 bl[30] br[30] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_31 bl[31] br[31] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_32 bl[32] br[32] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_33 bl[33] br[33] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_34 bl[34] br[34] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_35 bl[35] br[35] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_36 bl[36] br[36] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_37 bl[37] br[37] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_38 bl[38] br[38] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_39 bl[39] br[39] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_40 bl[40] br[40] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_41 bl[41] br[41] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_42 bl[42] br[42] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_43 bl[43] br[43] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_44 bl[44] br[44] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_45 bl[45] br[45] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_46 bl[46] br[46] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_47 bl[47] br[47] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_48 bl[48] br[48] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_49 bl[49] br[49] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_50 bl[50] br[50] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_51 bl[51] br[51] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_52 bl[52] br[52] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_53 bl[53] br[53] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_54 bl[54] br[54] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_55 bl[55] br[55] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_56 bl[56] br[56] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_57 bl[57] br[57] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_58 bl[58] br[58] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_59 bl[59] br[59] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_60 bl[60] br[60] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_61 bl[61] br[61] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_62 bl[62] br[62] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_63 bl[63] br[63] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_64 bl[64] br[64] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_65 bl[65] br[65] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_66 bl[66] br[66] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_67 bl[67] br[67] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_68 bl[68] br[68] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_69 bl[69] br[69] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_70 bl[70] br[70] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_71 bl[71] br[71] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_72 bl[72] br[72] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_73 bl[73] br[73] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_74 bl[74] br[74] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_75 bl[75] br[75] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_76 bl[76] br[76] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_77 bl[77] br[77] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_78 bl[78] br[78] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_79 bl[79] br[79] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_80 bl[80] br[80] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_81 bl[81] br[81] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_82 bl[82] br[82] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_83 bl[83] br[83] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_84 bl[84] br[84] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_85 bl[85] br[85] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_86 bl[86] br[86] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_87 bl[87] br[87] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_88 bl[88] br[88] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_89 bl[89] br[89] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_90 bl[90] br[90] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_91 bl[91] br[91] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_92 bl[92] br[92] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_93 bl[93] br[93] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_94 bl[94] br[94] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_95 bl[95] br[95] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_96 bl[96] br[96] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_97 bl[97] br[97] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_98 bl[98] br[98] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_99 bl[99] br[99] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_100 bl[100] br[100] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_101 bl[101] br[101] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_102 bl[102] br[102] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_103 bl[103] br[103] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_104 bl[104] br[104] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_105 bl[105] br[105] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_106 bl[106] br[106] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_107 bl[107] br[107] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_108 bl[108] br[108] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_109 bl[109] br[109] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_110 bl[110] br[110] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_111 bl[111] br[111] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_112 bl[112] br[112] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_113 bl[113] br[113] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_114 bl[114] br[114] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_115 bl[115] br[115] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_116 bl[116] br[116] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_117 bl[117] br[117] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_118 bl[118] br[118] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_119 bl[119] br[119] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_120 bl[120] br[120] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_121 bl[121] br[121] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_122 bl[122] br[122] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_123 bl[123] br[123] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_124 bl[124] br[124] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_125 bl[125] br[125] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_126 bl[126] br[126] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_127 bl[127] br[127] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_128 bl[128] br[128] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_129 bl[129] br[129] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_130 bl[130] br[130] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_131 bl[131] br[131] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_132 bl[132] br[132] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_133 bl[133] br[133] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_134 bl[134] br[134] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_135 bl[135] br[135] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_136 bl[136] br[136] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_137 bl[137] br[137] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_138 bl[138] br[138] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_139 bl[139] br[139] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_140 bl[140] br[140] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_141 bl[141] br[141] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_142 bl[142] br[142] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_143 bl[143] br[143] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_144 bl[144] br[144] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_145 bl[145] br[145] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_146 bl[146] br[146] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_147 bl[147] br[147] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_148 bl[148] br[148] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_149 bl[149] br[149] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_150 bl[150] br[150] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_151 bl[151] br[151] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_152 bl[152] br[152] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_153 bl[153] br[153] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_154 bl[154] br[154] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_155 bl[155] br[155] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_156 bl[156] br[156] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_157 bl[157] br[157] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_158 bl[158] br[158] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_159 bl[159] br[159] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_160 bl[160] br[160] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_161 bl[161] br[161] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_162 bl[162] br[162] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_163 bl[163] br[163] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_164 bl[164] br[164] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_165 bl[165] br[165] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_166 bl[166] br[166] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_167 bl[167] br[167] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_168 bl[168] br[168] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_169 bl[169] br[169] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_170 bl[170] br[170] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_171 bl[171] br[171] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_172 bl[172] br[172] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_173 bl[173] br[173] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_174 bl[174] br[174] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_175 bl[175] br[175] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_176 bl[176] br[176] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_177 bl[177] br[177] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_178 bl[178] br[178] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_179 bl[179] br[179] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_180 bl[180] br[180] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_181 bl[181] br[181] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_182 bl[182] br[182] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_183 bl[183] br[183] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_184 bl[184] br[184] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_185 bl[185] br[185] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_186 bl[186] br[186] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_187 bl[187] br[187] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_188 bl[188] br[188] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_189 bl[189] br[189] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_190 bl[190] br[190] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_191 bl[191] br[191] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_192 bl[192] br[192] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_193 bl[193] br[193] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_194 bl[194] br[194] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_195 bl[195] br[195] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_196 bl[196] br[196] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_197 bl[197] br[197] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_198 bl[198] br[198] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_199 bl[199] br[199] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_200 bl[200] br[200] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_201 bl[201] br[201] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_202 bl[202] br[202] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_203 bl[203] br[203] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_204 bl[204] br[204] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_205 bl[205] br[205] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_206 bl[206] br[206] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_207 bl[207] br[207] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_208 bl[208] br[208] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_209 bl[209] br[209] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_210 bl[210] br[210] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_211 bl[211] br[211] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_212 bl[212] br[212] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_213 bl[213] br[213] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_214 bl[214] br[214] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_215 bl[215] br[215] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_216 bl[216] br[216] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_217 bl[217] br[217] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_218 bl[218] br[218] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_219 bl[219] br[219] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_220 bl[220] br[220] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_221 bl[221] br[221] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_222 bl[222] br[222] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_223 bl[223] br[223] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_224 bl[224] br[224] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_225 bl[225] br[225] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_226 bl[226] br[226] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_227 bl[227] br[227] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_228 bl[228] br[228] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_229 bl[229] br[229] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_230 bl[230] br[230] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_231 bl[231] br[231] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_232 bl[232] br[232] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_233 bl[233] br[233] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_234 bl[234] br[234] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_235 bl[235] br[235] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_236 bl[236] br[236] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_237 bl[237] br[237] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_238 bl[238] br[238] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_239 bl[239] br[239] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_240 bl[240] br[240] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_241 bl[241] br[241] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_242 bl[242] br[242] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_243 bl[243] br[243] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_244 bl[244] br[244] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_245 bl[245] br[245] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_246 bl[246] br[246] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_247 bl[247] br[247] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_248 bl[248] br[248] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_249 bl[249] br[249] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_250 bl[250] br[250] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_251 bl[251] br[251] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_252 bl[252] br[252] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_253 bl[253] br[253] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_254 bl[254] br[254] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_255 bl[255] br[255] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_256 bl[256] br[256] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_257 bl[257] br[257] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_258 bl[258] br[258] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_259 bl[259] br[259] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_260 bl[260] br[260] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_261 bl[261] br[261] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_262 bl[262] br[262] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_263 bl[263] br[263] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_264 bl[264] br[264] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_265 bl[265] br[265] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_266 bl[266] br[266] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_267 bl[267] br[267] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_268 bl[268] br[268] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_269 bl[269] br[269] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_270 bl[270] br[270] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_271 bl[271] br[271] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_272 bl[272] br[272] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_273 bl[273] br[273] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_274 bl[274] br[274] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_275 bl[275] br[275] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_276 bl[276] br[276] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_277 bl[277] br[277] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_278 bl[278] br[278] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_279 bl[279] br[279] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_280 bl[280] br[280] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_281 bl[281] br[281] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_282 bl[282] br[282] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_283 bl[283] br[283] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_284 bl[284] br[284] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_285 bl[285] br[285] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_286 bl[286] br[286] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_287 bl[287] br[287] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_288 bl[288] br[288] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_289 bl[289] br[289] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_290 bl[290] br[290] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_291 bl[291] br[291] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_292 bl[292] br[292] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_293 bl[293] br[293] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_294 bl[294] br[294] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_295 bl[295] br[295] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_296 bl[296] br[296] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_297 bl[297] br[297] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_298 bl[298] br[298] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_299 bl[299] br[299] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_300 bl[300] br[300] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_301 bl[301] br[301] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_302 bl[302] br[302] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_303 bl[303] br[303] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_304 bl[304] br[304] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_305 bl[305] br[305] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_306 bl[306] br[306] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_307 bl[307] br[307] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_308 bl[308] br[308] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_309 bl[309] br[309] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_310 bl[310] br[310] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_311 bl[311] br[311] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_312 bl[312] br[312] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_313 bl[313] br[313] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_314 bl[314] br[314] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_315 bl[315] br[315] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_316 bl[316] br[316] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_317 bl[317] br[317] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_318 bl[318] br[318] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_319 bl[319] br[319] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_320 bl[320] br[320] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_321 bl[321] br[321] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_322 bl[322] br[322] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_323 bl[323] br[323] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_324 bl[324] br[324] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_325 bl[325] br[325] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_326 bl[326] br[326] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_327 bl[327] br[327] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_328 bl[328] br[328] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_329 bl[329] br[329] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_330 bl[330] br[330] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_331 bl[331] br[331] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_332 bl[332] br[332] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_333 bl[333] br[333] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_334 bl[334] br[334] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_335 bl[335] br[335] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_336 bl[336] br[336] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_337 bl[337] br[337] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_338 bl[338] br[338] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_339 bl[339] br[339] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_340 bl[340] br[340] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_341 bl[341] br[341] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_342 bl[342] br[342] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_343 bl[343] br[343] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_344 bl[344] br[344] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_345 bl[345] br[345] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_346 bl[346] br[346] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_347 bl[347] br[347] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_348 bl[348] br[348] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_349 bl[349] br[349] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_350 bl[350] br[350] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_351 bl[351] br[351] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_352 bl[352] br[352] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_353 bl[353] br[353] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_354 bl[354] br[354] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_355 bl[355] br[355] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_356 bl[356] br[356] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_357 bl[357] br[357] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_358 bl[358] br[358] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_359 bl[359] br[359] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_360 bl[360] br[360] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_361 bl[361] br[361] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_362 bl[362] br[362] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_363 bl[363] br[363] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_364 bl[364] br[364] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_365 bl[365] br[365] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_366 bl[366] br[366] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_367 bl[367] br[367] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_368 bl[368] br[368] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_369 bl[369] br[369] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_370 bl[370] br[370] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_371 bl[371] br[371] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_372 bl[372] br[372] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_373 bl[373] br[373] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_374 bl[374] br[374] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_375 bl[375] br[375] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_376 bl[376] br[376] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_377 bl[377] br[377] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_378 bl[378] br[378] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_379 bl[379] br[379] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_380 bl[380] br[380] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_381 bl[381] br[381] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_382 bl[382] br[382] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_383 bl[383] br[383] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_384 bl[384] br[384] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_385 bl[385] br[385] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_386 bl[386] br[386] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_387 bl[387] br[387] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_388 bl[388] br[388] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_389 bl[389] br[389] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_390 bl[390] br[390] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_391 bl[391] br[391] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_392 bl[392] br[392] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_393 bl[393] br[393] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_394 bl[394] br[394] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_395 bl[395] br[395] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_396 bl[396] br[396] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_397 bl[397] br[397] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_398 bl[398] br[398] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_399 bl[399] br[399] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_400 bl[400] br[400] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_401 bl[401] br[401] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_402 bl[402] br[402] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_403 bl[403] br[403] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_404 bl[404] br[404] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_405 bl[405] br[405] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_406 bl[406] br[406] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_407 bl[407] br[407] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_408 bl[408] br[408] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_409 bl[409] br[409] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_410 bl[410] br[410] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_411 bl[411] br[411] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_412 bl[412] br[412] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_413 bl[413] br[413] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_414 bl[414] br[414] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_415 bl[415] br[415] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_416 bl[416] br[416] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_417 bl[417] br[417] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_418 bl[418] br[418] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_419 bl[419] br[419] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_420 bl[420] br[420] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_421 bl[421] br[421] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_422 bl[422] br[422] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_423 bl[423] br[423] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_424 bl[424] br[424] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_425 bl[425] br[425] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_426 bl[426] br[426] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_427 bl[427] br[427] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_428 bl[428] br[428] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_429 bl[429] br[429] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_430 bl[430] br[430] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_431 bl[431] br[431] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_432 bl[432] br[432] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_433 bl[433] br[433] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_434 bl[434] br[434] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_435 bl[435] br[435] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_436 bl[436] br[436] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_437 bl[437] br[437] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_438 bl[438] br[438] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_439 bl[439] br[439] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_440 bl[440] br[440] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_441 bl[441] br[441] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_442 bl[442] br[442] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_443 bl[443] br[443] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_444 bl[444] br[444] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_445 bl[445] br[445] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_446 bl[446] br[446] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_447 bl[447] br[447] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_448 bl[448] br[448] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_449 bl[449] br[449] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_450 bl[450] br[450] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_451 bl[451] br[451] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_452 bl[452] br[452] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_453 bl[453] br[453] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_454 bl[454] br[454] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_455 bl[455] br[455] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_456 bl[456] br[456] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_457 bl[457] br[457] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_458 bl[458] br[458] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_459 bl[459] br[459] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_460 bl[460] br[460] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_461 bl[461] br[461] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_462 bl[462] br[462] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_463 bl[463] br[463] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_464 bl[464] br[464] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_465 bl[465] br[465] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_466 bl[466] br[466] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_467 bl[467] br[467] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_468 bl[468] br[468] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_469 bl[469] br[469] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_470 bl[470] br[470] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_471 bl[471] br[471] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_472 bl[472] br[472] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_473 bl[473] br[473] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_474 bl[474] br[474] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_475 bl[475] br[475] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_476 bl[476] br[476] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_477 bl[477] br[477] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_478 bl[478] br[478] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_479 bl[479] br[479] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_480 bl[480] br[480] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_481 bl[481] br[481] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_482 bl[482] br[482] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_483 bl[483] br[483] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_484 bl[484] br[484] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_485 bl[485] br[485] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_486 bl[486] br[486] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_487 bl[487] br[487] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_488 bl[488] br[488] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_489 bl[489] br[489] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_490 bl[490] br[490] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_491 bl[491] br[491] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_492 bl[492] br[492] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_493 bl[493] br[493] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_494 bl[494] br[494] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_495 bl[495] br[495] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_496 bl[496] br[496] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_497 bl[497] br[497] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_498 bl[498] br[498] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_499 bl[499] br[499] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_500 bl[500] br[500] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_501 bl[501] br[501] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_502 bl[502] br[502] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_503 bl[503] br[503] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_504 bl[504] br[504] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_505 bl[505] br[505] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_506 bl[506] br[506] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_507 bl[507] br[507] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_508 bl[508] br[508] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_509 bl[509] br[509] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_510 bl[510] br[510] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_44_511 bl[511] br[511] vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xcell_45_0 bl[0] br[0] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_1 bl[1] br[1] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_2 bl[2] br[2] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_3 bl[3] br[3] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_4 bl[4] br[4] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_5 bl[5] br[5] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_6 bl[6] br[6] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_7 bl[7] br[7] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_8 bl[8] br[8] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_9 bl[9] br[9] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_10 bl[10] br[10] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_11 bl[11] br[11] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_12 bl[12] br[12] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_13 bl[13] br[13] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_14 bl[14] br[14] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_15 bl[15] br[15] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_16 bl[16] br[16] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_17 bl[17] br[17] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_18 bl[18] br[18] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_19 bl[19] br[19] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_20 bl[20] br[20] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_21 bl[21] br[21] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_22 bl[22] br[22] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_23 bl[23] br[23] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_24 bl[24] br[24] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_25 bl[25] br[25] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_26 bl[26] br[26] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_27 bl[27] br[27] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_28 bl[28] br[28] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_29 bl[29] br[29] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_30 bl[30] br[30] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_31 bl[31] br[31] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_32 bl[32] br[32] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_33 bl[33] br[33] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_34 bl[34] br[34] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_35 bl[35] br[35] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_36 bl[36] br[36] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_37 bl[37] br[37] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_38 bl[38] br[38] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_39 bl[39] br[39] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_40 bl[40] br[40] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_41 bl[41] br[41] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_42 bl[42] br[42] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_43 bl[43] br[43] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_44 bl[44] br[44] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_45 bl[45] br[45] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_46 bl[46] br[46] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_47 bl[47] br[47] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_48 bl[48] br[48] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_49 bl[49] br[49] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_50 bl[50] br[50] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_51 bl[51] br[51] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_52 bl[52] br[52] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_53 bl[53] br[53] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_54 bl[54] br[54] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_55 bl[55] br[55] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_56 bl[56] br[56] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_57 bl[57] br[57] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_58 bl[58] br[58] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_59 bl[59] br[59] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_60 bl[60] br[60] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_61 bl[61] br[61] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_62 bl[62] br[62] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_63 bl[63] br[63] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_64 bl[64] br[64] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_65 bl[65] br[65] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_66 bl[66] br[66] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_67 bl[67] br[67] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_68 bl[68] br[68] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_69 bl[69] br[69] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_70 bl[70] br[70] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_71 bl[71] br[71] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_72 bl[72] br[72] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_73 bl[73] br[73] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_74 bl[74] br[74] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_75 bl[75] br[75] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_76 bl[76] br[76] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_77 bl[77] br[77] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_78 bl[78] br[78] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_79 bl[79] br[79] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_80 bl[80] br[80] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_81 bl[81] br[81] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_82 bl[82] br[82] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_83 bl[83] br[83] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_84 bl[84] br[84] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_85 bl[85] br[85] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_86 bl[86] br[86] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_87 bl[87] br[87] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_88 bl[88] br[88] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_89 bl[89] br[89] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_90 bl[90] br[90] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_91 bl[91] br[91] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_92 bl[92] br[92] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_93 bl[93] br[93] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_94 bl[94] br[94] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_95 bl[95] br[95] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_96 bl[96] br[96] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_97 bl[97] br[97] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_98 bl[98] br[98] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_99 bl[99] br[99] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_100 bl[100] br[100] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_101 bl[101] br[101] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_102 bl[102] br[102] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_103 bl[103] br[103] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_104 bl[104] br[104] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_105 bl[105] br[105] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_106 bl[106] br[106] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_107 bl[107] br[107] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_108 bl[108] br[108] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_109 bl[109] br[109] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_110 bl[110] br[110] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_111 bl[111] br[111] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_112 bl[112] br[112] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_113 bl[113] br[113] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_114 bl[114] br[114] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_115 bl[115] br[115] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_116 bl[116] br[116] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_117 bl[117] br[117] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_118 bl[118] br[118] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_119 bl[119] br[119] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_120 bl[120] br[120] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_121 bl[121] br[121] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_122 bl[122] br[122] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_123 bl[123] br[123] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_124 bl[124] br[124] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_125 bl[125] br[125] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_126 bl[126] br[126] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_127 bl[127] br[127] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_128 bl[128] br[128] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_129 bl[129] br[129] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_130 bl[130] br[130] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_131 bl[131] br[131] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_132 bl[132] br[132] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_133 bl[133] br[133] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_134 bl[134] br[134] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_135 bl[135] br[135] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_136 bl[136] br[136] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_137 bl[137] br[137] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_138 bl[138] br[138] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_139 bl[139] br[139] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_140 bl[140] br[140] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_141 bl[141] br[141] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_142 bl[142] br[142] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_143 bl[143] br[143] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_144 bl[144] br[144] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_145 bl[145] br[145] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_146 bl[146] br[146] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_147 bl[147] br[147] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_148 bl[148] br[148] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_149 bl[149] br[149] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_150 bl[150] br[150] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_151 bl[151] br[151] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_152 bl[152] br[152] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_153 bl[153] br[153] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_154 bl[154] br[154] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_155 bl[155] br[155] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_156 bl[156] br[156] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_157 bl[157] br[157] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_158 bl[158] br[158] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_159 bl[159] br[159] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_160 bl[160] br[160] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_161 bl[161] br[161] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_162 bl[162] br[162] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_163 bl[163] br[163] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_164 bl[164] br[164] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_165 bl[165] br[165] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_166 bl[166] br[166] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_167 bl[167] br[167] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_168 bl[168] br[168] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_169 bl[169] br[169] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_170 bl[170] br[170] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_171 bl[171] br[171] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_172 bl[172] br[172] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_173 bl[173] br[173] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_174 bl[174] br[174] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_175 bl[175] br[175] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_176 bl[176] br[176] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_177 bl[177] br[177] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_178 bl[178] br[178] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_179 bl[179] br[179] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_180 bl[180] br[180] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_181 bl[181] br[181] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_182 bl[182] br[182] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_183 bl[183] br[183] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_184 bl[184] br[184] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_185 bl[185] br[185] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_186 bl[186] br[186] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_187 bl[187] br[187] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_188 bl[188] br[188] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_189 bl[189] br[189] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_190 bl[190] br[190] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_191 bl[191] br[191] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_192 bl[192] br[192] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_193 bl[193] br[193] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_194 bl[194] br[194] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_195 bl[195] br[195] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_196 bl[196] br[196] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_197 bl[197] br[197] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_198 bl[198] br[198] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_199 bl[199] br[199] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_200 bl[200] br[200] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_201 bl[201] br[201] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_202 bl[202] br[202] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_203 bl[203] br[203] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_204 bl[204] br[204] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_205 bl[205] br[205] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_206 bl[206] br[206] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_207 bl[207] br[207] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_208 bl[208] br[208] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_209 bl[209] br[209] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_210 bl[210] br[210] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_211 bl[211] br[211] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_212 bl[212] br[212] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_213 bl[213] br[213] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_214 bl[214] br[214] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_215 bl[215] br[215] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_216 bl[216] br[216] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_217 bl[217] br[217] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_218 bl[218] br[218] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_219 bl[219] br[219] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_220 bl[220] br[220] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_221 bl[221] br[221] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_222 bl[222] br[222] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_223 bl[223] br[223] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_224 bl[224] br[224] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_225 bl[225] br[225] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_226 bl[226] br[226] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_227 bl[227] br[227] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_228 bl[228] br[228] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_229 bl[229] br[229] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_230 bl[230] br[230] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_231 bl[231] br[231] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_232 bl[232] br[232] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_233 bl[233] br[233] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_234 bl[234] br[234] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_235 bl[235] br[235] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_236 bl[236] br[236] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_237 bl[237] br[237] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_238 bl[238] br[238] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_239 bl[239] br[239] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_240 bl[240] br[240] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_241 bl[241] br[241] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_242 bl[242] br[242] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_243 bl[243] br[243] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_244 bl[244] br[244] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_245 bl[245] br[245] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_246 bl[246] br[246] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_247 bl[247] br[247] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_248 bl[248] br[248] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_249 bl[249] br[249] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_250 bl[250] br[250] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_251 bl[251] br[251] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_252 bl[252] br[252] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_253 bl[253] br[253] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_254 bl[254] br[254] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_255 bl[255] br[255] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_256 bl[256] br[256] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_257 bl[257] br[257] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_258 bl[258] br[258] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_259 bl[259] br[259] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_260 bl[260] br[260] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_261 bl[261] br[261] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_262 bl[262] br[262] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_263 bl[263] br[263] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_264 bl[264] br[264] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_265 bl[265] br[265] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_266 bl[266] br[266] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_267 bl[267] br[267] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_268 bl[268] br[268] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_269 bl[269] br[269] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_270 bl[270] br[270] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_271 bl[271] br[271] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_272 bl[272] br[272] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_273 bl[273] br[273] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_274 bl[274] br[274] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_275 bl[275] br[275] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_276 bl[276] br[276] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_277 bl[277] br[277] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_278 bl[278] br[278] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_279 bl[279] br[279] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_280 bl[280] br[280] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_281 bl[281] br[281] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_282 bl[282] br[282] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_283 bl[283] br[283] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_284 bl[284] br[284] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_285 bl[285] br[285] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_286 bl[286] br[286] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_287 bl[287] br[287] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_288 bl[288] br[288] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_289 bl[289] br[289] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_290 bl[290] br[290] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_291 bl[291] br[291] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_292 bl[292] br[292] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_293 bl[293] br[293] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_294 bl[294] br[294] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_295 bl[295] br[295] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_296 bl[296] br[296] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_297 bl[297] br[297] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_298 bl[298] br[298] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_299 bl[299] br[299] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_300 bl[300] br[300] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_301 bl[301] br[301] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_302 bl[302] br[302] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_303 bl[303] br[303] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_304 bl[304] br[304] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_305 bl[305] br[305] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_306 bl[306] br[306] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_307 bl[307] br[307] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_308 bl[308] br[308] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_309 bl[309] br[309] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_310 bl[310] br[310] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_311 bl[311] br[311] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_312 bl[312] br[312] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_313 bl[313] br[313] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_314 bl[314] br[314] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_315 bl[315] br[315] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_316 bl[316] br[316] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_317 bl[317] br[317] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_318 bl[318] br[318] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_319 bl[319] br[319] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_320 bl[320] br[320] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_321 bl[321] br[321] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_322 bl[322] br[322] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_323 bl[323] br[323] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_324 bl[324] br[324] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_325 bl[325] br[325] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_326 bl[326] br[326] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_327 bl[327] br[327] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_328 bl[328] br[328] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_329 bl[329] br[329] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_330 bl[330] br[330] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_331 bl[331] br[331] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_332 bl[332] br[332] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_333 bl[333] br[333] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_334 bl[334] br[334] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_335 bl[335] br[335] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_336 bl[336] br[336] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_337 bl[337] br[337] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_338 bl[338] br[338] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_339 bl[339] br[339] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_340 bl[340] br[340] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_341 bl[341] br[341] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_342 bl[342] br[342] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_343 bl[343] br[343] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_344 bl[344] br[344] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_345 bl[345] br[345] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_346 bl[346] br[346] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_347 bl[347] br[347] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_348 bl[348] br[348] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_349 bl[349] br[349] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_350 bl[350] br[350] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_351 bl[351] br[351] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_352 bl[352] br[352] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_353 bl[353] br[353] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_354 bl[354] br[354] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_355 bl[355] br[355] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_356 bl[356] br[356] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_357 bl[357] br[357] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_358 bl[358] br[358] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_359 bl[359] br[359] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_360 bl[360] br[360] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_361 bl[361] br[361] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_362 bl[362] br[362] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_363 bl[363] br[363] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_364 bl[364] br[364] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_365 bl[365] br[365] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_366 bl[366] br[366] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_367 bl[367] br[367] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_368 bl[368] br[368] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_369 bl[369] br[369] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_370 bl[370] br[370] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_371 bl[371] br[371] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_372 bl[372] br[372] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_373 bl[373] br[373] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_374 bl[374] br[374] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_375 bl[375] br[375] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_376 bl[376] br[376] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_377 bl[377] br[377] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_378 bl[378] br[378] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_379 bl[379] br[379] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_380 bl[380] br[380] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_381 bl[381] br[381] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_382 bl[382] br[382] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_383 bl[383] br[383] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_384 bl[384] br[384] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_385 bl[385] br[385] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_386 bl[386] br[386] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_387 bl[387] br[387] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_388 bl[388] br[388] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_389 bl[389] br[389] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_390 bl[390] br[390] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_391 bl[391] br[391] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_392 bl[392] br[392] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_393 bl[393] br[393] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_394 bl[394] br[394] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_395 bl[395] br[395] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_396 bl[396] br[396] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_397 bl[397] br[397] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_398 bl[398] br[398] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_399 bl[399] br[399] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_400 bl[400] br[400] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_401 bl[401] br[401] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_402 bl[402] br[402] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_403 bl[403] br[403] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_404 bl[404] br[404] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_405 bl[405] br[405] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_406 bl[406] br[406] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_407 bl[407] br[407] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_408 bl[408] br[408] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_409 bl[409] br[409] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_410 bl[410] br[410] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_411 bl[411] br[411] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_412 bl[412] br[412] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_413 bl[413] br[413] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_414 bl[414] br[414] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_415 bl[415] br[415] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_416 bl[416] br[416] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_417 bl[417] br[417] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_418 bl[418] br[418] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_419 bl[419] br[419] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_420 bl[420] br[420] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_421 bl[421] br[421] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_422 bl[422] br[422] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_423 bl[423] br[423] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_424 bl[424] br[424] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_425 bl[425] br[425] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_426 bl[426] br[426] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_427 bl[427] br[427] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_428 bl[428] br[428] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_429 bl[429] br[429] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_430 bl[430] br[430] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_431 bl[431] br[431] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_432 bl[432] br[432] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_433 bl[433] br[433] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_434 bl[434] br[434] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_435 bl[435] br[435] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_436 bl[436] br[436] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_437 bl[437] br[437] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_438 bl[438] br[438] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_439 bl[439] br[439] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_440 bl[440] br[440] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_441 bl[441] br[441] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_442 bl[442] br[442] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_443 bl[443] br[443] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_444 bl[444] br[444] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_445 bl[445] br[445] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_446 bl[446] br[446] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_447 bl[447] br[447] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_448 bl[448] br[448] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_449 bl[449] br[449] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_450 bl[450] br[450] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_451 bl[451] br[451] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_452 bl[452] br[452] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_453 bl[453] br[453] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_454 bl[454] br[454] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_455 bl[455] br[455] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_456 bl[456] br[456] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_457 bl[457] br[457] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_458 bl[458] br[458] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_459 bl[459] br[459] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_460 bl[460] br[460] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_461 bl[461] br[461] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_462 bl[462] br[462] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_463 bl[463] br[463] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_464 bl[464] br[464] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_465 bl[465] br[465] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_466 bl[466] br[466] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_467 bl[467] br[467] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_468 bl[468] br[468] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_469 bl[469] br[469] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_470 bl[470] br[470] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_471 bl[471] br[471] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_472 bl[472] br[472] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_473 bl[473] br[473] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_474 bl[474] br[474] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_475 bl[475] br[475] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_476 bl[476] br[476] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_477 bl[477] br[477] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_478 bl[478] br[478] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_479 bl[479] br[479] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_480 bl[480] br[480] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_481 bl[481] br[481] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_482 bl[482] br[482] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_483 bl[483] br[483] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_484 bl[484] br[484] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_485 bl[485] br[485] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_486 bl[486] br[486] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_487 bl[487] br[487] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_488 bl[488] br[488] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_489 bl[489] br[489] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_490 bl[490] br[490] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_491 bl[491] br[491] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_492 bl[492] br[492] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_493 bl[493] br[493] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_494 bl[494] br[494] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_495 bl[495] br[495] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_496 bl[496] br[496] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_497 bl[497] br[497] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_498 bl[498] br[498] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_499 bl[499] br[499] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_500 bl[500] br[500] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_501 bl[501] br[501] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_502 bl[502] br[502] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_503 bl[503] br[503] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_504 bl[504] br[504] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_505 bl[505] br[505] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_506 bl[506] br[506] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_507 bl[507] br[507] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_508 bl[508] br[508] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_509 bl[509] br[509] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_510 bl[510] br[510] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_45_511 bl[511] br[511] vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xcell_46_0 bl[0] br[0] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_1 bl[1] br[1] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_2 bl[2] br[2] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_3 bl[3] br[3] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_4 bl[4] br[4] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_5 bl[5] br[5] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_6 bl[6] br[6] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_7 bl[7] br[7] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_8 bl[8] br[8] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_9 bl[9] br[9] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_10 bl[10] br[10] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_11 bl[11] br[11] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_12 bl[12] br[12] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_13 bl[13] br[13] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_14 bl[14] br[14] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_15 bl[15] br[15] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_16 bl[16] br[16] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_17 bl[17] br[17] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_18 bl[18] br[18] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_19 bl[19] br[19] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_20 bl[20] br[20] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_21 bl[21] br[21] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_22 bl[22] br[22] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_23 bl[23] br[23] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_24 bl[24] br[24] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_25 bl[25] br[25] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_26 bl[26] br[26] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_27 bl[27] br[27] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_28 bl[28] br[28] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_29 bl[29] br[29] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_30 bl[30] br[30] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_31 bl[31] br[31] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_32 bl[32] br[32] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_33 bl[33] br[33] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_34 bl[34] br[34] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_35 bl[35] br[35] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_36 bl[36] br[36] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_37 bl[37] br[37] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_38 bl[38] br[38] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_39 bl[39] br[39] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_40 bl[40] br[40] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_41 bl[41] br[41] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_42 bl[42] br[42] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_43 bl[43] br[43] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_44 bl[44] br[44] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_45 bl[45] br[45] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_46 bl[46] br[46] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_47 bl[47] br[47] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_48 bl[48] br[48] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_49 bl[49] br[49] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_50 bl[50] br[50] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_51 bl[51] br[51] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_52 bl[52] br[52] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_53 bl[53] br[53] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_54 bl[54] br[54] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_55 bl[55] br[55] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_56 bl[56] br[56] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_57 bl[57] br[57] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_58 bl[58] br[58] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_59 bl[59] br[59] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_60 bl[60] br[60] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_61 bl[61] br[61] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_62 bl[62] br[62] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_63 bl[63] br[63] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_64 bl[64] br[64] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_65 bl[65] br[65] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_66 bl[66] br[66] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_67 bl[67] br[67] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_68 bl[68] br[68] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_69 bl[69] br[69] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_70 bl[70] br[70] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_71 bl[71] br[71] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_72 bl[72] br[72] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_73 bl[73] br[73] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_74 bl[74] br[74] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_75 bl[75] br[75] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_76 bl[76] br[76] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_77 bl[77] br[77] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_78 bl[78] br[78] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_79 bl[79] br[79] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_80 bl[80] br[80] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_81 bl[81] br[81] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_82 bl[82] br[82] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_83 bl[83] br[83] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_84 bl[84] br[84] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_85 bl[85] br[85] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_86 bl[86] br[86] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_87 bl[87] br[87] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_88 bl[88] br[88] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_89 bl[89] br[89] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_90 bl[90] br[90] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_91 bl[91] br[91] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_92 bl[92] br[92] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_93 bl[93] br[93] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_94 bl[94] br[94] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_95 bl[95] br[95] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_96 bl[96] br[96] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_97 bl[97] br[97] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_98 bl[98] br[98] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_99 bl[99] br[99] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_100 bl[100] br[100] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_101 bl[101] br[101] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_102 bl[102] br[102] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_103 bl[103] br[103] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_104 bl[104] br[104] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_105 bl[105] br[105] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_106 bl[106] br[106] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_107 bl[107] br[107] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_108 bl[108] br[108] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_109 bl[109] br[109] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_110 bl[110] br[110] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_111 bl[111] br[111] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_112 bl[112] br[112] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_113 bl[113] br[113] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_114 bl[114] br[114] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_115 bl[115] br[115] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_116 bl[116] br[116] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_117 bl[117] br[117] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_118 bl[118] br[118] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_119 bl[119] br[119] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_120 bl[120] br[120] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_121 bl[121] br[121] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_122 bl[122] br[122] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_123 bl[123] br[123] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_124 bl[124] br[124] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_125 bl[125] br[125] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_126 bl[126] br[126] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_127 bl[127] br[127] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_128 bl[128] br[128] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_129 bl[129] br[129] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_130 bl[130] br[130] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_131 bl[131] br[131] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_132 bl[132] br[132] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_133 bl[133] br[133] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_134 bl[134] br[134] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_135 bl[135] br[135] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_136 bl[136] br[136] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_137 bl[137] br[137] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_138 bl[138] br[138] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_139 bl[139] br[139] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_140 bl[140] br[140] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_141 bl[141] br[141] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_142 bl[142] br[142] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_143 bl[143] br[143] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_144 bl[144] br[144] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_145 bl[145] br[145] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_146 bl[146] br[146] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_147 bl[147] br[147] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_148 bl[148] br[148] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_149 bl[149] br[149] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_150 bl[150] br[150] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_151 bl[151] br[151] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_152 bl[152] br[152] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_153 bl[153] br[153] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_154 bl[154] br[154] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_155 bl[155] br[155] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_156 bl[156] br[156] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_157 bl[157] br[157] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_158 bl[158] br[158] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_159 bl[159] br[159] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_160 bl[160] br[160] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_161 bl[161] br[161] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_162 bl[162] br[162] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_163 bl[163] br[163] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_164 bl[164] br[164] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_165 bl[165] br[165] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_166 bl[166] br[166] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_167 bl[167] br[167] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_168 bl[168] br[168] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_169 bl[169] br[169] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_170 bl[170] br[170] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_171 bl[171] br[171] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_172 bl[172] br[172] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_173 bl[173] br[173] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_174 bl[174] br[174] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_175 bl[175] br[175] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_176 bl[176] br[176] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_177 bl[177] br[177] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_178 bl[178] br[178] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_179 bl[179] br[179] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_180 bl[180] br[180] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_181 bl[181] br[181] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_182 bl[182] br[182] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_183 bl[183] br[183] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_184 bl[184] br[184] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_185 bl[185] br[185] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_186 bl[186] br[186] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_187 bl[187] br[187] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_188 bl[188] br[188] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_189 bl[189] br[189] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_190 bl[190] br[190] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_191 bl[191] br[191] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_192 bl[192] br[192] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_193 bl[193] br[193] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_194 bl[194] br[194] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_195 bl[195] br[195] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_196 bl[196] br[196] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_197 bl[197] br[197] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_198 bl[198] br[198] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_199 bl[199] br[199] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_200 bl[200] br[200] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_201 bl[201] br[201] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_202 bl[202] br[202] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_203 bl[203] br[203] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_204 bl[204] br[204] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_205 bl[205] br[205] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_206 bl[206] br[206] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_207 bl[207] br[207] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_208 bl[208] br[208] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_209 bl[209] br[209] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_210 bl[210] br[210] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_211 bl[211] br[211] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_212 bl[212] br[212] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_213 bl[213] br[213] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_214 bl[214] br[214] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_215 bl[215] br[215] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_216 bl[216] br[216] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_217 bl[217] br[217] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_218 bl[218] br[218] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_219 bl[219] br[219] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_220 bl[220] br[220] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_221 bl[221] br[221] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_222 bl[222] br[222] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_223 bl[223] br[223] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_224 bl[224] br[224] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_225 bl[225] br[225] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_226 bl[226] br[226] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_227 bl[227] br[227] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_228 bl[228] br[228] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_229 bl[229] br[229] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_230 bl[230] br[230] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_231 bl[231] br[231] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_232 bl[232] br[232] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_233 bl[233] br[233] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_234 bl[234] br[234] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_235 bl[235] br[235] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_236 bl[236] br[236] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_237 bl[237] br[237] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_238 bl[238] br[238] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_239 bl[239] br[239] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_240 bl[240] br[240] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_241 bl[241] br[241] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_242 bl[242] br[242] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_243 bl[243] br[243] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_244 bl[244] br[244] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_245 bl[245] br[245] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_246 bl[246] br[246] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_247 bl[247] br[247] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_248 bl[248] br[248] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_249 bl[249] br[249] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_250 bl[250] br[250] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_251 bl[251] br[251] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_252 bl[252] br[252] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_253 bl[253] br[253] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_254 bl[254] br[254] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_255 bl[255] br[255] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_256 bl[256] br[256] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_257 bl[257] br[257] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_258 bl[258] br[258] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_259 bl[259] br[259] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_260 bl[260] br[260] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_261 bl[261] br[261] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_262 bl[262] br[262] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_263 bl[263] br[263] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_264 bl[264] br[264] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_265 bl[265] br[265] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_266 bl[266] br[266] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_267 bl[267] br[267] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_268 bl[268] br[268] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_269 bl[269] br[269] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_270 bl[270] br[270] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_271 bl[271] br[271] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_272 bl[272] br[272] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_273 bl[273] br[273] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_274 bl[274] br[274] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_275 bl[275] br[275] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_276 bl[276] br[276] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_277 bl[277] br[277] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_278 bl[278] br[278] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_279 bl[279] br[279] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_280 bl[280] br[280] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_281 bl[281] br[281] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_282 bl[282] br[282] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_283 bl[283] br[283] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_284 bl[284] br[284] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_285 bl[285] br[285] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_286 bl[286] br[286] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_287 bl[287] br[287] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_288 bl[288] br[288] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_289 bl[289] br[289] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_290 bl[290] br[290] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_291 bl[291] br[291] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_292 bl[292] br[292] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_293 bl[293] br[293] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_294 bl[294] br[294] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_295 bl[295] br[295] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_296 bl[296] br[296] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_297 bl[297] br[297] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_298 bl[298] br[298] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_299 bl[299] br[299] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_300 bl[300] br[300] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_301 bl[301] br[301] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_302 bl[302] br[302] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_303 bl[303] br[303] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_304 bl[304] br[304] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_305 bl[305] br[305] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_306 bl[306] br[306] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_307 bl[307] br[307] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_308 bl[308] br[308] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_309 bl[309] br[309] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_310 bl[310] br[310] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_311 bl[311] br[311] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_312 bl[312] br[312] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_313 bl[313] br[313] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_314 bl[314] br[314] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_315 bl[315] br[315] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_316 bl[316] br[316] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_317 bl[317] br[317] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_318 bl[318] br[318] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_319 bl[319] br[319] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_320 bl[320] br[320] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_321 bl[321] br[321] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_322 bl[322] br[322] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_323 bl[323] br[323] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_324 bl[324] br[324] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_325 bl[325] br[325] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_326 bl[326] br[326] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_327 bl[327] br[327] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_328 bl[328] br[328] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_329 bl[329] br[329] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_330 bl[330] br[330] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_331 bl[331] br[331] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_332 bl[332] br[332] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_333 bl[333] br[333] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_334 bl[334] br[334] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_335 bl[335] br[335] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_336 bl[336] br[336] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_337 bl[337] br[337] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_338 bl[338] br[338] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_339 bl[339] br[339] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_340 bl[340] br[340] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_341 bl[341] br[341] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_342 bl[342] br[342] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_343 bl[343] br[343] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_344 bl[344] br[344] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_345 bl[345] br[345] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_346 bl[346] br[346] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_347 bl[347] br[347] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_348 bl[348] br[348] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_349 bl[349] br[349] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_350 bl[350] br[350] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_351 bl[351] br[351] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_352 bl[352] br[352] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_353 bl[353] br[353] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_354 bl[354] br[354] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_355 bl[355] br[355] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_356 bl[356] br[356] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_357 bl[357] br[357] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_358 bl[358] br[358] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_359 bl[359] br[359] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_360 bl[360] br[360] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_361 bl[361] br[361] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_362 bl[362] br[362] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_363 bl[363] br[363] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_364 bl[364] br[364] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_365 bl[365] br[365] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_366 bl[366] br[366] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_367 bl[367] br[367] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_368 bl[368] br[368] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_369 bl[369] br[369] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_370 bl[370] br[370] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_371 bl[371] br[371] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_372 bl[372] br[372] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_373 bl[373] br[373] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_374 bl[374] br[374] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_375 bl[375] br[375] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_376 bl[376] br[376] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_377 bl[377] br[377] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_378 bl[378] br[378] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_379 bl[379] br[379] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_380 bl[380] br[380] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_381 bl[381] br[381] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_382 bl[382] br[382] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_383 bl[383] br[383] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_384 bl[384] br[384] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_385 bl[385] br[385] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_386 bl[386] br[386] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_387 bl[387] br[387] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_388 bl[388] br[388] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_389 bl[389] br[389] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_390 bl[390] br[390] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_391 bl[391] br[391] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_392 bl[392] br[392] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_393 bl[393] br[393] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_394 bl[394] br[394] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_395 bl[395] br[395] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_396 bl[396] br[396] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_397 bl[397] br[397] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_398 bl[398] br[398] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_399 bl[399] br[399] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_400 bl[400] br[400] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_401 bl[401] br[401] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_402 bl[402] br[402] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_403 bl[403] br[403] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_404 bl[404] br[404] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_405 bl[405] br[405] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_406 bl[406] br[406] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_407 bl[407] br[407] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_408 bl[408] br[408] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_409 bl[409] br[409] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_410 bl[410] br[410] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_411 bl[411] br[411] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_412 bl[412] br[412] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_413 bl[413] br[413] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_414 bl[414] br[414] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_415 bl[415] br[415] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_416 bl[416] br[416] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_417 bl[417] br[417] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_418 bl[418] br[418] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_419 bl[419] br[419] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_420 bl[420] br[420] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_421 bl[421] br[421] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_422 bl[422] br[422] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_423 bl[423] br[423] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_424 bl[424] br[424] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_425 bl[425] br[425] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_426 bl[426] br[426] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_427 bl[427] br[427] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_428 bl[428] br[428] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_429 bl[429] br[429] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_430 bl[430] br[430] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_431 bl[431] br[431] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_432 bl[432] br[432] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_433 bl[433] br[433] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_434 bl[434] br[434] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_435 bl[435] br[435] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_436 bl[436] br[436] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_437 bl[437] br[437] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_438 bl[438] br[438] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_439 bl[439] br[439] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_440 bl[440] br[440] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_441 bl[441] br[441] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_442 bl[442] br[442] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_443 bl[443] br[443] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_444 bl[444] br[444] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_445 bl[445] br[445] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_446 bl[446] br[446] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_447 bl[447] br[447] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_448 bl[448] br[448] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_449 bl[449] br[449] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_450 bl[450] br[450] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_451 bl[451] br[451] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_452 bl[452] br[452] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_453 bl[453] br[453] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_454 bl[454] br[454] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_455 bl[455] br[455] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_456 bl[456] br[456] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_457 bl[457] br[457] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_458 bl[458] br[458] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_459 bl[459] br[459] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_460 bl[460] br[460] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_461 bl[461] br[461] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_462 bl[462] br[462] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_463 bl[463] br[463] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_464 bl[464] br[464] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_465 bl[465] br[465] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_466 bl[466] br[466] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_467 bl[467] br[467] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_468 bl[468] br[468] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_469 bl[469] br[469] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_470 bl[470] br[470] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_471 bl[471] br[471] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_472 bl[472] br[472] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_473 bl[473] br[473] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_474 bl[474] br[474] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_475 bl[475] br[475] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_476 bl[476] br[476] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_477 bl[477] br[477] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_478 bl[478] br[478] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_479 bl[479] br[479] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_480 bl[480] br[480] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_481 bl[481] br[481] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_482 bl[482] br[482] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_483 bl[483] br[483] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_484 bl[484] br[484] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_485 bl[485] br[485] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_486 bl[486] br[486] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_487 bl[487] br[487] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_488 bl[488] br[488] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_489 bl[489] br[489] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_490 bl[490] br[490] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_491 bl[491] br[491] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_492 bl[492] br[492] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_493 bl[493] br[493] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_494 bl[494] br[494] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_495 bl[495] br[495] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_496 bl[496] br[496] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_497 bl[497] br[497] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_498 bl[498] br[498] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_499 bl[499] br[499] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_500 bl[500] br[500] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_501 bl[501] br[501] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_502 bl[502] br[502] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_503 bl[503] br[503] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_504 bl[504] br[504] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_505 bl[505] br[505] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_506 bl[506] br[506] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_507 bl[507] br[507] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_508 bl[508] br[508] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_509 bl[509] br[509] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_510 bl[510] br[510] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_46_511 bl[511] br[511] vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xcell_47_0 bl[0] br[0] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_1 bl[1] br[1] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_2 bl[2] br[2] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_3 bl[3] br[3] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_4 bl[4] br[4] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_5 bl[5] br[5] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_6 bl[6] br[6] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_7 bl[7] br[7] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_8 bl[8] br[8] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_9 bl[9] br[9] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_10 bl[10] br[10] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_11 bl[11] br[11] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_12 bl[12] br[12] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_13 bl[13] br[13] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_14 bl[14] br[14] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_15 bl[15] br[15] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_16 bl[16] br[16] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_17 bl[17] br[17] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_18 bl[18] br[18] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_19 bl[19] br[19] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_20 bl[20] br[20] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_21 bl[21] br[21] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_22 bl[22] br[22] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_23 bl[23] br[23] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_24 bl[24] br[24] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_25 bl[25] br[25] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_26 bl[26] br[26] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_27 bl[27] br[27] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_28 bl[28] br[28] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_29 bl[29] br[29] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_30 bl[30] br[30] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_31 bl[31] br[31] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_32 bl[32] br[32] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_33 bl[33] br[33] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_34 bl[34] br[34] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_35 bl[35] br[35] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_36 bl[36] br[36] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_37 bl[37] br[37] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_38 bl[38] br[38] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_39 bl[39] br[39] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_40 bl[40] br[40] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_41 bl[41] br[41] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_42 bl[42] br[42] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_43 bl[43] br[43] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_44 bl[44] br[44] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_45 bl[45] br[45] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_46 bl[46] br[46] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_47 bl[47] br[47] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_48 bl[48] br[48] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_49 bl[49] br[49] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_50 bl[50] br[50] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_51 bl[51] br[51] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_52 bl[52] br[52] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_53 bl[53] br[53] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_54 bl[54] br[54] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_55 bl[55] br[55] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_56 bl[56] br[56] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_57 bl[57] br[57] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_58 bl[58] br[58] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_59 bl[59] br[59] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_60 bl[60] br[60] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_61 bl[61] br[61] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_62 bl[62] br[62] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_63 bl[63] br[63] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_64 bl[64] br[64] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_65 bl[65] br[65] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_66 bl[66] br[66] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_67 bl[67] br[67] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_68 bl[68] br[68] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_69 bl[69] br[69] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_70 bl[70] br[70] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_71 bl[71] br[71] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_72 bl[72] br[72] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_73 bl[73] br[73] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_74 bl[74] br[74] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_75 bl[75] br[75] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_76 bl[76] br[76] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_77 bl[77] br[77] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_78 bl[78] br[78] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_79 bl[79] br[79] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_80 bl[80] br[80] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_81 bl[81] br[81] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_82 bl[82] br[82] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_83 bl[83] br[83] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_84 bl[84] br[84] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_85 bl[85] br[85] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_86 bl[86] br[86] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_87 bl[87] br[87] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_88 bl[88] br[88] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_89 bl[89] br[89] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_90 bl[90] br[90] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_91 bl[91] br[91] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_92 bl[92] br[92] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_93 bl[93] br[93] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_94 bl[94] br[94] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_95 bl[95] br[95] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_96 bl[96] br[96] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_97 bl[97] br[97] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_98 bl[98] br[98] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_99 bl[99] br[99] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_100 bl[100] br[100] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_101 bl[101] br[101] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_102 bl[102] br[102] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_103 bl[103] br[103] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_104 bl[104] br[104] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_105 bl[105] br[105] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_106 bl[106] br[106] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_107 bl[107] br[107] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_108 bl[108] br[108] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_109 bl[109] br[109] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_110 bl[110] br[110] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_111 bl[111] br[111] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_112 bl[112] br[112] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_113 bl[113] br[113] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_114 bl[114] br[114] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_115 bl[115] br[115] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_116 bl[116] br[116] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_117 bl[117] br[117] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_118 bl[118] br[118] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_119 bl[119] br[119] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_120 bl[120] br[120] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_121 bl[121] br[121] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_122 bl[122] br[122] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_123 bl[123] br[123] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_124 bl[124] br[124] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_125 bl[125] br[125] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_126 bl[126] br[126] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_127 bl[127] br[127] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_128 bl[128] br[128] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_129 bl[129] br[129] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_130 bl[130] br[130] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_131 bl[131] br[131] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_132 bl[132] br[132] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_133 bl[133] br[133] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_134 bl[134] br[134] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_135 bl[135] br[135] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_136 bl[136] br[136] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_137 bl[137] br[137] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_138 bl[138] br[138] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_139 bl[139] br[139] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_140 bl[140] br[140] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_141 bl[141] br[141] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_142 bl[142] br[142] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_143 bl[143] br[143] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_144 bl[144] br[144] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_145 bl[145] br[145] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_146 bl[146] br[146] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_147 bl[147] br[147] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_148 bl[148] br[148] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_149 bl[149] br[149] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_150 bl[150] br[150] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_151 bl[151] br[151] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_152 bl[152] br[152] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_153 bl[153] br[153] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_154 bl[154] br[154] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_155 bl[155] br[155] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_156 bl[156] br[156] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_157 bl[157] br[157] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_158 bl[158] br[158] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_159 bl[159] br[159] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_160 bl[160] br[160] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_161 bl[161] br[161] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_162 bl[162] br[162] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_163 bl[163] br[163] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_164 bl[164] br[164] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_165 bl[165] br[165] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_166 bl[166] br[166] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_167 bl[167] br[167] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_168 bl[168] br[168] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_169 bl[169] br[169] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_170 bl[170] br[170] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_171 bl[171] br[171] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_172 bl[172] br[172] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_173 bl[173] br[173] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_174 bl[174] br[174] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_175 bl[175] br[175] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_176 bl[176] br[176] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_177 bl[177] br[177] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_178 bl[178] br[178] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_179 bl[179] br[179] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_180 bl[180] br[180] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_181 bl[181] br[181] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_182 bl[182] br[182] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_183 bl[183] br[183] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_184 bl[184] br[184] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_185 bl[185] br[185] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_186 bl[186] br[186] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_187 bl[187] br[187] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_188 bl[188] br[188] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_189 bl[189] br[189] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_190 bl[190] br[190] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_191 bl[191] br[191] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_192 bl[192] br[192] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_193 bl[193] br[193] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_194 bl[194] br[194] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_195 bl[195] br[195] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_196 bl[196] br[196] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_197 bl[197] br[197] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_198 bl[198] br[198] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_199 bl[199] br[199] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_200 bl[200] br[200] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_201 bl[201] br[201] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_202 bl[202] br[202] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_203 bl[203] br[203] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_204 bl[204] br[204] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_205 bl[205] br[205] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_206 bl[206] br[206] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_207 bl[207] br[207] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_208 bl[208] br[208] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_209 bl[209] br[209] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_210 bl[210] br[210] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_211 bl[211] br[211] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_212 bl[212] br[212] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_213 bl[213] br[213] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_214 bl[214] br[214] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_215 bl[215] br[215] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_216 bl[216] br[216] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_217 bl[217] br[217] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_218 bl[218] br[218] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_219 bl[219] br[219] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_220 bl[220] br[220] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_221 bl[221] br[221] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_222 bl[222] br[222] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_223 bl[223] br[223] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_224 bl[224] br[224] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_225 bl[225] br[225] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_226 bl[226] br[226] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_227 bl[227] br[227] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_228 bl[228] br[228] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_229 bl[229] br[229] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_230 bl[230] br[230] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_231 bl[231] br[231] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_232 bl[232] br[232] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_233 bl[233] br[233] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_234 bl[234] br[234] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_235 bl[235] br[235] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_236 bl[236] br[236] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_237 bl[237] br[237] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_238 bl[238] br[238] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_239 bl[239] br[239] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_240 bl[240] br[240] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_241 bl[241] br[241] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_242 bl[242] br[242] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_243 bl[243] br[243] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_244 bl[244] br[244] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_245 bl[245] br[245] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_246 bl[246] br[246] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_247 bl[247] br[247] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_248 bl[248] br[248] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_249 bl[249] br[249] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_250 bl[250] br[250] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_251 bl[251] br[251] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_252 bl[252] br[252] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_253 bl[253] br[253] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_254 bl[254] br[254] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_255 bl[255] br[255] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_256 bl[256] br[256] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_257 bl[257] br[257] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_258 bl[258] br[258] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_259 bl[259] br[259] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_260 bl[260] br[260] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_261 bl[261] br[261] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_262 bl[262] br[262] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_263 bl[263] br[263] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_264 bl[264] br[264] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_265 bl[265] br[265] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_266 bl[266] br[266] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_267 bl[267] br[267] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_268 bl[268] br[268] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_269 bl[269] br[269] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_270 bl[270] br[270] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_271 bl[271] br[271] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_272 bl[272] br[272] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_273 bl[273] br[273] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_274 bl[274] br[274] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_275 bl[275] br[275] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_276 bl[276] br[276] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_277 bl[277] br[277] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_278 bl[278] br[278] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_279 bl[279] br[279] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_280 bl[280] br[280] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_281 bl[281] br[281] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_282 bl[282] br[282] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_283 bl[283] br[283] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_284 bl[284] br[284] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_285 bl[285] br[285] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_286 bl[286] br[286] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_287 bl[287] br[287] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_288 bl[288] br[288] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_289 bl[289] br[289] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_290 bl[290] br[290] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_291 bl[291] br[291] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_292 bl[292] br[292] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_293 bl[293] br[293] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_294 bl[294] br[294] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_295 bl[295] br[295] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_296 bl[296] br[296] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_297 bl[297] br[297] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_298 bl[298] br[298] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_299 bl[299] br[299] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_300 bl[300] br[300] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_301 bl[301] br[301] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_302 bl[302] br[302] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_303 bl[303] br[303] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_304 bl[304] br[304] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_305 bl[305] br[305] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_306 bl[306] br[306] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_307 bl[307] br[307] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_308 bl[308] br[308] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_309 bl[309] br[309] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_310 bl[310] br[310] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_311 bl[311] br[311] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_312 bl[312] br[312] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_313 bl[313] br[313] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_314 bl[314] br[314] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_315 bl[315] br[315] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_316 bl[316] br[316] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_317 bl[317] br[317] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_318 bl[318] br[318] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_319 bl[319] br[319] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_320 bl[320] br[320] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_321 bl[321] br[321] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_322 bl[322] br[322] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_323 bl[323] br[323] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_324 bl[324] br[324] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_325 bl[325] br[325] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_326 bl[326] br[326] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_327 bl[327] br[327] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_328 bl[328] br[328] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_329 bl[329] br[329] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_330 bl[330] br[330] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_331 bl[331] br[331] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_332 bl[332] br[332] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_333 bl[333] br[333] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_334 bl[334] br[334] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_335 bl[335] br[335] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_336 bl[336] br[336] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_337 bl[337] br[337] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_338 bl[338] br[338] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_339 bl[339] br[339] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_340 bl[340] br[340] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_341 bl[341] br[341] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_342 bl[342] br[342] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_343 bl[343] br[343] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_344 bl[344] br[344] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_345 bl[345] br[345] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_346 bl[346] br[346] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_347 bl[347] br[347] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_348 bl[348] br[348] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_349 bl[349] br[349] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_350 bl[350] br[350] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_351 bl[351] br[351] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_352 bl[352] br[352] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_353 bl[353] br[353] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_354 bl[354] br[354] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_355 bl[355] br[355] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_356 bl[356] br[356] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_357 bl[357] br[357] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_358 bl[358] br[358] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_359 bl[359] br[359] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_360 bl[360] br[360] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_361 bl[361] br[361] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_362 bl[362] br[362] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_363 bl[363] br[363] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_364 bl[364] br[364] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_365 bl[365] br[365] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_366 bl[366] br[366] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_367 bl[367] br[367] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_368 bl[368] br[368] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_369 bl[369] br[369] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_370 bl[370] br[370] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_371 bl[371] br[371] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_372 bl[372] br[372] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_373 bl[373] br[373] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_374 bl[374] br[374] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_375 bl[375] br[375] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_376 bl[376] br[376] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_377 bl[377] br[377] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_378 bl[378] br[378] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_379 bl[379] br[379] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_380 bl[380] br[380] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_381 bl[381] br[381] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_382 bl[382] br[382] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_383 bl[383] br[383] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_384 bl[384] br[384] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_385 bl[385] br[385] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_386 bl[386] br[386] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_387 bl[387] br[387] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_388 bl[388] br[388] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_389 bl[389] br[389] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_390 bl[390] br[390] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_391 bl[391] br[391] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_392 bl[392] br[392] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_393 bl[393] br[393] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_394 bl[394] br[394] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_395 bl[395] br[395] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_396 bl[396] br[396] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_397 bl[397] br[397] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_398 bl[398] br[398] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_399 bl[399] br[399] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_400 bl[400] br[400] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_401 bl[401] br[401] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_402 bl[402] br[402] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_403 bl[403] br[403] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_404 bl[404] br[404] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_405 bl[405] br[405] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_406 bl[406] br[406] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_407 bl[407] br[407] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_408 bl[408] br[408] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_409 bl[409] br[409] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_410 bl[410] br[410] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_411 bl[411] br[411] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_412 bl[412] br[412] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_413 bl[413] br[413] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_414 bl[414] br[414] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_415 bl[415] br[415] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_416 bl[416] br[416] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_417 bl[417] br[417] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_418 bl[418] br[418] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_419 bl[419] br[419] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_420 bl[420] br[420] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_421 bl[421] br[421] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_422 bl[422] br[422] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_423 bl[423] br[423] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_424 bl[424] br[424] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_425 bl[425] br[425] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_426 bl[426] br[426] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_427 bl[427] br[427] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_428 bl[428] br[428] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_429 bl[429] br[429] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_430 bl[430] br[430] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_431 bl[431] br[431] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_432 bl[432] br[432] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_433 bl[433] br[433] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_434 bl[434] br[434] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_435 bl[435] br[435] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_436 bl[436] br[436] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_437 bl[437] br[437] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_438 bl[438] br[438] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_439 bl[439] br[439] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_440 bl[440] br[440] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_441 bl[441] br[441] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_442 bl[442] br[442] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_443 bl[443] br[443] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_444 bl[444] br[444] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_445 bl[445] br[445] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_446 bl[446] br[446] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_447 bl[447] br[447] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_448 bl[448] br[448] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_449 bl[449] br[449] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_450 bl[450] br[450] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_451 bl[451] br[451] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_452 bl[452] br[452] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_453 bl[453] br[453] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_454 bl[454] br[454] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_455 bl[455] br[455] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_456 bl[456] br[456] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_457 bl[457] br[457] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_458 bl[458] br[458] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_459 bl[459] br[459] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_460 bl[460] br[460] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_461 bl[461] br[461] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_462 bl[462] br[462] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_463 bl[463] br[463] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_464 bl[464] br[464] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_465 bl[465] br[465] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_466 bl[466] br[466] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_467 bl[467] br[467] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_468 bl[468] br[468] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_469 bl[469] br[469] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_470 bl[470] br[470] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_471 bl[471] br[471] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_472 bl[472] br[472] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_473 bl[473] br[473] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_474 bl[474] br[474] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_475 bl[475] br[475] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_476 bl[476] br[476] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_477 bl[477] br[477] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_478 bl[478] br[478] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_479 bl[479] br[479] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_480 bl[480] br[480] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_481 bl[481] br[481] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_482 bl[482] br[482] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_483 bl[483] br[483] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_484 bl[484] br[484] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_485 bl[485] br[485] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_486 bl[486] br[486] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_487 bl[487] br[487] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_488 bl[488] br[488] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_489 bl[489] br[489] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_490 bl[490] br[490] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_491 bl[491] br[491] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_492 bl[492] br[492] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_493 bl[493] br[493] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_494 bl[494] br[494] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_495 bl[495] br[495] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_496 bl[496] br[496] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_497 bl[497] br[497] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_498 bl[498] br[498] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_499 bl[499] br[499] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_500 bl[500] br[500] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_501 bl[501] br[501] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_502 bl[502] br[502] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_503 bl[503] br[503] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_504 bl[504] br[504] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_505 bl[505] br[505] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_506 bl[506] br[506] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_507 bl[507] br[507] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_508 bl[508] br[508] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_509 bl[509] br[509] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_510 bl[510] br[510] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_47_511 bl[511] br[511] vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xcell_48_0 bl[0] br[0] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_1 bl[1] br[1] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_2 bl[2] br[2] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_3 bl[3] br[3] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_4 bl[4] br[4] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_5 bl[5] br[5] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_6 bl[6] br[6] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_7 bl[7] br[7] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_8 bl[8] br[8] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_9 bl[9] br[9] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_10 bl[10] br[10] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_11 bl[11] br[11] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_12 bl[12] br[12] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_13 bl[13] br[13] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_14 bl[14] br[14] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_15 bl[15] br[15] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_16 bl[16] br[16] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_17 bl[17] br[17] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_18 bl[18] br[18] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_19 bl[19] br[19] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_20 bl[20] br[20] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_21 bl[21] br[21] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_22 bl[22] br[22] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_23 bl[23] br[23] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_24 bl[24] br[24] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_25 bl[25] br[25] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_26 bl[26] br[26] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_27 bl[27] br[27] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_28 bl[28] br[28] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_29 bl[29] br[29] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_30 bl[30] br[30] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_31 bl[31] br[31] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_32 bl[32] br[32] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_33 bl[33] br[33] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_34 bl[34] br[34] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_35 bl[35] br[35] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_36 bl[36] br[36] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_37 bl[37] br[37] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_38 bl[38] br[38] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_39 bl[39] br[39] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_40 bl[40] br[40] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_41 bl[41] br[41] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_42 bl[42] br[42] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_43 bl[43] br[43] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_44 bl[44] br[44] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_45 bl[45] br[45] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_46 bl[46] br[46] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_47 bl[47] br[47] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_48 bl[48] br[48] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_49 bl[49] br[49] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_50 bl[50] br[50] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_51 bl[51] br[51] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_52 bl[52] br[52] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_53 bl[53] br[53] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_54 bl[54] br[54] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_55 bl[55] br[55] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_56 bl[56] br[56] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_57 bl[57] br[57] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_58 bl[58] br[58] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_59 bl[59] br[59] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_60 bl[60] br[60] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_61 bl[61] br[61] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_62 bl[62] br[62] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_63 bl[63] br[63] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_64 bl[64] br[64] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_65 bl[65] br[65] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_66 bl[66] br[66] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_67 bl[67] br[67] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_68 bl[68] br[68] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_69 bl[69] br[69] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_70 bl[70] br[70] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_71 bl[71] br[71] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_72 bl[72] br[72] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_73 bl[73] br[73] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_74 bl[74] br[74] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_75 bl[75] br[75] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_76 bl[76] br[76] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_77 bl[77] br[77] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_78 bl[78] br[78] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_79 bl[79] br[79] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_80 bl[80] br[80] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_81 bl[81] br[81] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_82 bl[82] br[82] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_83 bl[83] br[83] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_84 bl[84] br[84] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_85 bl[85] br[85] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_86 bl[86] br[86] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_87 bl[87] br[87] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_88 bl[88] br[88] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_89 bl[89] br[89] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_90 bl[90] br[90] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_91 bl[91] br[91] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_92 bl[92] br[92] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_93 bl[93] br[93] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_94 bl[94] br[94] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_95 bl[95] br[95] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_96 bl[96] br[96] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_97 bl[97] br[97] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_98 bl[98] br[98] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_99 bl[99] br[99] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_100 bl[100] br[100] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_101 bl[101] br[101] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_102 bl[102] br[102] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_103 bl[103] br[103] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_104 bl[104] br[104] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_105 bl[105] br[105] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_106 bl[106] br[106] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_107 bl[107] br[107] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_108 bl[108] br[108] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_109 bl[109] br[109] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_110 bl[110] br[110] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_111 bl[111] br[111] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_112 bl[112] br[112] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_113 bl[113] br[113] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_114 bl[114] br[114] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_115 bl[115] br[115] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_116 bl[116] br[116] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_117 bl[117] br[117] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_118 bl[118] br[118] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_119 bl[119] br[119] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_120 bl[120] br[120] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_121 bl[121] br[121] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_122 bl[122] br[122] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_123 bl[123] br[123] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_124 bl[124] br[124] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_125 bl[125] br[125] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_126 bl[126] br[126] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_127 bl[127] br[127] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_128 bl[128] br[128] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_129 bl[129] br[129] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_130 bl[130] br[130] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_131 bl[131] br[131] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_132 bl[132] br[132] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_133 bl[133] br[133] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_134 bl[134] br[134] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_135 bl[135] br[135] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_136 bl[136] br[136] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_137 bl[137] br[137] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_138 bl[138] br[138] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_139 bl[139] br[139] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_140 bl[140] br[140] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_141 bl[141] br[141] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_142 bl[142] br[142] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_143 bl[143] br[143] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_144 bl[144] br[144] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_145 bl[145] br[145] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_146 bl[146] br[146] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_147 bl[147] br[147] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_148 bl[148] br[148] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_149 bl[149] br[149] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_150 bl[150] br[150] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_151 bl[151] br[151] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_152 bl[152] br[152] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_153 bl[153] br[153] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_154 bl[154] br[154] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_155 bl[155] br[155] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_156 bl[156] br[156] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_157 bl[157] br[157] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_158 bl[158] br[158] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_159 bl[159] br[159] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_160 bl[160] br[160] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_161 bl[161] br[161] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_162 bl[162] br[162] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_163 bl[163] br[163] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_164 bl[164] br[164] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_165 bl[165] br[165] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_166 bl[166] br[166] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_167 bl[167] br[167] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_168 bl[168] br[168] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_169 bl[169] br[169] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_170 bl[170] br[170] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_171 bl[171] br[171] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_172 bl[172] br[172] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_173 bl[173] br[173] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_174 bl[174] br[174] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_175 bl[175] br[175] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_176 bl[176] br[176] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_177 bl[177] br[177] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_178 bl[178] br[178] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_179 bl[179] br[179] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_180 bl[180] br[180] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_181 bl[181] br[181] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_182 bl[182] br[182] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_183 bl[183] br[183] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_184 bl[184] br[184] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_185 bl[185] br[185] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_186 bl[186] br[186] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_187 bl[187] br[187] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_188 bl[188] br[188] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_189 bl[189] br[189] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_190 bl[190] br[190] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_191 bl[191] br[191] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_192 bl[192] br[192] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_193 bl[193] br[193] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_194 bl[194] br[194] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_195 bl[195] br[195] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_196 bl[196] br[196] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_197 bl[197] br[197] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_198 bl[198] br[198] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_199 bl[199] br[199] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_200 bl[200] br[200] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_201 bl[201] br[201] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_202 bl[202] br[202] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_203 bl[203] br[203] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_204 bl[204] br[204] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_205 bl[205] br[205] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_206 bl[206] br[206] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_207 bl[207] br[207] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_208 bl[208] br[208] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_209 bl[209] br[209] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_210 bl[210] br[210] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_211 bl[211] br[211] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_212 bl[212] br[212] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_213 bl[213] br[213] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_214 bl[214] br[214] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_215 bl[215] br[215] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_216 bl[216] br[216] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_217 bl[217] br[217] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_218 bl[218] br[218] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_219 bl[219] br[219] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_220 bl[220] br[220] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_221 bl[221] br[221] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_222 bl[222] br[222] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_223 bl[223] br[223] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_224 bl[224] br[224] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_225 bl[225] br[225] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_226 bl[226] br[226] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_227 bl[227] br[227] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_228 bl[228] br[228] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_229 bl[229] br[229] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_230 bl[230] br[230] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_231 bl[231] br[231] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_232 bl[232] br[232] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_233 bl[233] br[233] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_234 bl[234] br[234] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_235 bl[235] br[235] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_236 bl[236] br[236] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_237 bl[237] br[237] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_238 bl[238] br[238] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_239 bl[239] br[239] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_240 bl[240] br[240] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_241 bl[241] br[241] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_242 bl[242] br[242] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_243 bl[243] br[243] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_244 bl[244] br[244] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_245 bl[245] br[245] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_246 bl[246] br[246] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_247 bl[247] br[247] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_248 bl[248] br[248] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_249 bl[249] br[249] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_250 bl[250] br[250] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_251 bl[251] br[251] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_252 bl[252] br[252] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_253 bl[253] br[253] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_254 bl[254] br[254] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_255 bl[255] br[255] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_256 bl[256] br[256] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_257 bl[257] br[257] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_258 bl[258] br[258] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_259 bl[259] br[259] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_260 bl[260] br[260] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_261 bl[261] br[261] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_262 bl[262] br[262] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_263 bl[263] br[263] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_264 bl[264] br[264] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_265 bl[265] br[265] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_266 bl[266] br[266] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_267 bl[267] br[267] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_268 bl[268] br[268] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_269 bl[269] br[269] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_270 bl[270] br[270] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_271 bl[271] br[271] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_272 bl[272] br[272] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_273 bl[273] br[273] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_274 bl[274] br[274] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_275 bl[275] br[275] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_276 bl[276] br[276] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_277 bl[277] br[277] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_278 bl[278] br[278] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_279 bl[279] br[279] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_280 bl[280] br[280] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_281 bl[281] br[281] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_282 bl[282] br[282] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_283 bl[283] br[283] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_284 bl[284] br[284] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_285 bl[285] br[285] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_286 bl[286] br[286] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_287 bl[287] br[287] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_288 bl[288] br[288] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_289 bl[289] br[289] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_290 bl[290] br[290] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_291 bl[291] br[291] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_292 bl[292] br[292] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_293 bl[293] br[293] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_294 bl[294] br[294] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_295 bl[295] br[295] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_296 bl[296] br[296] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_297 bl[297] br[297] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_298 bl[298] br[298] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_299 bl[299] br[299] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_300 bl[300] br[300] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_301 bl[301] br[301] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_302 bl[302] br[302] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_303 bl[303] br[303] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_304 bl[304] br[304] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_305 bl[305] br[305] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_306 bl[306] br[306] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_307 bl[307] br[307] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_308 bl[308] br[308] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_309 bl[309] br[309] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_310 bl[310] br[310] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_311 bl[311] br[311] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_312 bl[312] br[312] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_313 bl[313] br[313] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_314 bl[314] br[314] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_315 bl[315] br[315] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_316 bl[316] br[316] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_317 bl[317] br[317] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_318 bl[318] br[318] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_319 bl[319] br[319] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_320 bl[320] br[320] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_321 bl[321] br[321] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_322 bl[322] br[322] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_323 bl[323] br[323] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_324 bl[324] br[324] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_325 bl[325] br[325] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_326 bl[326] br[326] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_327 bl[327] br[327] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_328 bl[328] br[328] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_329 bl[329] br[329] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_330 bl[330] br[330] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_331 bl[331] br[331] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_332 bl[332] br[332] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_333 bl[333] br[333] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_334 bl[334] br[334] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_335 bl[335] br[335] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_336 bl[336] br[336] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_337 bl[337] br[337] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_338 bl[338] br[338] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_339 bl[339] br[339] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_340 bl[340] br[340] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_341 bl[341] br[341] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_342 bl[342] br[342] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_343 bl[343] br[343] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_344 bl[344] br[344] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_345 bl[345] br[345] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_346 bl[346] br[346] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_347 bl[347] br[347] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_348 bl[348] br[348] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_349 bl[349] br[349] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_350 bl[350] br[350] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_351 bl[351] br[351] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_352 bl[352] br[352] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_353 bl[353] br[353] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_354 bl[354] br[354] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_355 bl[355] br[355] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_356 bl[356] br[356] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_357 bl[357] br[357] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_358 bl[358] br[358] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_359 bl[359] br[359] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_360 bl[360] br[360] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_361 bl[361] br[361] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_362 bl[362] br[362] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_363 bl[363] br[363] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_364 bl[364] br[364] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_365 bl[365] br[365] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_366 bl[366] br[366] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_367 bl[367] br[367] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_368 bl[368] br[368] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_369 bl[369] br[369] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_370 bl[370] br[370] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_371 bl[371] br[371] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_372 bl[372] br[372] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_373 bl[373] br[373] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_374 bl[374] br[374] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_375 bl[375] br[375] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_376 bl[376] br[376] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_377 bl[377] br[377] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_378 bl[378] br[378] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_379 bl[379] br[379] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_380 bl[380] br[380] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_381 bl[381] br[381] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_382 bl[382] br[382] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_383 bl[383] br[383] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_384 bl[384] br[384] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_385 bl[385] br[385] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_386 bl[386] br[386] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_387 bl[387] br[387] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_388 bl[388] br[388] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_389 bl[389] br[389] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_390 bl[390] br[390] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_391 bl[391] br[391] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_392 bl[392] br[392] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_393 bl[393] br[393] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_394 bl[394] br[394] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_395 bl[395] br[395] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_396 bl[396] br[396] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_397 bl[397] br[397] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_398 bl[398] br[398] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_399 bl[399] br[399] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_400 bl[400] br[400] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_401 bl[401] br[401] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_402 bl[402] br[402] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_403 bl[403] br[403] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_404 bl[404] br[404] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_405 bl[405] br[405] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_406 bl[406] br[406] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_407 bl[407] br[407] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_408 bl[408] br[408] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_409 bl[409] br[409] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_410 bl[410] br[410] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_411 bl[411] br[411] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_412 bl[412] br[412] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_413 bl[413] br[413] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_414 bl[414] br[414] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_415 bl[415] br[415] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_416 bl[416] br[416] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_417 bl[417] br[417] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_418 bl[418] br[418] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_419 bl[419] br[419] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_420 bl[420] br[420] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_421 bl[421] br[421] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_422 bl[422] br[422] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_423 bl[423] br[423] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_424 bl[424] br[424] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_425 bl[425] br[425] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_426 bl[426] br[426] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_427 bl[427] br[427] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_428 bl[428] br[428] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_429 bl[429] br[429] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_430 bl[430] br[430] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_431 bl[431] br[431] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_432 bl[432] br[432] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_433 bl[433] br[433] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_434 bl[434] br[434] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_435 bl[435] br[435] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_436 bl[436] br[436] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_437 bl[437] br[437] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_438 bl[438] br[438] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_439 bl[439] br[439] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_440 bl[440] br[440] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_441 bl[441] br[441] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_442 bl[442] br[442] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_443 bl[443] br[443] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_444 bl[444] br[444] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_445 bl[445] br[445] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_446 bl[446] br[446] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_447 bl[447] br[447] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_448 bl[448] br[448] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_449 bl[449] br[449] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_450 bl[450] br[450] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_451 bl[451] br[451] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_452 bl[452] br[452] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_453 bl[453] br[453] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_454 bl[454] br[454] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_455 bl[455] br[455] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_456 bl[456] br[456] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_457 bl[457] br[457] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_458 bl[458] br[458] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_459 bl[459] br[459] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_460 bl[460] br[460] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_461 bl[461] br[461] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_462 bl[462] br[462] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_463 bl[463] br[463] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_464 bl[464] br[464] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_465 bl[465] br[465] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_466 bl[466] br[466] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_467 bl[467] br[467] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_468 bl[468] br[468] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_469 bl[469] br[469] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_470 bl[470] br[470] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_471 bl[471] br[471] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_472 bl[472] br[472] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_473 bl[473] br[473] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_474 bl[474] br[474] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_475 bl[475] br[475] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_476 bl[476] br[476] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_477 bl[477] br[477] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_478 bl[478] br[478] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_479 bl[479] br[479] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_480 bl[480] br[480] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_481 bl[481] br[481] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_482 bl[482] br[482] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_483 bl[483] br[483] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_484 bl[484] br[484] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_485 bl[485] br[485] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_486 bl[486] br[486] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_487 bl[487] br[487] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_488 bl[488] br[488] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_489 bl[489] br[489] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_490 bl[490] br[490] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_491 bl[491] br[491] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_492 bl[492] br[492] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_493 bl[493] br[493] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_494 bl[494] br[494] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_495 bl[495] br[495] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_496 bl[496] br[496] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_497 bl[497] br[497] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_498 bl[498] br[498] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_499 bl[499] br[499] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_500 bl[500] br[500] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_501 bl[501] br[501] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_502 bl[502] br[502] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_503 bl[503] br[503] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_504 bl[504] br[504] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_505 bl[505] br[505] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_506 bl[506] br[506] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_507 bl[507] br[507] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_508 bl[508] br[508] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_509 bl[509] br[509] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_510 bl[510] br[510] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_48_511 bl[511] br[511] vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xcell_49_0 bl[0] br[0] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_1 bl[1] br[1] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_2 bl[2] br[2] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_3 bl[3] br[3] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_4 bl[4] br[4] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_5 bl[5] br[5] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_6 bl[6] br[6] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_7 bl[7] br[7] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_8 bl[8] br[8] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_9 bl[9] br[9] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_10 bl[10] br[10] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_11 bl[11] br[11] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_12 bl[12] br[12] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_13 bl[13] br[13] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_14 bl[14] br[14] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_15 bl[15] br[15] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_16 bl[16] br[16] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_17 bl[17] br[17] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_18 bl[18] br[18] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_19 bl[19] br[19] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_20 bl[20] br[20] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_21 bl[21] br[21] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_22 bl[22] br[22] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_23 bl[23] br[23] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_24 bl[24] br[24] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_25 bl[25] br[25] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_26 bl[26] br[26] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_27 bl[27] br[27] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_28 bl[28] br[28] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_29 bl[29] br[29] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_30 bl[30] br[30] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_31 bl[31] br[31] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_32 bl[32] br[32] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_33 bl[33] br[33] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_34 bl[34] br[34] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_35 bl[35] br[35] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_36 bl[36] br[36] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_37 bl[37] br[37] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_38 bl[38] br[38] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_39 bl[39] br[39] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_40 bl[40] br[40] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_41 bl[41] br[41] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_42 bl[42] br[42] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_43 bl[43] br[43] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_44 bl[44] br[44] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_45 bl[45] br[45] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_46 bl[46] br[46] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_47 bl[47] br[47] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_48 bl[48] br[48] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_49 bl[49] br[49] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_50 bl[50] br[50] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_51 bl[51] br[51] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_52 bl[52] br[52] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_53 bl[53] br[53] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_54 bl[54] br[54] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_55 bl[55] br[55] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_56 bl[56] br[56] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_57 bl[57] br[57] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_58 bl[58] br[58] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_59 bl[59] br[59] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_60 bl[60] br[60] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_61 bl[61] br[61] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_62 bl[62] br[62] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_63 bl[63] br[63] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_64 bl[64] br[64] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_65 bl[65] br[65] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_66 bl[66] br[66] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_67 bl[67] br[67] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_68 bl[68] br[68] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_69 bl[69] br[69] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_70 bl[70] br[70] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_71 bl[71] br[71] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_72 bl[72] br[72] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_73 bl[73] br[73] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_74 bl[74] br[74] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_75 bl[75] br[75] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_76 bl[76] br[76] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_77 bl[77] br[77] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_78 bl[78] br[78] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_79 bl[79] br[79] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_80 bl[80] br[80] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_81 bl[81] br[81] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_82 bl[82] br[82] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_83 bl[83] br[83] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_84 bl[84] br[84] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_85 bl[85] br[85] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_86 bl[86] br[86] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_87 bl[87] br[87] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_88 bl[88] br[88] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_89 bl[89] br[89] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_90 bl[90] br[90] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_91 bl[91] br[91] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_92 bl[92] br[92] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_93 bl[93] br[93] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_94 bl[94] br[94] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_95 bl[95] br[95] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_96 bl[96] br[96] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_97 bl[97] br[97] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_98 bl[98] br[98] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_99 bl[99] br[99] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_100 bl[100] br[100] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_101 bl[101] br[101] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_102 bl[102] br[102] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_103 bl[103] br[103] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_104 bl[104] br[104] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_105 bl[105] br[105] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_106 bl[106] br[106] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_107 bl[107] br[107] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_108 bl[108] br[108] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_109 bl[109] br[109] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_110 bl[110] br[110] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_111 bl[111] br[111] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_112 bl[112] br[112] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_113 bl[113] br[113] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_114 bl[114] br[114] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_115 bl[115] br[115] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_116 bl[116] br[116] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_117 bl[117] br[117] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_118 bl[118] br[118] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_119 bl[119] br[119] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_120 bl[120] br[120] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_121 bl[121] br[121] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_122 bl[122] br[122] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_123 bl[123] br[123] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_124 bl[124] br[124] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_125 bl[125] br[125] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_126 bl[126] br[126] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_127 bl[127] br[127] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_128 bl[128] br[128] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_129 bl[129] br[129] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_130 bl[130] br[130] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_131 bl[131] br[131] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_132 bl[132] br[132] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_133 bl[133] br[133] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_134 bl[134] br[134] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_135 bl[135] br[135] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_136 bl[136] br[136] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_137 bl[137] br[137] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_138 bl[138] br[138] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_139 bl[139] br[139] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_140 bl[140] br[140] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_141 bl[141] br[141] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_142 bl[142] br[142] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_143 bl[143] br[143] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_144 bl[144] br[144] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_145 bl[145] br[145] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_146 bl[146] br[146] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_147 bl[147] br[147] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_148 bl[148] br[148] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_149 bl[149] br[149] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_150 bl[150] br[150] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_151 bl[151] br[151] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_152 bl[152] br[152] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_153 bl[153] br[153] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_154 bl[154] br[154] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_155 bl[155] br[155] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_156 bl[156] br[156] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_157 bl[157] br[157] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_158 bl[158] br[158] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_159 bl[159] br[159] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_160 bl[160] br[160] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_161 bl[161] br[161] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_162 bl[162] br[162] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_163 bl[163] br[163] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_164 bl[164] br[164] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_165 bl[165] br[165] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_166 bl[166] br[166] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_167 bl[167] br[167] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_168 bl[168] br[168] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_169 bl[169] br[169] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_170 bl[170] br[170] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_171 bl[171] br[171] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_172 bl[172] br[172] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_173 bl[173] br[173] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_174 bl[174] br[174] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_175 bl[175] br[175] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_176 bl[176] br[176] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_177 bl[177] br[177] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_178 bl[178] br[178] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_179 bl[179] br[179] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_180 bl[180] br[180] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_181 bl[181] br[181] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_182 bl[182] br[182] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_183 bl[183] br[183] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_184 bl[184] br[184] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_185 bl[185] br[185] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_186 bl[186] br[186] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_187 bl[187] br[187] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_188 bl[188] br[188] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_189 bl[189] br[189] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_190 bl[190] br[190] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_191 bl[191] br[191] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_192 bl[192] br[192] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_193 bl[193] br[193] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_194 bl[194] br[194] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_195 bl[195] br[195] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_196 bl[196] br[196] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_197 bl[197] br[197] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_198 bl[198] br[198] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_199 bl[199] br[199] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_200 bl[200] br[200] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_201 bl[201] br[201] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_202 bl[202] br[202] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_203 bl[203] br[203] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_204 bl[204] br[204] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_205 bl[205] br[205] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_206 bl[206] br[206] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_207 bl[207] br[207] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_208 bl[208] br[208] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_209 bl[209] br[209] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_210 bl[210] br[210] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_211 bl[211] br[211] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_212 bl[212] br[212] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_213 bl[213] br[213] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_214 bl[214] br[214] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_215 bl[215] br[215] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_216 bl[216] br[216] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_217 bl[217] br[217] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_218 bl[218] br[218] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_219 bl[219] br[219] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_220 bl[220] br[220] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_221 bl[221] br[221] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_222 bl[222] br[222] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_223 bl[223] br[223] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_224 bl[224] br[224] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_225 bl[225] br[225] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_226 bl[226] br[226] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_227 bl[227] br[227] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_228 bl[228] br[228] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_229 bl[229] br[229] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_230 bl[230] br[230] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_231 bl[231] br[231] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_232 bl[232] br[232] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_233 bl[233] br[233] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_234 bl[234] br[234] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_235 bl[235] br[235] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_236 bl[236] br[236] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_237 bl[237] br[237] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_238 bl[238] br[238] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_239 bl[239] br[239] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_240 bl[240] br[240] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_241 bl[241] br[241] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_242 bl[242] br[242] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_243 bl[243] br[243] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_244 bl[244] br[244] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_245 bl[245] br[245] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_246 bl[246] br[246] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_247 bl[247] br[247] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_248 bl[248] br[248] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_249 bl[249] br[249] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_250 bl[250] br[250] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_251 bl[251] br[251] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_252 bl[252] br[252] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_253 bl[253] br[253] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_254 bl[254] br[254] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_255 bl[255] br[255] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_256 bl[256] br[256] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_257 bl[257] br[257] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_258 bl[258] br[258] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_259 bl[259] br[259] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_260 bl[260] br[260] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_261 bl[261] br[261] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_262 bl[262] br[262] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_263 bl[263] br[263] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_264 bl[264] br[264] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_265 bl[265] br[265] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_266 bl[266] br[266] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_267 bl[267] br[267] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_268 bl[268] br[268] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_269 bl[269] br[269] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_270 bl[270] br[270] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_271 bl[271] br[271] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_272 bl[272] br[272] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_273 bl[273] br[273] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_274 bl[274] br[274] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_275 bl[275] br[275] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_276 bl[276] br[276] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_277 bl[277] br[277] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_278 bl[278] br[278] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_279 bl[279] br[279] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_280 bl[280] br[280] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_281 bl[281] br[281] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_282 bl[282] br[282] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_283 bl[283] br[283] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_284 bl[284] br[284] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_285 bl[285] br[285] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_286 bl[286] br[286] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_287 bl[287] br[287] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_288 bl[288] br[288] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_289 bl[289] br[289] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_290 bl[290] br[290] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_291 bl[291] br[291] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_292 bl[292] br[292] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_293 bl[293] br[293] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_294 bl[294] br[294] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_295 bl[295] br[295] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_296 bl[296] br[296] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_297 bl[297] br[297] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_298 bl[298] br[298] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_299 bl[299] br[299] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_300 bl[300] br[300] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_301 bl[301] br[301] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_302 bl[302] br[302] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_303 bl[303] br[303] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_304 bl[304] br[304] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_305 bl[305] br[305] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_306 bl[306] br[306] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_307 bl[307] br[307] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_308 bl[308] br[308] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_309 bl[309] br[309] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_310 bl[310] br[310] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_311 bl[311] br[311] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_312 bl[312] br[312] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_313 bl[313] br[313] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_314 bl[314] br[314] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_315 bl[315] br[315] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_316 bl[316] br[316] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_317 bl[317] br[317] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_318 bl[318] br[318] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_319 bl[319] br[319] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_320 bl[320] br[320] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_321 bl[321] br[321] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_322 bl[322] br[322] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_323 bl[323] br[323] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_324 bl[324] br[324] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_325 bl[325] br[325] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_326 bl[326] br[326] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_327 bl[327] br[327] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_328 bl[328] br[328] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_329 bl[329] br[329] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_330 bl[330] br[330] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_331 bl[331] br[331] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_332 bl[332] br[332] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_333 bl[333] br[333] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_334 bl[334] br[334] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_335 bl[335] br[335] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_336 bl[336] br[336] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_337 bl[337] br[337] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_338 bl[338] br[338] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_339 bl[339] br[339] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_340 bl[340] br[340] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_341 bl[341] br[341] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_342 bl[342] br[342] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_343 bl[343] br[343] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_344 bl[344] br[344] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_345 bl[345] br[345] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_346 bl[346] br[346] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_347 bl[347] br[347] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_348 bl[348] br[348] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_349 bl[349] br[349] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_350 bl[350] br[350] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_351 bl[351] br[351] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_352 bl[352] br[352] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_353 bl[353] br[353] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_354 bl[354] br[354] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_355 bl[355] br[355] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_356 bl[356] br[356] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_357 bl[357] br[357] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_358 bl[358] br[358] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_359 bl[359] br[359] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_360 bl[360] br[360] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_361 bl[361] br[361] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_362 bl[362] br[362] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_363 bl[363] br[363] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_364 bl[364] br[364] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_365 bl[365] br[365] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_366 bl[366] br[366] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_367 bl[367] br[367] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_368 bl[368] br[368] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_369 bl[369] br[369] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_370 bl[370] br[370] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_371 bl[371] br[371] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_372 bl[372] br[372] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_373 bl[373] br[373] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_374 bl[374] br[374] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_375 bl[375] br[375] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_376 bl[376] br[376] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_377 bl[377] br[377] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_378 bl[378] br[378] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_379 bl[379] br[379] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_380 bl[380] br[380] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_381 bl[381] br[381] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_382 bl[382] br[382] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_383 bl[383] br[383] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_384 bl[384] br[384] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_385 bl[385] br[385] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_386 bl[386] br[386] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_387 bl[387] br[387] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_388 bl[388] br[388] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_389 bl[389] br[389] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_390 bl[390] br[390] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_391 bl[391] br[391] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_392 bl[392] br[392] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_393 bl[393] br[393] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_394 bl[394] br[394] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_395 bl[395] br[395] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_396 bl[396] br[396] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_397 bl[397] br[397] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_398 bl[398] br[398] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_399 bl[399] br[399] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_400 bl[400] br[400] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_401 bl[401] br[401] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_402 bl[402] br[402] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_403 bl[403] br[403] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_404 bl[404] br[404] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_405 bl[405] br[405] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_406 bl[406] br[406] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_407 bl[407] br[407] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_408 bl[408] br[408] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_409 bl[409] br[409] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_410 bl[410] br[410] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_411 bl[411] br[411] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_412 bl[412] br[412] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_413 bl[413] br[413] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_414 bl[414] br[414] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_415 bl[415] br[415] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_416 bl[416] br[416] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_417 bl[417] br[417] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_418 bl[418] br[418] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_419 bl[419] br[419] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_420 bl[420] br[420] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_421 bl[421] br[421] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_422 bl[422] br[422] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_423 bl[423] br[423] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_424 bl[424] br[424] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_425 bl[425] br[425] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_426 bl[426] br[426] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_427 bl[427] br[427] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_428 bl[428] br[428] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_429 bl[429] br[429] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_430 bl[430] br[430] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_431 bl[431] br[431] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_432 bl[432] br[432] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_433 bl[433] br[433] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_434 bl[434] br[434] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_435 bl[435] br[435] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_436 bl[436] br[436] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_437 bl[437] br[437] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_438 bl[438] br[438] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_439 bl[439] br[439] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_440 bl[440] br[440] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_441 bl[441] br[441] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_442 bl[442] br[442] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_443 bl[443] br[443] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_444 bl[444] br[444] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_445 bl[445] br[445] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_446 bl[446] br[446] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_447 bl[447] br[447] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_448 bl[448] br[448] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_449 bl[449] br[449] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_450 bl[450] br[450] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_451 bl[451] br[451] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_452 bl[452] br[452] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_453 bl[453] br[453] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_454 bl[454] br[454] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_455 bl[455] br[455] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_456 bl[456] br[456] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_457 bl[457] br[457] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_458 bl[458] br[458] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_459 bl[459] br[459] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_460 bl[460] br[460] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_461 bl[461] br[461] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_462 bl[462] br[462] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_463 bl[463] br[463] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_464 bl[464] br[464] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_465 bl[465] br[465] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_466 bl[466] br[466] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_467 bl[467] br[467] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_468 bl[468] br[468] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_469 bl[469] br[469] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_470 bl[470] br[470] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_471 bl[471] br[471] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_472 bl[472] br[472] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_473 bl[473] br[473] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_474 bl[474] br[474] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_475 bl[475] br[475] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_476 bl[476] br[476] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_477 bl[477] br[477] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_478 bl[478] br[478] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_479 bl[479] br[479] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_480 bl[480] br[480] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_481 bl[481] br[481] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_482 bl[482] br[482] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_483 bl[483] br[483] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_484 bl[484] br[484] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_485 bl[485] br[485] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_486 bl[486] br[486] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_487 bl[487] br[487] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_488 bl[488] br[488] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_489 bl[489] br[489] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_490 bl[490] br[490] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_491 bl[491] br[491] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_492 bl[492] br[492] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_493 bl[493] br[493] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_494 bl[494] br[494] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_495 bl[495] br[495] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_496 bl[496] br[496] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_497 bl[497] br[497] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_498 bl[498] br[498] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_499 bl[499] br[499] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_500 bl[500] br[500] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_501 bl[501] br[501] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_502 bl[502] br[502] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_503 bl[503] br[503] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_504 bl[504] br[504] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_505 bl[505] br[505] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_506 bl[506] br[506] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_507 bl[507] br[507] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_508 bl[508] br[508] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_509 bl[509] br[509] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_510 bl[510] br[510] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_49_511 bl[511] br[511] vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xcell_50_0 bl[0] br[0] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_1 bl[1] br[1] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_2 bl[2] br[2] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_3 bl[3] br[3] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_4 bl[4] br[4] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_5 bl[5] br[5] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_6 bl[6] br[6] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_7 bl[7] br[7] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_8 bl[8] br[8] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_9 bl[9] br[9] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_10 bl[10] br[10] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_11 bl[11] br[11] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_12 bl[12] br[12] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_13 bl[13] br[13] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_14 bl[14] br[14] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_15 bl[15] br[15] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_16 bl[16] br[16] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_17 bl[17] br[17] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_18 bl[18] br[18] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_19 bl[19] br[19] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_20 bl[20] br[20] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_21 bl[21] br[21] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_22 bl[22] br[22] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_23 bl[23] br[23] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_24 bl[24] br[24] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_25 bl[25] br[25] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_26 bl[26] br[26] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_27 bl[27] br[27] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_28 bl[28] br[28] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_29 bl[29] br[29] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_30 bl[30] br[30] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_31 bl[31] br[31] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_32 bl[32] br[32] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_33 bl[33] br[33] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_34 bl[34] br[34] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_35 bl[35] br[35] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_36 bl[36] br[36] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_37 bl[37] br[37] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_38 bl[38] br[38] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_39 bl[39] br[39] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_40 bl[40] br[40] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_41 bl[41] br[41] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_42 bl[42] br[42] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_43 bl[43] br[43] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_44 bl[44] br[44] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_45 bl[45] br[45] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_46 bl[46] br[46] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_47 bl[47] br[47] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_48 bl[48] br[48] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_49 bl[49] br[49] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_50 bl[50] br[50] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_51 bl[51] br[51] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_52 bl[52] br[52] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_53 bl[53] br[53] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_54 bl[54] br[54] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_55 bl[55] br[55] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_56 bl[56] br[56] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_57 bl[57] br[57] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_58 bl[58] br[58] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_59 bl[59] br[59] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_60 bl[60] br[60] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_61 bl[61] br[61] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_62 bl[62] br[62] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_63 bl[63] br[63] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_64 bl[64] br[64] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_65 bl[65] br[65] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_66 bl[66] br[66] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_67 bl[67] br[67] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_68 bl[68] br[68] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_69 bl[69] br[69] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_70 bl[70] br[70] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_71 bl[71] br[71] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_72 bl[72] br[72] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_73 bl[73] br[73] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_74 bl[74] br[74] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_75 bl[75] br[75] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_76 bl[76] br[76] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_77 bl[77] br[77] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_78 bl[78] br[78] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_79 bl[79] br[79] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_80 bl[80] br[80] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_81 bl[81] br[81] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_82 bl[82] br[82] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_83 bl[83] br[83] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_84 bl[84] br[84] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_85 bl[85] br[85] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_86 bl[86] br[86] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_87 bl[87] br[87] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_88 bl[88] br[88] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_89 bl[89] br[89] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_90 bl[90] br[90] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_91 bl[91] br[91] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_92 bl[92] br[92] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_93 bl[93] br[93] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_94 bl[94] br[94] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_95 bl[95] br[95] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_96 bl[96] br[96] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_97 bl[97] br[97] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_98 bl[98] br[98] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_99 bl[99] br[99] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_100 bl[100] br[100] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_101 bl[101] br[101] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_102 bl[102] br[102] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_103 bl[103] br[103] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_104 bl[104] br[104] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_105 bl[105] br[105] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_106 bl[106] br[106] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_107 bl[107] br[107] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_108 bl[108] br[108] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_109 bl[109] br[109] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_110 bl[110] br[110] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_111 bl[111] br[111] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_112 bl[112] br[112] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_113 bl[113] br[113] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_114 bl[114] br[114] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_115 bl[115] br[115] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_116 bl[116] br[116] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_117 bl[117] br[117] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_118 bl[118] br[118] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_119 bl[119] br[119] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_120 bl[120] br[120] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_121 bl[121] br[121] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_122 bl[122] br[122] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_123 bl[123] br[123] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_124 bl[124] br[124] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_125 bl[125] br[125] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_126 bl[126] br[126] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_127 bl[127] br[127] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_128 bl[128] br[128] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_129 bl[129] br[129] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_130 bl[130] br[130] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_131 bl[131] br[131] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_132 bl[132] br[132] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_133 bl[133] br[133] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_134 bl[134] br[134] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_135 bl[135] br[135] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_136 bl[136] br[136] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_137 bl[137] br[137] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_138 bl[138] br[138] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_139 bl[139] br[139] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_140 bl[140] br[140] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_141 bl[141] br[141] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_142 bl[142] br[142] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_143 bl[143] br[143] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_144 bl[144] br[144] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_145 bl[145] br[145] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_146 bl[146] br[146] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_147 bl[147] br[147] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_148 bl[148] br[148] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_149 bl[149] br[149] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_150 bl[150] br[150] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_151 bl[151] br[151] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_152 bl[152] br[152] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_153 bl[153] br[153] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_154 bl[154] br[154] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_155 bl[155] br[155] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_156 bl[156] br[156] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_157 bl[157] br[157] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_158 bl[158] br[158] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_159 bl[159] br[159] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_160 bl[160] br[160] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_161 bl[161] br[161] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_162 bl[162] br[162] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_163 bl[163] br[163] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_164 bl[164] br[164] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_165 bl[165] br[165] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_166 bl[166] br[166] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_167 bl[167] br[167] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_168 bl[168] br[168] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_169 bl[169] br[169] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_170 bl[170] br[170] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_171 bl[171] br[171] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_172 bl[172] br[172] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_173 bl[173] br[173] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_174 bl[174] br[174] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_175 bl[175] br[175] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_176 bl[176] br[176] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_177 bl[177] br[177] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_178 bl[178] br[178] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_179 bl[179] br[179] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_180 bl[180] br[180] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_181 bl[181] br[181] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_182 bl[182] br[182] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_183 bl[183] br[183] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_184 bl[184] br[184] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_185 bl[185] br[185] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_186 bl[186] br[186] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_187 bl[187] br[187] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_188 bl[188] br[188] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_189 bl[189] br[189] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_190 bl[190] br[190] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_191 bl[191] br[191] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_192 bl[192] br[192] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_193 bl[193] br[193] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_194 bl[194] br[194] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_195 bl[195] br[195] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_196 bl[196] br[196] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_197 bl[197] br[197] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_198 bl[198] br[198] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_199 bl[199] br[199] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_200 bl[200] br[200] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_201 bl[201] br[201] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_202 bl[202] br[202] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_203 bl[203] br[203] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_204 bl[204] br[204] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_205 bl[205] br[205] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_206 bl[206] br[206] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_207 bl[207] br[207] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_208 bl[208] br[208] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_209 bl[209] br[209] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_210 bl[210] br[210] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_211 bl[211] br[211] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_212 bl[212] br[212] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_213 bl[213] br[213] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_214 bl[214] br[214] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_215 bl[215] br[215] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_216 bl[216] br[216] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_217 bl[217] br[217] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_218 bl[218] br[218] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_219 bl[219] br[219] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_220 bl[220] br[220] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_221 bl[221] br[221] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_222 bl[222] br[222] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_223 bl[223] br[223] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_224 bl[224] br[224] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_225 bl[225] br[225] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_226 bl[226] br[226] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_227 bl[227] br[227] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_228 bl[228] br[228] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_229 bl[229] br[229] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_230 bl[230] br[230] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_231 bl[231] br[231] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_232 bl[232] br[232] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_233 bl[233] br[233] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_234 bl[234] br[234] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_235 bl[235] br[235] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_236 bl[236] br[236] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_237 bl[237] br[237] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_238 bl[238] br[238] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_239 bl[239] br[239] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_240 bl[240] br[240] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_241 bl[241] br[241] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_242 bl[242] br[242] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_243 bl[243] br[243] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_244 bl[244] br[244] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_245 bl[245] br[245] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_246 bl[246] br[246] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_247 bl[247] br[247] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_248 bl[248] br[248] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_249 bl[249] br[249] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_250 bl[250] br[250] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_251 bl[251] br[251] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_252 bl[252] br[252] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_253 bl[253] br[253] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_254 bl[254] br[254] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_255 bl[255] br[255] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_256 bl[256] br[256] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_257 bl[257] br[257] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_258 bl[258] br[258] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_259 bl[259] br[259] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_260 bl[260] br[260] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_261 bl[261] br[261] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_262 bl[262] br[262] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_263 bl[263] br[263] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_264 bl[264] br[264] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_265 bl[265] br[265] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_266 bl[266] br[266] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_267 bl[267] br[267] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_268 bl[268] br[268] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_269 bl[269] br[269] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_270 bl[270] br[270] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_271 bl[271] br[271] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_272 bl[272] br[272] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_273 bl[273] br[273] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_274 bl[274] br[274] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_275 bl[275] br[275] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_276 bl[276] br[276] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_277 bl[277] br[277] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_278 bl[278] br[278] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_279 bl[279] br[279] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_280 bl[280] br[280] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_281 bl[281] br[281] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_282 bl[282] br[282] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_283 bl[283] br[283] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_284 bl[284] br[284] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_285 bl[285] br[285] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_286 bl[286] br[286] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_287 bl[287] br[287] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_288 bl[288] br[288] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_289 bl[289] br[289] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_290 bl[290] br[290] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_291 bl[291] br[291] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_292 bl[292] br[292] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_293 bl[293] br[293] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_294 bl[294] br[294] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_295 bl[295] br[295] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_296 bl[296] br[296] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_297 bl[297] br[297] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_298 bl[298] br[298] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_299 bl[299] br[299] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_300 bl[300] br[300] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_301 bl[301] br[301] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_302 bl[302] br[302] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_303 bl[303] br[303] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_304 bl[304] br[304] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_305 bl[305] br[305] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_306 bl[306] br[306] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_307 bl[307] br[307] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_308 bl[308] br[308] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_309 bl[309] br[309] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_310 bl[310] br[310] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_311 bl[311] br[311] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_312 bl[312] br[312] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_313 bl[313] br[313] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_314 bl[314] br[314] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_315 bl[315] br[315] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_316 bl[316] br[316] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_317 bl[317] br[317] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_318 bl[318] br[318] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_319 bl[319] br[319] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_320 bl[320] br[320] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_321 bl[321] br[321] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_322 bl[322] br[322] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_323 bl[323] br[323] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_324 bl[324] br[324] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_325 bl[325] br[325] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_326 bl[326] br[326] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_327 bl[327] br[327] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_328 bl[328] br[328] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_329 bl[329] br[329] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_330 bl[330] br[330] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_331 bl[331] br[331] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_332 bl[332] br[332] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_333 bl[333] br[333] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_334 bl[334] br[334] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_335 bl[335] br[335] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_336 bl[336] br[336] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_337 bl[337] br[337] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_338 bl[338] br[338] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_339 bl[339] br[339] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_340 bl[340] br[340] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_341 bl[341] br[341] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_342 bl[342] br[342] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_343 bl[343] br[343] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_344 bl[344] br[344] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_345 bl[345] br[345] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_346 bl[346] br[346] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_347 bl[347] br[347] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_348 bl[348] br[348] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_349 bl[349] br[349] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_350 bl[350] br[350] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_351 bl[351] br[351] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_352 bl[352] br[352] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_353 bl[353] br[353] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_354 bl[354] br[354] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_355 bl[355] br[355] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_356 bl[356] br[356] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_357 bl[357] br[357] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_358 bl[358] br[358] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_359 bl[359] br[359] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_360 bl[360] br[360] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_361 bl[361] br[361] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_362 bl[362] br[362] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_363 bl[363] br[363] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_364 bl[364] br[364] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_365 bl[365] br[365] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_366 bl[366] br[366] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_367 bl[367] br[367] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_368 bl[368] br[368] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_369 bl[369] br[369] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_370 bl[370] br[370] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_371 bl[371] br[371] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_372 bl[372] br[372] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_373 bl[373] br[373] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_374 bl[374] br[374] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_375 bl[375] br[375] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_376 bl[376] br[376] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_377 bl[377] br[377] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_378 bl[378] br[378] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_379 bl[379] br[379] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_380 bl[380] br[380] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_381 bl[381] br[381] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_382 bl[382] br[382] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_383 bl[383] br[383] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_384 bl[384] br[384] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_385 bl[385] br[385] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_386 bl[386] br[386] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_387 bl[387] br[387] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_388 bl[388] br[388] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_389 bl[389] br[389] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_390 bl[390] br[390] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_391 bl[391] br[391] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_392 bl[392] br[392] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_393 bl[393] br[393] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_394 bl[394] br[394] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_395 bl[395] br[395] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_396 bl[396] br[396] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_397 bl[397] br[397] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_398 bl[398] br[398] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_399 bl[399] br[399] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_400 bl[400] br[400] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_401 bl[401] br[401] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_402 bl[402] br[402] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_403 bl[403] br[403] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_404 bl[404] br[404] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_405 bl[405] br[405] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_406 bl[406] br[406] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_407 bl[407] br[407] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_408 bl[408] br[408] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_409 bl[409] br[409] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_410 bl[410] br[410] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_411 bl[411] br[411] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_412 bl[412] br[412] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_413 bl[413] br[413] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_414 bl[414] br[414] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_415 bl[415] br[415] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_416 bl[416] br[416] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_417 bl[417] br[417] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_418 bl[418] br[418] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_419 bl[419] br[419] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_420 bl[420] br[420] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_421 bl[421] br[421] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_422 bl[422] br[422] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_423 bl[423] br[423] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_424 bl[424] br[424] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_425 bl[425] br[425] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_426 bl[426] br[426] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_427 bl[427] br[427] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_428 bl[428] br[428] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_429 bl[429] br[429] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_430 bl[430] br[430] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_431 bl[431] br[431] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_432 bl[432] br[432] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_433 bl[433] br[433] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_434 bl[434] br[434] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_435 bl[435] br[435] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_436 bl[436] br[436] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_437 bl[437] br[437] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_438 bl[438] br[438] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_439 bl[439] br[439] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_440 bl[440] br[440] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_441 bl[441] br[441] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_442 bl[442] br[442] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_443 bl[443] br[443] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_444 bl[444] br[444] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_445 bl[445] br[445] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_446 bl[446] br[446] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_447 bl[447] br[447] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_448 bl[448] br[448] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_449 bl[449] br[449] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_450 bl[450] br[450] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_451 bl[451] br[451] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_452 bl[452] br[452] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_453 bl[453] br[453] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_454 bl[454] br[454] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_455 bl[455] br[455] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_456 bl[456] br[456] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_457 bl[457] br[457] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_458 bl[458] br[458] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_459 bl[459] br[459] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_460 bl[460] br[460] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_461 bl[461] br[461] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_462 bl[462] br[462] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_463 bl[463] br[463] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_464 bl[464] br[464] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_465 bl[465] br[465] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_466 bl[466] br[466] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_467 bl[467] br[467] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_468 bl[468] br[468] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_469 bl[469] br[469] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_470 bl[470] br[470] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_471 bl[471] br[471] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_472 bl[472] br[472] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_473 bl[473] br[473] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_474 bl[474] br[474] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_475 bl[475] br[475] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_476 bl[476] br[476] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_477 bl[477] br[477] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_478 bl[478] br[478] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_479 bl[479] br[479] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_480 bl[480] br[480] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_481 bl[481] br[481] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_482 bl[482] br[482] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_483 bl[483] br[483] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_484 bl[484] br[484] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_485 bl[485] br[485] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_486 bl[486] br[486] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_487 bl[487] br[487] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_488 bl[488] br[488] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_489 bl[489] br[489] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_490 bl[490] br[490] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_491 bl[491] br[491] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_492 bl[492] br[492] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_493 bl[493] br[493] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_494 bl[494] br[494] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_495 bl[495] br[495] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_496 bl[496] br[496] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_497 bl[497] br[497] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_498 bl[498] br[498] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_499 bl[499] br[499] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_500 bl[500] br[500] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_501 bl[501] br[501] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_502 bl[502] br[502] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_503 bl[503] br[503] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_504 bl[504] br[504] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_505 bl[505] br[505] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_506 bl[506] br[506] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_507 bl[507] br[507] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_508 bl[508] br[508] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_509 bl[509] br[509] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_510 bl[510] br[510] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_50_511 bl[511] br[511] vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xcell_51_0 bl[0] br[0] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_1 bl[1] br[1] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_2 bl[2] br[2] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_3 bl[3] br[3] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_4 bl[4] br[4] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_5 bl[5] br[5] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_6 bl[6] br[6] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_7 bl[7] br[7] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_8 bl[8] br[8] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_9 bl[9] br[9] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_10 bl[10] br[10] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_11 bl[11] br[11] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_12 bl[12] br[12] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_13 bl[13] br[13] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_14 bl[14] br[14] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_15 bl[15] br[15] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_16 bl[16] br[16] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_17 bl[17] br[17] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_18 bl[18] br[18] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_19 bl[19] br[19] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_20 bl[20] br[20] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_21 bl[21] br[21] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_22 bl[22] br[22] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_23 bl[23] br[23] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_24 bl[24] br[24] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_25 bl[25] br[25] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_26 bl[26] br[26] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_27 bl[27] br[27] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_28 bl[28] br[28] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_29 bl[29] br[29] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_30 bl[30] br[30] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_31 bl[31] br[31] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_32 bl[32] br[32] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_33 bl[33] br[33] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_34 bl[34] br[34] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_35 bl[35] br[35] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_36 bl[36] br[36] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_37 bl[37] br[37] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_38 bl[38] br[38] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_39 bl[39] br[39] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_40 bl[40] br[40] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_41 bl[41] br[41] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_42 bl[42] br[42] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_43 bl[43] br[43] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_44 bl[44] br[44] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_45 bl[45] br[45] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_46 bl[46] br[46] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_47 bl[47] br[47] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_48 bl[48] br[48] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_49 bl[49] br[49] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_50 bl[50] br[50] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_51 bl[51] br[51] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_52 bl[52] br[52] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_53 bl[53] br[53] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_54 bl[54] br[54] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_55 bl[55] br[55] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_56 bl[56] br[56] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_57 bl[57] br[57] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_58 bl[58] br[58] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_59 bl[59] br[59] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_60 bl[60] br[60] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_61 bl[61] br[61] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_62 bl[62] br[62] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_63 bl[63] br[63] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_64 bl[64] br[64] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_65 bl[65] br[65] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_66 bl[66] br[66] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_67 bl[67] br[67] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_68 bl[68] br[68] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_69 bl[69] br[69] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_70 bl[70] br[70] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_71 bl[71] br[71] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_72 bl[72] br[72] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_73 bl[73] br[73] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_74 bl[74] br[74] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_75 bl[75] br[75] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_76 bl[76] br[76] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_77 bl[77] br[77] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_78 bl[78] br[78] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_79 bl[79] br[79] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_80 bl[80] br[80] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_81 bl[81] br[81] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_82 bl[82] br[82] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_83 bl[83] br[83] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_84 bl[84] br[84] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_85 bl[85] br[85] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_86 bl[86] br[86] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_87 bl[87] br[87] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_88 bl[88] br[88] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_89 bl[89] br[89] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_90 bl[90] br[90] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_91 bl[91] br[91] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_92 bl[92] br[92] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_93 bl[93] br[93] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_94 bl[94] br[94] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_95 bl[95] br[95] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_96 bl[96] br[96] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_97 bl[97] br[97] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_98 bl[98] br[98] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_99 bl[99] br[99] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_100 bl[100] br[100] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_101 bl[101] br[101] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_102 bl[102] br[102] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_103 bl[103] br[103] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_104 bl[104] br[104] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_105 bl[105] br[105] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_106 bl[106] br[106] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_107 bl[107] br[107] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_108 bl[108] br[108] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_109 bl[109] br[109] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_110 bl[110] br[110] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_111 bl[111] br[111] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_112 bl[112] br[112] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_113 bl[113] br[113] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_114 bl[114] br[114] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_115 bl[115] br[115] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_116 bl[116] br[116] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_117 bl[117] br[117] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_118 bl[118] br[118] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_119 bl[119] br[119] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_120 bl[120] br[120] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_121 bl[121] br[121] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_122 bl[122] br[122] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_123 bl[123] br[123] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_124 bl[124] br[124] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_125 bl[125] br[125] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_126 bl[126] br[126] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_127 bl[127] br[127] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_128 bl[128] br[128] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_129 bl[129] br[129] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_130 bl[130] br[130] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_131 bl[131] br[131] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_132 bl[132] br[132] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_133 bl[133] br[133] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_134 bl[134] br[134] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_135 bl[135] br[135] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_136 bl[136] br[136] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_137 bl[137] br[137] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_138 bl[138] br[138] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_139 bl[139] br[139] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_140 bl[140] br[140] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_141 bl[141] br[141] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_142 bl[142] br[142] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_143 bl[143] br[143] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_144 bl[144] br[144] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_145 bl[145] br[145] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_146 bl[146] br[146] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_147 bl[147] br[147] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_148 bl[148] br[148] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_149 bl[149] br[149] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_150 bl[150] br[150] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_151 bl[151] br[151] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_152 bl[152] br[152] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_153 bl[153] br[153] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_154 bl[154] br[154] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_155 bl[155] br[155] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_156 bl[156] br[156] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_157 bl[157] br[157] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_158 bl[158] br[158] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_159 bl[159] br[159] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_160 bl[160] br[160] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_161 bl[161] br[161] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_162 bl[162] br[162] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_163 bl[163] br[163] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_164 bl[164] br[164] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_165 bl[165] br[165] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_166 bl[166] br[166] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_167 bl[167] br[167] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_168 bl[168] br[168] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_169 bl[169] br[169] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_170 bl[170] br[170] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_171 bl[171] br[171] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_172 bl[172] br[172] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_173 bl[173] br[173] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_174 bl[174] br[174] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_175 bl[175] br[175] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_176 bl[176] br[176] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_177 bl[177] br[177] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_178 bl[178] br[178] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_179 bl[179] br[179] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_180 bl[180] br[180] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_181 bl[181] br[181] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_182 bl[182] br[182] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_183 bl[183] br[183] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_184 bl[184] br[184] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_185 bl[185] br[185] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_186 bl[186] br[186] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_187 bl[187] br[187] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_188 bl[188] br[188] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_189 bl[189] br[189] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_190 bl[190] br[190] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_191 bl[191] br[191] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_192 bl[192] br[192] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_193 bl[193] br[193] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_194 bl[194] br[194] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_195 bl[195] br[195] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_196 bl[196] br[196] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_197 bl[197] br[197] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_198 bl[198] br[198] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_199 bl[199] br[199] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_200 bl[200] br[200] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_201 bl[201] br[201] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_202 bl[202] br[202] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_203 bl[203] br[203] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_204 bl[204] br[204] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_205 bl[205] br[205] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_206 bl[206] br[206] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_207 bl[207] br[207] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_208 bl[208] br[208] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_209 bl[209] br[209] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_210 bl[210] br[210] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_211 bl[211] br[211] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_212 bl[212] br[212] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_213 bl[213] br[213] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_214 bl[214] br[214] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_215 bl[215] br[215] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_216 bl[216] br[216] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_217 bl[217] br[217] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_218 bl[218] br[218] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_219 bl[219] br[219] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_220 bl[220] br[220] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_221 bl[221] br[221] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_222 bl[222] br[222] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_223 bl[223] br[223] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_224 bl[224] br[224] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_225 bl[225] br[225] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_226 bl[226] br[226] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_227 bl[227] br[227] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_228 bl[228] br[228] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_229 bl[229] br[229] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_230 bl[230] br[230] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_231 bl[231] br[231] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_232 bl[232] br[232] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_233 bl[233] br[233] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_234 bl[234] br[234] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_235 bl[235] br[235] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_236 bl[236] br[236] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_237 bl[237] br[237] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_238 bl[238] br[238] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_239 bl[239] br[239] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_240 bl[240] br[240] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_241 bl[241] br[241] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_242 bl[242] br[242] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_243 bl[243] br[243] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_244 bl[244] br[244] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_245 bl[245] br[245] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_246 bl[246] br[246] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_247 bl[247] br[247] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_248 bl[248] br[248] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_249 bl[249] br[249] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_250 bl[250] br[250] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_251 bl[251] br[251] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_252 bl[252] br[252] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_253 bl[253] br[253] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_254 bl[254] br[254] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_255 bl[255] br[255] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_256 bl[256] br[256] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_257 bl[257] br[257] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_258 bl[258] br[258] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_259 bl[259] br[259] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_260 bl[260] br[260] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_261 bl[261] br[261] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_262 bl[262] br[262] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_263 bl[263] br[263] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_264 bl[264] br[264] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_265 bl[265] br[265] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_266 bl[266] br[266] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_267 bl[267] br[267] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_268 bl[268] br[268] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_269 bl[269] br[269] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_270 bl[270] br[270] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_271 bl[271] br[271] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_272 bl[272] br[272] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_273 bl[273] br[273] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_274 bl[274] br[274] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_275 bl[275] br[275] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_276 bl[276] br[276] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_277 bl[277] br[277] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_278 bl[278] br[278] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_279 bl[279] br[279] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_280 bl[280] br[280] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_281 bl[281] br[281] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_282 bl[282] br[282] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_283 bl[283] br[283] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_284 bl[284] br[284] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_285 bl[285] br[285] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_286 bl[286] br[286] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_287 bl[287] br[287] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_288 bl[288] br[288] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_289 bl[289] br[289] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_290 bl[290] br[290] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_291 bl[291] br[291] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_292 bl[292] br[292] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_293 bl[293] br[293] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_294 bl[294] br[294] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_295 bl[295] br[295] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_296 bl[296] br[296] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_297 bl[297] br[297] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_298 bl[298] br[298] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_299 bl[299] br[299] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_300 bl[300] br[300] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_301 bl[301] br[301] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_302 bl[302] br[302] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_303 bl[303] br[303] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_304 bl[304] br[304] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_305 bl[305] br[305] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_306 bl[306] br[306] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_307 bl[307] br[307] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_308 bl[308] br[308] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_309 bl[309] br[309] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_310 bl[310] br[310] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_311 bl[311] br[311] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_312 bl[312] br[312] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_313 bl[313] br[313] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_314 bl[314] br[314] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_315 bl[315] br[315] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_316 bl[316] br[316] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_317 bl[317] br[317] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_318 bl[318] br[318] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_319 bl[319] br[319] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_320 bl[320] br[320] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_321 bl[321] br[321] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_322 bl[322] br[322] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_323 bl[323] br[323] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_324 bl[324] br[324] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_325 bl[325] br[325] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_326 bl[326] br[326] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_327 bl[327] br[327] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_328 bl[328] br[328] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_329 bl[329] br[329] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_330 bl[330] br[330] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_331 bl[331] br[331] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_332 bl[332] br[332] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_333 bl[333] br[333] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_334 bl[334] br[334] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_335 bl[335] br[335] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_336 bl[336] br[336] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_337 bl[337] br[337] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_338 bl[338] br[338] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_339 bl[339] br[339] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_340 bl[340] br[340] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_341 bl[341] br[341] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_342 bl[342] br[342] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_343 bl[343] br[343] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_344 bl[344] br[344] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_345 bl[345] br[345] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_346 bl[346] br[346] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_347 bl[347] br[347] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_348 bl[348] br[348] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_349 bl[349] br[349] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_350 bl[350] br[350] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_351 bl[351] br[351] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_352 bl[352] br[352] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_353 bl[353] br[353] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_354 bl[354] br[354] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_355 bl[355] br[355] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_356 bl[356] br[356] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_357 bl[357] br[357] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_358 bl[358] br[358] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_359 bl[359] br[359] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_360 bl[360] br[360] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_361 bl[361] br[361] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_362 bl[362] br[362] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_363 bl[363] br[363] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_364 bl[364] br[364] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_365 bl[365] br[365] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_366 bl[366] br[366] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_367 bl[367] br[367] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_368 bl[368] br[368] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_369 bl[369] br[369] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_370 bl[370] br[370] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_371 bl[371] br[371] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_372 bl[372] br[372] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_373 bl[373] br[373] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_374 bl[374] br[374] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_375 bl[375] br[375] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_376 bl[376] br[376] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_377 bl[377] br[377] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_378 bl[378] br[378] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_379 bl[379] br[379] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_380 bl[380] br[380] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_381 bl[381] br[381] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_382 bl[382] br[382] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_383 bl[383] br[383] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_384 bl[384] br[384] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_385 bl[385] br[385] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_386 bl[386] br[386] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_387 bl[387] br[387] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_388 bl[388] br[388] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_389 bl[389] br[389] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_390 bl[390] br[390] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_391 bl[391] br[391] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_392 bl[392] br[392] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_393 bl[393] br[393] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_394 bl[394] br[394] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_395 bl[395] br[395] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_396 bl[396] br[396] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_397 bl[397] br[397] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_398 bl[398] br[398] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_399 bl[399] br[399] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_400 bl[400] br[400] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_401 bl[401] br[401] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_402 bl[402] br[402] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_403 bl[403] br[403] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_404 bl[404] br[404] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_405 bl[405] br[405] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_406 bl[406] br[406] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_407 bl[407] br[407] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_408 bl[408] br[408] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_409 bl[409] br[409] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_410 bl[410] br[410] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_411 bl[411] br[411] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_412 bl[412] br[412] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_413 bl[413] br[413] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_414 bl[414] br[414] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_415 bl[415] br[415] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_416 bl[416] br[416] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_417 bl[417] br[417] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_418 bl[418] br[418] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_419 bl[419] br[419] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_420 bl[420] br[420] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_421 bl[421] br[421] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_422 bl[422] br[422] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_423 bl[423] br[423] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_424 bl[424] br[424] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_425 bl[425] br[425] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_426 bl[426] br[426] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_427 bl[427] br[427] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_428 bl[428] br[428] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_429 bl[429] br[429] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_430 bl[430] br[430] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_431 bl[431] br[431] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_432 bl[432] br[432] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_433 bl[433] br[433] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_434 bl[434] br[434] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_435 bl[435] br[435] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_436 bl[436] br[436] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_437 bl[437] br[437] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_438 bl[438] br[438] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_439 bl[439] br[439] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_440 bl[440] br[440] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_441 bl[441] br[441] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_442 bl[442] br[442] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_443 bl[443] br[443] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_444 bl[444] br[444] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_445 bl[445] br[445] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_446 bl[446] br[446] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_447 bl[447] br[447] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_448 bl[448] br[448] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_449 bl[449] br[449] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_450 bl[450] br[450] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_451 bl[451] br[451] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_452 bl[452] br[452] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_453 bl[453] br[453] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_454 bl[454] br[454] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_455 bl[455] br[455] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_456 bl[456] br[456] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_457 bl[457] br[457] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_458 bl[458] br[458] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_459 bl[459] br[459] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_460 bl[460] br[460] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_461 bl[461] br[461] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_462 bl[462] br[462] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_463 bl[463] br[463] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_464 bl[464] br[464] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_465 bl[465] br[465] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_466 bl[466] br[466] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_467 bl[467] br[467] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_468 bl[468] br[468] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_469 bl[469] br[469] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_470 bl[470] br[470] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_471 bl[471] br[471] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_472 bl[472] br[472] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_473 bl[473] br[473] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_474 bl[474] br[474] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_475 bl[475] br[475] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_476 bl[476] br[476] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_477 bl[477] br[477] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_478 bl[478] br[478] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_479 bl[479] br[479] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_480 bl[480] br[480] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_481 bl[481] br[481] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_482 bl[482] br[482] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_483 bl[483] br[483] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_484 bl[484] br[484] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_485 bl[485] br[485] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_486 bl[486] br[486] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_487 bl[487] br[487] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_488 bl[488] br[488] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_489 bl[489] br[489] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_490 bl[490] br[490] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_491 bl[491] br[491] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_492 bl[492] br[492] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_493 bl[493] br[493] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_494 bl[494] br[494] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_495 bl[495] br[495] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_496 bl[496] br[496] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_497 bl[497] br[497] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_498 bl[498] br[498] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_499 bl[499] br[499] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_500 bl[500] br[500] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_501 bl[501] br[501] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_502 bl[502] br[502] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_503 bl[503] br[503] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_504 bl[504] br[504] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_505 bl[505] br[505] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_506 bl[506] br[506] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_507 bl[507] br[507] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_508 bl[508] br[508] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_509 bl[509] br[509] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_510 bl[510] br[510] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_51_511 bl[511] br[511] vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xcell_52_0 bl[0] br[0] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_1 bl[1] br[1] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_2 bl[2] br[2] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_3 bl[3] br[3] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_4 bl[4] br[4] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_5 bl[5] br[5] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_6 bl[6] br[6] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_7 bl[7] br[7] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_8 bl[8] br[8] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_9 bl[9] br[9] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_10 bl[10] br[10] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_11 bl[11] br[11] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_12 bl[12] br[12] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_13 bl[13] br[13] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_14 bl[14] br[14] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_15 bl[15] br[15] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_16 bl[16] br[16] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_17 bl[17] br[17] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_18 bl[18] br[18] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_19 bl[19] br[19] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_20 bl[20] br[20] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_21 bl[21] br[21] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_22 bl[22] br[22] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_23 bl[23] br[23] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_24 bl[24] br[24] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_25 bl[25] br[25] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_26 bl[26] br[26] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_27 bl[27] br[27] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_28 bl[28] br[28] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_29 bl[29] br[29] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_30 bl[30] br[30] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_31 bl[31] br[31] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_32 bl[32] br[32] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_33 bl[33] br[33] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_34 bl[34] br[34] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_35 bl[35] br[35] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_36 bl[36] br[36] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_37 bl[37] br[37] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_38 bl[38] br[38] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_39 bl[39] br[39] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_40 bl[40] br[40] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_41 bl[41] br[41] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_42 bl[42] br[42] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_43 bl[43] br[43] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_44 bl[44] br[44] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_45 bl[45] br[45] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_46 bl[46] br[46] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_47 bl[47] br[47] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_48 bl[48] br[48] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_49 bl[49] br[49] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_50 bl[50] br[50] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_51 bl[51] br[51] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_52 bl[52] br[52] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_53 bl[53] br[53] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_54 bl[54] br[54] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_55 bl[55] br[55] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_56 bl[56] br[56] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_57 bl[57] br[57] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_58 bl[58] br[58] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_59 bl[59] br[59] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_60 bl[60] br[60] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_61 bl[61] br[61] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_62 bl[62] br[62] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_63 bl[63] br[63] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_64 bl[64] br[64] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_65 bl[65] br[65] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_66 bl[66] br[66] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_67 bl[67] br[67] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_68 bl[68] br[68] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_69 bl[69] br[69] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_70 bl[70] br[70] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_71 bl[71] br[71] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_72 bl[72] br[72] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_73 bl[73] br[73] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_74 bl[74] br[74] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_75 bl[75] br[75] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_76 bl[76] br[76] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_77 bl[77] br[77] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_78 bl[78] br[78] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_79 bl[79] br[79] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_80 bl[80] br[80] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_81 bl[81] br[81] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_82 bl[82] br[82] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_83 bl[83] br[83] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_84 bl[84] br[84] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_85 bl[85] br[85] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_86 bl[86] br[86] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_87 bl[87] br[87] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_88 bl[88] br[88] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_89 bl[89] br[89] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_90 bl[90] br[90] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_91 bl[91] br[91] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_92 bl[92] br[92] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_93 bl[93] br[93] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_94 bl[94] br[94] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_95 bl[95] br[95] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_96 bl[96] br[96] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_97 bl[97] br[97] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_98 bl[98] br[98] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_99 bl[99] br[99] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_100 bl[100] br[100] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_101 bl[101] br[101] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_102 bl[102] br[102] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_103 bl[103] br[103] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_104 bl[104] br[104] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_105 bl[105] br[105] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_106 bl[106] br[106] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_107 bl[107] br[107] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_108 bl[108] br[108] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_109 bl[109] br[109] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_110 bl[110] br[110] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_111 bl[111] br[111] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_112 bl[112] br[112] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_113 bl[113] br[113] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_114 bl[114] br[114] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_115 bl[115] br[115] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_116 bl[116] br[116] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_117 bl[117] br[117] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_118 bl[118] br[118] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_119 bl[119] br[119] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_120 bl[120] br[120] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_121 bl[121] br[121] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_122 bl[122] br[122] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_123 bl[123] br[123] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_124 bl[124] br[124] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_125 bl[125] br[125] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_126 bl[126] br[126] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_127 bl[127] br[127] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_128 bl[128] br[128] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_129 bl[129] br[129] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_130 bl[130] br[130] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_131 bl[131] br[131] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_132 bl[132] br[132] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_133 bl[133] br[133] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_134 bl[134] br[134] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_135 bl[135] br[135] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_136 bl[136] br[136] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_137 bl[137] br[137] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_138 bl[138] br[138] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_139 bl[139] br[139] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_140 bl[140] br[140] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_141 bl[141] br[141] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_142 bl[142] br[142] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_143 bl[143] br[143] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_144 bl[144] br[144] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_145 bl[145] br[145] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_146 bl[146] br[146] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_147 bl[147] br[147] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_148 bl[148] br[148] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_149 bl[149] br[149] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_150 bl[150] br[150] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_151 bl[151] br[151] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_152 bl[152] br[152] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_153 bl[153] br[153] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_154 bl[154] br[154] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_155 bl[155] br[155] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_156 bl[156] br[156] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_157 bl[157] br[157] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_158 bl[158] br[158] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_159 bl[159] br[159] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_160 bl[160] br[160] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_161 bl[161] br[161] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_162 bl[162] br[162] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_163 bl[163] br[163] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_164 bl[164] br[164] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_165 bl[165] br[165] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_166 bl[166] br[166] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_167 bl[167] br[167] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_168 bl[168] br[168] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_169 bl[169] br[169] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_170 bl[170] br[170] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_171 bl[171] br[171] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_172 bl[172] br[172] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_173 bl[173] br[173] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_174 bl[174] br[174] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_175 bl[175] br[175] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_176 bl[176] br[176] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_177 bl[177] br[177] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_178 bl[178] br[178] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_179 bl[179] br[179] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_180 bl[180] br[180] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_181 bl[181] br[181] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_182 bl[182] br[182] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_183 bl[183] br[183] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_184 bl[184] br[184] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_185 bl[185] br[185] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_186 bl[186] br[186] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_187 bl[187] br[187] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_188 bl[188] br[188] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_189 bl[189] br[189] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_190 bl[190] br[190] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_191 bl[191] br[191] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_192 bl[192] br[192] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_193 bl[193] br[193] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_194 bl[194] br[194] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_195 bl[195] br[195] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_196 bl[196] br[196] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_197 bl[197] br[197] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_198 bl[198] br[198] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_199 bl[199] br[199] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_200 bl[200] br[200] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_201 bl[201] br[201] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_202 bl[202] br[202] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_203 bl[203] br[203] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_204 bl[204] br[204] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_205 bl[205] br[205] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_206 bl[206] br[206] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_207 bl[207] br[207] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_208 bl[208] br[208] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_209 bl[209] br[209] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_210 bl[210] br[210] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_211 bl[211] br[211] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_212 bl[212] br[212] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_213 bl[213] br[213] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_214 bl[214] br[214] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_215 bl[215] br[215] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_216 bl[216] br[216] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_217 bl[217] br[217] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_218 bl[218] br[218] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_219 bl[219] br[219] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_220 bl[220] br[220] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_221 bl[221] br[221] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_222 bl[222] br[222] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_223 bl[223] br[223] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_224 bl[224] br[224] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_225 bl[225] br[225] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_226 bl[226] br[226] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_227 bl[227] br[227] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_228 bl[228] br[228] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_229 bl[229] br[229] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_230 bl[230] br[230] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_231 bl[231] br[231] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_232 bl[232] br[232] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_233 bl[233] br[233] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_234 bl[234] br[234] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_235 bl[235] br[235] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_236 bl[236] br[236] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_237 bl[237] br[237] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_238 bl[238] br[238] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_239 bl[239] br[239] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_240 bl[240] br[240] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_241 bl[241] br[241] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_242 bl[242] br[242] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_243 bl[243] br[243] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_244 bl[244] br[244] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_245 bl[245] br[245] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_246 bl[246] br[246] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_247 bl[247] br[247] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_248 bl[248] br[248] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_249 bl[249] br[249] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_250 bl[250] br[250] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_251 bl[251] br[251] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_252 bl[252] br[252] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_253 bl[253] br[253] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_254 bl[254] br[254] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_255 bl[255] br[255] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_256 bl[256] br[256] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_257 bl[257] br[257] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_258 bl[258] br[258] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_259 bl[259] br[259] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_260 bl[260] br[260] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_261 bl[261] br[261] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_262 bl[262] br[262] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_263 bl[263] br[263] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_264 bl[264] br[264] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_265 bl[265] br[265] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_266 bl[266] br[266] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_267 bl[267] br[267] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_268 bl[268] br[268] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_269 bl[269] br[269] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_270 bl[270] br[270] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_271 bl[271] br[271] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_272 bl[272] br[272] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_273 bl[273] br[273] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_274 bl[274] br[274] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_275 bl[275] br[275] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_276 bl[276] br[276] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_277 bl[277] br[277] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_278 bl[278] br[278] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_279 bl[279] br[279] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_280 bl[280] br[280] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_281 bl[281] br[281] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_282 bl[282] br[282] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_283 bl[283] br[283] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_284 bl[284] br[284] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_285 bl[285] br[285] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_286 bl[286] br[286] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_287 bl[287] br[287] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_288 bl[288] br[288] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_289 bl[289] br[289] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_290 bl[290] br[290] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_291 bl[291] br[291] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_292 bl[292] br[292] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_293 bl[293] br[293] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_294 bl[294] br[294] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_295 bl[295] br[295] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_296 bl[296] br[296] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_297 bl[297] br[297] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_298 bl[298] br[298] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_299 bl[299] br[299] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_300 bl[300] br[300] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_301 bl[301] br[301] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_302 bl[302] br[302] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_303 bl[303] br[303] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_304 bl[304] br[304] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_305 bl[305] br[305] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_306 bl[306] br[306] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_307 bl[307] br[307] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_308 bl[308] br[308] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_309 bl[309] br[309] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_310 bl[310] br[310] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_311 bl[311] br[311] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_312 bl[312] br[312] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_313 bl[313] br[313] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_314 bl[314] br[314] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_315 bl[315] br[315] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_316 bl[316] br[316] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_317 bl[317] br[317] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_318 bl[318] br[318] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_319 bl[319] br[319] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_320 bl[320] br[320] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_321 bl[321] br[321] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_322 bl[322] br[322] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_323 bl[323] br[323] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_324 bl[324] br[324] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_325 bl[325] br[325] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_326 bl[326] br[326] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_327 bl[327] br[327] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_328 bl[328] br[328] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_329 bl[329] br[329] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_330 bl[330] br[330] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_331 bl[331] br[331] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_332 bl[332] br[332] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_333 bl[333] br[333] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_334 bl[334] br[334] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_335 bl[335] br[335] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_336 bl[336] br[336] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_337 bl[337] br[337] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_338 bl[338] br[338] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_339 bl[339] br[339] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_340 bl[340] br[340] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_341 bl[341] br[341] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_342 bl[342] br[342] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_343 bl[343] br[343] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_344 bl[344] br[344] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_345 bl[345] br[345] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_346 bl[346] br[346] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_347 bl[347] br[347] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_348 bl[348] br[348] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_349 bl[349] br[349] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_350 bl[350] br[350] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_351 bl[351] br[351] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_352 bl[352] br[352] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_353 bl[353] br[353] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_354 bl[354] br[354] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_355 bl[355] br[355] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_356 bl[356] br[356] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_357 bl[357] br[357] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_358 bl[358] br[358] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_359 bl[359] br[359] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_360 bl[360] br[360] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_361 bl[361] br[361] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_362 bl[362] br[362] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_363 bl[363] br[363] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_364 bl[364] br[364] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_365 bl[365] br[365] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_366 bl[366] br[366] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_367 bl[367] br[367] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_368 bl[368] br[368] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_369 bl[369] br[369] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_370 bl[370] br[370] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_371 bl[371] br[371] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_372 bl[372] br[372] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_373 bl[373] br[373] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_374 bl[374] br[374] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_375 bl[375] br[375] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_376 bl[376] br[376] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_377 bl[377] br[377] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_378 bl[378] br[378] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_379 bl[379] br[379] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_380 bl[380] br[380] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_381 bl[381] br[381] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_382 bl[382] br[382] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_383 bl[383] br[383] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_384 bl[384] br[384] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_385 bl[385] br[385] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_386 bl[386] br[386] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_387 bl[387] br[387] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_388 bl[388] br[388] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_389 bl[389] br[389] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_390 bl[390] br[390] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_391 bl[391] br[391] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_392 bl[392] br[392] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_393 bl[393] br[393] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_394 bl[394] br[394] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_395 bl[395] br[395] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_396 bl[396] br[396] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_397 bl[397] br[397] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_398 bl[398] br[398] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_399 bl[399] br[399] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_400 bl[400] br[400] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_401 bl[401] br[401] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_402 bl[402] br[402] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_403 bl[403] br[403] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_404 bl[404] br[404] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_405 bl[405] br[405] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_406 bl[406] br[406] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_407 bl[407] br[407] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_408 bl[408] br[408] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_409 bl[409] br[409] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_410 bl[410] br[410] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_411 bl[411] br[411] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_412 bl[412] br[412] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_413 bl[413] br[413] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_414 bl[414] br[414] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_415 bl[415] br[415] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_416 bl[416] br[416] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_417 bl[417] br[417] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_418 bl[418] br[418] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_419 bl[419] br[419] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_420 bl[420] br[420] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_421 bl[421] br[421] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_422 bl[422] br[422] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_423 bl[423] br[423] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_424 bl[424] br[424] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_425 bl[425] br[425] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_426 bl[426] br[426] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_427 bl[427] br[427] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_428 bl[428] br[428] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_429 bl[429] br[429] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_430 bl[430] br[430] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_431 bl[431] br[431] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_432 bl[432] br[432] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_433 bl[433] br[433] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_434 bl[434] br[434] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_435 bl[435] br[435] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_436 bl[436] br[436] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_437 bl[437] br[437] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_438 bl[438] br[438] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_439 bl[439] br[439] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_440 bl[440] br[440] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_441 bl[441] br[441] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_442 bl[442] br[442] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_443 bl[443] br[443] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_444 bl[444] br[444] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_445 bl[445] br[445] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_446 bl[446] br[446] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_447 bl[447] br[447] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_448 bl[448] br[448] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_449 bl[449] br[449] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_450 bl[450] br[450] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_451 bl[451] br[451] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_452 bl[452] br[452] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_453 bl[453] br[453] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_454 bl[454] br[454] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_455 bl[455] br[455] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_456 bl[456] br[456] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_457 bl[457] br[457] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_458 bl[458] br[458] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_459 bl[459] br[459] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_460 bl[460] br[460] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_461 bl[461] br[461] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_462 bl[462] br[462] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_463 bl[463] br[463] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_464 bl[464] br[464] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_465 bl[465] br[465] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_466 bl[466] br[466] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_467 bl[467] br[467] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_468 bl[468] br[468] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_469 bl[469] br[469] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_470 bl[470] br[470] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_471 bl[471] br[471] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_472 bl[472] br[472] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_473 bl[473] br[473] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_474 bl[474] br[474] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_475 bl[475] br[475] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_476 bl[476] br[476] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_477 bl[477] br[477] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_478 bl[478] br[478] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_479 bl[479] br[479] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_480 bl[480] br[480] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_481 bl[481] br[481] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_482 bl[482] br[482] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_483 bl[483] br[483] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_484 bl[484] br[484] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_485 bl[485] br[485] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_486 bl[486] br[486] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_487 bl[487] br[487] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_488 bl[488] br[488] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_489 bl[489] br[489] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_490 bl[490] br[490] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_491 bl[491] br[491] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_492 bl[492] br[492] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_493 bl[493] br[493] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_494 bl[494] br[494] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_495 bl[495] br[495] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_496 bl[496] br[496] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_497 bl[497] br[497] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_498 bl[498] br[498] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_499 bl[499] br[499] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_500 bl[500] br[500] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_501 bl[501] br[501] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_502 bl[502] br[502] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_503 bl[503] br[503] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_504 bl[504] br[504] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_505 bl[505] br[505] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_506 bl[506] br[506] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_507 bl[507] br[507] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_508 bl[508] br[508] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_509 bl[509] br[509] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_510 bl[510] br[510] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_52_511 bl[511] br[511] vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xcell_53_0 bl[0] br[0] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_1 bl[1] br[1] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_2 bl[2] br[2] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_3 bl[3] br[3] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_4 bl[4] br[4] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_5 bl[5] br[5] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_6 bl[6] br[6] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_7 bl[7] br[7] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_8 bl[8] br[8] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_9 bl[9] br[9] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_10 bl[10] br[10] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_11 bl[11] br[11] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_12 bl[12] br[12] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_13 bl[13] br[13] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_14 bl[14] br[14] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_15 bl[15] br[15] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_16 bl[16] br[16] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_17 bl[17] br[17] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_18 bl[18] br[18] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_19 bl[19] br[19] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_20 bl[20] br[20] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_21 bl[21] br[21] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_22 bl[22] br[22] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_23 bl[23] br[23] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_24 bl[24] br[24] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_25 bl[25] br[25] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_26 bl[26] br[26] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_27 bl[27] br[27] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_28 bl[28] br[28] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_29 bl[29] br[29] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_30 bl[30] br[30] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_31 bl[31] br[31] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_32 bl[32] br[32] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_33 bl[33] br[33] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_34 bl[34] br[34] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_35 bl[35] br[35] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_36 bl[36] br[36] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_37 bl[37] br[37] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_38 bl[38] br[38] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_39 bl[39] br[39] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_40 bl[40] br[40] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_41 bl[41] br[41] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_42 bl[42] br[42] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_43 bl[43] br[43] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_44 bl[44] br[44] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_45 bl[45] br[45] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_46 bl[46] br[46] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_47 bl[47] br[47] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_48 bl[48] br[48] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_49 bl[49] br[49] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_50 bl[50] br[50] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_51 bl[51] br[51] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_52 bl[52] br[52] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_53 bl[53] br[53] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_54 bl[54] br[54] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_55 bl[55] br[55] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_56 bl[56] br[56] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_57 bl[57] br[57] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_58 bl[58] br[58] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_59 bl[59] br[59] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_60 bl[60] br[60] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_61 bl[61] br[61] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_62 bl[62] br[62] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_63 bl[63] br[63] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_64 bl[64] br[64] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_65 bl[65] br[65] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_66 bl[66] br[66] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_67 bl[67] br[67] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_68 bl[68] br[68] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_69 bl[69] br[69] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_70 bl[70] br[70] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_71 bl[71] br[71] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_72 bl[72] br[72] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_73 bl[73] br[73] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_74 bl[74] br[74] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_75 bl[75] br[75] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_76 bl[76] br[76] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_77 bl[77] br[77] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_78 bl[78] br[78] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_79 bl[79] br[79] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_80 bl[80] br[80] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_81 bl[81] br[81] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_82 bl[82] br[82] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_83 bl[83] br[83] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_84 bl[84] br[84] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_85 bl[85] br[85] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_86 bl[86] br[86] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_87 bl[87] br[87] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_88 bl[88] br[88] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_89 bl[89] br[89] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_90 bl[90] br[90] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_91 bl[91] br[91] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_92 bl[92] br[92] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_93 bl[93] br[93] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_94 bl[94] br[94] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_95 bl[95] br[95] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_96 bl[96] br[96] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_97 bl[97] br[97] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_98 bl[98] br[98] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_99 bl[99] br[99] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_100 bl[100] br[100] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_101 bl[101] br[101] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_102 bl[102] br[102] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_103 bl[103] br[103] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_104 bl[104] br[104] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_105 bl[105] br[105] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_106 bl[106] br[106] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_107 bl[107] br[107] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_108 bl[108] br[108] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_109 bl[109] br[109] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_110 bl[110] br[110] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_111 bl[111] br[111] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_112 bl[112] br[112] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_113 bl[113] br[113] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_114 bl[114] br[114] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_115 bl[115] br[115] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_116 bl[116] br[116] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_117 bl[117] br[117] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_118 bl[118] br[118] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_119 bl[119] br[119] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_120 bl[120] br[120] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_121 bl[121] br[121] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_122 bl[122] br[122] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_123 bl[123] br[123] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_124 bl[124] br[124] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_125 bl[125] br[125] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_126 bl[126] br[126] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_127 bl[127] br[127] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_128 bl[128] br[128] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_129 bl[129] br[129] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_130 bl[130] br[130] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_131 bl[131] br[131] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_132 bl[132] br[132] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_133 bl[133] br[133] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_134 bl[134] br[134] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_135 bl[135] br[135] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_136 bl[136] br[136] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_137 bl[137] br[137] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_138 bl[138] br[138] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_139 bl[139] br[139] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_140 bl[140] br[140] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_141 bl[141] br[141] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_142 bl[142] br[142] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_143 bl[143] br[143] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_144 bl[144] br[144] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_145 bl[145] br[145] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_146 bl[146] br[146] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_147 bl[147] br[147] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_148 bl[148] br[148] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_149 bl[149] br[149] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_150 bl[150] br[150] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_151 bl[151] br[151] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_152 bl[152] br[152] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_153 bl[153] br[153] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_154 bl[154] br[154] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_155 bl[155] br[155] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_156 bl[156] br[156] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_157 bl[157] br[157] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_158 bl[158] br[158] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_159 bl[159] br[159] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_160 bl[160] br[160] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_161 bl[161] br[161] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_162 bl[162] br[162] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_163 bl[163] br[163] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_164 bl[164] br[164] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_165 bl[165] br[165] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_166 bl[166] br[166] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_167 bl[167] br[167] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_168 bl[168] br[168] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_169 bl[169] br[169] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_170 bl[170] br[170] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_171 bl[171] br[171] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_172 bl[172] br[172] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_173 bl[173] br[173] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_174 bl[174] br[174] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_175 bl[175] br[175] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_176 bl[176] br[176] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_177 bl[177] br[177] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_178 bl[178] br[178] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_179 bl[179] br[179] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_180 bl[180] br[180] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_181 bl[181] br[181] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_182 bl[182] br[182] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_183 bl[183] br[183] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_184 bl[184] br[184] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_185 bl[185] br[185] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_186 bl[186] br[186] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_187 bl[187] br[187] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_188 bl[188] br[188] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_189 bl[189] br[189] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_190 bl[190] br[190] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_191 bl[191] br[191] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_192 bl[192] br[192] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_193 bl[193] br[193] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_194 bl[194] br[194] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_195 bl[195] br[195] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_196 bl[196] br[196] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_197 bl[197] br[197] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_198 bl[198] br[198] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_199 bl[199] br[199] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_200 bl[200] br[200] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_201 bl[201] br[201] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_202 bl[202] br[202] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_203 bl[203] br[203] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_204 bl[204] br[204] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_205 bl[205] br[205] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_206 bl[206] br[206] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_207 bl[207] br[207] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_208 bl[208] br[208] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_209 bl[209] br[209] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_210 bl[210] br[210] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_211 bl[211] br[211] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_212 bl[212] br[212] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_213 bl[213] br[213] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_214 bl[214] br[214] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_215 bl[215] br[215] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_216 bl[216] br[216] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_217 bl[217] br[217] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_218 bl[218] br[218] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_219 bl[219] br[219] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_220 bl[220] br[220] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_221 bl[221] br[221] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_222 bl[222] br[222] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_223 bl[223] br[223] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_224 bl[224] br[224] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_225 bl[225] br[225] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_226 bl[226] br[226] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_227 bl[227] br[227] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_228 bl[228] br[228] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_229 bl[229] br[229] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_230 bl[230] br[230] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_231 bl[231] br[231] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_232 bl[232] br[232] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_233 bl[233] br[233] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_234 bl[234] br[234] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_235 bl[235] br[235] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_236 bl[236] br[236] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_237 bl[237] br[237] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_238 bl[238] br[238] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_239 bl[239] br[239] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_240 bl[240] br[240] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_241 bl[241] br[241] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_242 bl[242] br[242] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_243 bl[243] br[243] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_244 bl[244] br[244] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_245 bl[245] br[245] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_246 bl[246] br[246] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_247 bl[247] br[247] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_248 bl[248] br[248] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_249 bl[249] br[249] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_250 bl[250] br[250] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_251 bl[251] br[251] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_252 bl[252] br[252] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_253 bl[253] br[253] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_254 bl[254] br[254] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_255 bl[255] br[255] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_256 bl[256] br[256] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_257 bl[257] br[257] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_258 bl[258] br[258] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_259 bl[259] br[259] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_260 bl[260] br[260] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_261 bl[261] br[261] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_262 bl[262] br[262] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_263 bl[263] br[263] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_264 bl[264] br[264] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_265 bl[265] br[265] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_266 bl[266] br[266] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_267 bl[267] br[267] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_268 bl[268] br[268] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_269 bl[269] br[269] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_270 bl[270] br[270] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_271 bl[271] br[271] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_272 bl[272] br[272] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_273 bl[273] br[273] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_274 bl[274] br[274] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_275 bl[275] br[275] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_276 bl[276] br[276] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_277 bl[277] br[277] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_278 bl[278] br[278] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_279 bl[279] br[279] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_280 bl[280] br[280] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_281 bl[281] br[281] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_282 bl[282] br[282] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_283 bl[283] br[283] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_284 bl[284] br[284] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_285 bl[285] br[285] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_286 bl[286] br[286] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_287 bl[287] br[287] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_288 bl[288] br[288] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_289 bl[289] br[289] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_290 bl[290] br[290] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_291 bl[291] br[291] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_292 bl[292] br[292] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_293 bl[293] br[293] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_294 bl[294] br[294] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_295 bl[295] br[295] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_296 bl[296] br[296] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_297 bl[297] br[297] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_298 bl[298] br[298] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_299 bl[299] br[299] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_300 bl[300] br[300] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_301 bl[301] br[301] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_302 bl[302] br[302] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_303 bl[303] br[303] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_304 bl[304] br[304] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_305 bl[305] br[305] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_306 bl[306] br[306] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_307 bl[307] br[307] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_308 bl[308] br[308] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_309 bl[309] br[309] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_310 bl[310] br[310] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_311 bl[311] br[311] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_312 bl[312] br[312] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_313 bl[313] br[313] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_314 bl[314] br[314] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_315 bl[315] br[315] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_316 bl[316] br[316] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_317 bl[317] br[317] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_318 bl[318] br[318] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_319 bl[319] br[319] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_320 bl[320] br[320] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_321 bl[321] br[321] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_322 bl[322] br[322] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_323 bl[323] br[323] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_324 bl[324] br[324] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_325 bl[325] br[325] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_326 bl[326] br[326] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_327 bl[327] br[327] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_328 bl[328] br[328] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_329 bl[329] br[329] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_330 bl[330] br[330] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_331 bl[331] br[331] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_332 bl[332] br[332] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_333 bl[333] br[333] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_334 bl[334] br[334] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_335 bl[335] br[335] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_336 bl[336] br[336] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_337 bl[337] br[337] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_338 bl[338] br[338] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_339 bl[339] br[339] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_340 bl[340] br[340] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_341 bl[341] br[341] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_342 bl[342] br[342] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_343 bl[343] br[343] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_344 bl[344] br[344] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_345 bl[345] br[345] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_346 bl[346] br[346] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_347 bl[347] br[347] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_348 bl[348] br[348] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_349 bl[349] br[349] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_350 bl[350] br[350] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_351 bl[351] br[351] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_352 bl[352] br[352] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_353 bl[353] br[353] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_354 bl[354] br[354] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_355 bl[355] br[355] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_356 bl[356] br[356] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_357 bl[357] br[357] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_358 bl[358] br[358] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_359 bl[359] br[359] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_360 bl[360] br[360] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_361 bl[361] br[361] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_362 bl[362] br[362] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_363 bl[363] br[363] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_364 bl[364] br[364] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_365 bl[365] br[365] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_366 bl[366] br[366] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_367 bl[367] br[367] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_368 bl[368] br[368] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_369 bl[369] br[369] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_370 bl[370] br[370] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_371 bl[371] br[371] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_372 bl[372] br[372] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_373 bl[373] br[373] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_374 bl[374] br[374] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_375 bl[375] br[375] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_376 bl[376] br[376] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_377 bl[377] br[377] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_378 bl[378] br[378] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_379 bl[379] br[379] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_380 bl[380] br[380] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_381 bl[381] br[381] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_382 bl[382] br[382] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_383 bl[383] br[383] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_384 bl[384] br[384] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_385 bl[385] br[385] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_386 bl[386] br[386] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_387 bl[387] br[387] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_388 bl[388] br[388] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_389 bl[389] br[389] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_390 bl[390] br[390] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_391 bl[391] br[391] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_392 bl[392] br[392] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_393 bl[393] br[393] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_394 bl[394] br[394] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_395 bl[395] br[395] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_396 bl[396] br[396] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_397 bl[397] br[397] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_398 bl[398] br[398] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_399 bl[399] br[399] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_400 bl[400] br[400] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_401 bl[401] br[401] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_402 bl[402] br[402] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_403 bl[403] br[403] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_404 bl[404] br[404] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_405 bl[405] br[405] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_406 bl[406] br[406] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_407 bl[407] br[407] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_408 bl[408] br[408] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_409 bl[409] br[409] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_410 bl[410] br[410] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_411 bl[411] br[411] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_412 bl[412] br[412] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_413 bl[413] br[413] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_414 bl[414] br[414] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_415 bl[415] br[415] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_416 bl[416] br[416] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_417 bl[417] br[417] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_418 bl[418] br[418] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_419 bl[419] br[419] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_420 bl[420] br[420] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_421 bl[421] br[421] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_422 bl[422] br[422] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_423 bl[423] br[423] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_424 bl[424] br[424] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_425 bl[425] br[425] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_426 bl[426] br[426] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_427 bl[427] br[427] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_428 bl[428] br[428] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_429 bl[429] br[429] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_430 bl[430] br[430] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_431 bl[431] br[431] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_432 bl[432] br[432] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_433 bl[433] br[433] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_434 bl[434] br[434] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_435 bl[435] br[435] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_436 bl[436] br[436] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_437 bl[437] br[437] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_438 bl[438] br[438] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_439 bl[439] br[439] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_440 bl[440] br[440] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_441 bl[441] br[441] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_442 bl[442] br[442] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_443 bl[443] br[443] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_444 bl[444] br[444] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_445 bl[445] br[445] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_446 bl[446] br[446] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_447 bl[447] br[447] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_448 bl[448] br[448] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_449 bl[449] br[449] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_450 bl[450] br[450] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_451 bl[451] br[451] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_452 bl[452] br[452] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_453 bl[453] br[453] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_454 bl[454] br[454] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_455 bl[455] br[455] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_456 bl[456] br[456] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_457 bl[457] br[457] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_458 bl[458] br[458] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_459 bl[459] br[459] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_460 bl[460] br[460] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_461 bl[461] br[461] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_462 bl[462] br[462] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_463 bl[463] br[463] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_464 bl[464] br[464] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_465 bl[465] br[465] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_466 bl[466] br[466] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_467 bl[467] br[467] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_468 bl[468] br[468] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_469 bl[469] br[469] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_470 bl[470] br[470] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_471 bl[471] br[471] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_472 bl[472] br[472] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_473 bl[473] br[473] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_474 bl[474] br[474] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_475 bl[475] br[475] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_476 bl[476] br[476] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_477 bl[477] br[477] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_478 bl[478] br[478] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_479 bl[479] br[479] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_480 bl[480] br[480] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_481 bl[481] br[481] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_482 bl[482] br[482] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_483 bl[483] br[483] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_484 bl[484] br[484] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_485 bl[485] br[485] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_486 bl[486] br[486] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_487 bl[487] br[487] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_488 bl[488] br[488] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_489 bl[489] br[489] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_490 bl[490] br[490] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_491 bl[491] br[491] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_492 bl[492] br[492] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_493 bl[493] br[493] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_494 bl[494] br[494] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_495 bl[495] br[495] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_496 bl[496] br[496] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_497 bl[497] br[497] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_498 bl[498] br[498] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_499 bl[499] br[499] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_500 bl[500] br[500] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_501 bl[501] br[501] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_502 bl[502] br[502] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_503 bl[503] br[503] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_504 bl[504] br[504] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_505 bl[505] br[505] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_506 bl[506] br[506] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_507 bl[507] br[507] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_508 bl[508] br[508] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_509 bl[509] br[509] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_510 bl[510] br[510] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_53_511 bl[511] br[511] vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xcell_54_0 bl[0] br[0] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_1 bl[1] br[1] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_2 bl[2] br[2] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_3 bl[3] br[3] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_4 bl[4] br[4] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_5 bl[5] br[5] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_6 bl[6] br[6] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_7 bl[7] br[7] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_8 bl[8] br[8] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_9 bl[9] br[9] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_10 bl[10] br[10] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_11 bl[11] br[11] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_12 bl[12] br[12] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_13 bl[13] br[13] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_14 bl[14] br[14] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_15 bl[15] br[15] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_16 bl[16] br[16] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_17 bl[17] br[17] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_18 bl[18] br[18] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_19 bl[19] br[19] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_20 bl[20] br[20] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_21 bl[21] br[21] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_22 bl[22] br[22] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_23 bl[23] br[23] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_24 bl[24] br[24] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_25 bl[25] br[25] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_26 bl[26] br[26] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_27 bl[27] br[27] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_28 bl[28] br[28] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_29 bl[29] br[29] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_30 bl[30] br[30] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_31 bl[31] br[31] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_32 bl[32] br[32] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_33 bl[33] br[33] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_34 bl[34] br[34] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_35 bl[35] br[35] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_36 bl[36] br[36] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_37 bl[37] br[37] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_38 bl[38] br[38] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_39 bl[39] br[39] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_40 bl[40] br[40] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_41 bl[41] br[41] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_42 bl[42] br[42] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_43 bl[43] br[43] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_44 bl[44] br[44] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_45 bl[45] br[45] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_46 bl[46] br[46] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_47 bl[47] br[47] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_48 bl[48] br[48] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_49 bl[49] br[49] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_50 bl[50] br[50] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_51 bl[51] br[51] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_52 bl[52] br[52] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_53 bl[53] br[53] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_54 bl[54] br[54] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_55 bl[55] br[55] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_56 bl[56] br[56] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_57 bl[57] br[57] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_58 bl[58] br[58] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_59 bl[59] br[59] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_60 bl[60] br[60] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_61 bl[61] br[61] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_62 bl[62] br[62] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_63 bl[63] br[63] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_64 bl[64] br[64] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_65 bl[65] br[65] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_66 bl[66] br[66] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_67 bl[67] br[67] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_68 bl[68] br[68] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_69 bl[69] br[69] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_70 bl[70] br[70] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_71 bl[71] br[71] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_72 bl[72] br[72] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_73 bl[73] br[73] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_74 bl[74] br[74] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_75 bl[75] br[75] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_76 bl[76] br[76] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_77 bl[77] br[77] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_78 bl[78] br[78] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_79 bl[79] br[79] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_80 bl[80] br[80] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_81 bl[81] br[81] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_82 bl[82] br[82] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_83 bl[83] br[83] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_84 bl[84] br[84] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_85 bl[85] br[85] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_86 bl[86] br[86] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_87 bl[87] br[87] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_88 bl[88] br[88] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_89 bl[89] br[89] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_90 bl[90] br[90] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_91 bl[91] br[91] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_92 bl[92] br[92] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_93 bl[93] br[93] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_94 bl[94] br[94] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_95 bl[95] br[95] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_96 bl[96] br[96] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_97 bl[97] br[97] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_98 bl[98] br[98] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_99 bl[99] br[99] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_100 bl[100] br[100] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_101 bl[101] br[101] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_102 bl[102] br[102] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_103 bl[103] br[103] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_104 bl[104] br[104] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_105 bl[105] br[105] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_106 bl[106] br[106] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_107 bl[107] br[107] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_108 bl[108] br[108] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_109 bl[109] br[109] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_110 bl[110] br[110] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_111 bl[111] br[111] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_112 bl[112] br[112] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_113 bl[113] br[113] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_114 bl[114] br[114] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_115 bl[115] br[115] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_116 bl[116] br[116] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_117 bl[117] br[117] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_118 bl[118] br[118] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_119 bl[119] br[119] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_120 bl[120] br[120] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_121 bl[121] br[121] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_122 bl[122] br[122] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_123 bl[123] br[123] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_124 bl[124] br[124] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_125 bl[125] br[125] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_126 bl[126] br[126] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_127 bl[127] br[127] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_128 bl[128] br[128] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_129 bl[129] br[129] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_130 bl[130] br[130] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_131 bl[131] br[131] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_132 bl[132] br[132] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_133 bl[133] br[133] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_134 bl[134] br[134] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_135 bl[135] br[135] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_136 bl[136] br[136] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_137 bl[137] br[137] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_138 bl[138] br[138] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_139 bl[139] br[139] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_140 bl[140] br[140] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_141 bl[141] br[141] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_142 bl[142] br[142] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_143 bl[143] br[143] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_144 bl[144] br[144] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_145 bl[145] br[145] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_146 bl[146] br[146] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_147 bl[147] br[147] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_148 bl[148] br[148] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_149 bl[149] br[149] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_150 bl[150] br[150] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_151 bl[151] br[151] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_152 bl[152] br[152] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_153 bl[153] br[153] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_154 bl[154] br[154] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_155 bl[155] br[155] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_156 bl[156] br[156] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_157 bl[157] br[157] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_158 bl[158] br[158] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_159 bl[159] br[159] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_160 bl[160] br[160] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_161 bl[161] br[161] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_162 bl[162] br[162] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_163 bl[163] br[163] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_164 bl[164] br[164] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_165 bl[165] br[165] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_166 bl[166] br[166] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_167 bl[167] br[167] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_168 bl[168] br[168] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_169 bl[169] br[169] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_170 bl[170] br[170] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_171 bl[171] br[171] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_172 bl[172] br[172] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_173 bl[173] br[173] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_174 bl[174] br[174] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_175 bl[175] br[175] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_176 bl[176] br[176] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_177 bl[177] br[177] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_178 bl[178] br[178] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_179 bl[179] br[179] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_180 bl[180] br[180] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_181 bl[181] br[181] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_182 bl[182] br[182] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_183 bl[183] br[183] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_184 bl[184] br[184] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_185 bl[185] br[185] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_186 bl[186] br[186] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_187 bl[187] br[187] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_188 bl[188] br[188] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_189 bl[189] br[189] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_190 bl[190] br[190] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_191 bl[191] br[191] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_192 bl[192] br[192] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_193 bl[193] br[193] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_194 bl[194] br[194] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_195 bl[195] br[195] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_196 bl[196] br[196] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_197 bl[197] br[197] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_198 bl[198] br[198] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_199 bl[199] br[199] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_200 bl[200] br[200] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_201 bl[201] br[201] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_202 bl[202] br[202] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_203 bl[203] br[203] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_204 bl[204] br[204] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_205 bl[205] br[205] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_206 bl[206] br[206] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_207 bl[207] br[207] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_208 bl[208] br[208] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_209 bl[209] br[209] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_210 bl[210] br[210] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_211 bl[211] br[211] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_212 bl[212] br[212] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_213 bl[213] br[213] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_214 bl[214] br[214] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_215 bl[215] br[215] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_216 bl[216] br[216] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_217 bl[217] br[217] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_218 bl[218] br[218] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_219 bl[219] br[219] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_220 bl[220] br[220] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_221 bl[221] br[221] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_222 bl[222] br[222] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_223 bl[223] br[223] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_224 bl[224] br[224] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_225 bl[225] br[225] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_226 bl[226] br[226] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_227 bl[227] br[227] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_228 bl[228] br[228] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_229 bl[229] br[229] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_230 bl[230] br[230] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_231 bl[231] br[231] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_232 bl[232] br[232] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_233 bl[233] br[233] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_234 bl[234] br[234] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_235 bl[235] br[235] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_236 bl[236] br[236] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_237 bl[237] br[237] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_238 bl[238] br[238] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_239 bl[239] br[239] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_240 bl[240] br[240] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_241 bl[241] br[241] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_242 bl[242] br[242] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_243 bl[243] br[243] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_244 bl[244] br[244] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_245 bl[245] br[245] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_246 bl[246] br[246] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_247 bl[247] br[247] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_248 bl[248] br[248] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_249 bl[249] br[249] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_250 bl[250] br[250] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_251 bl[251] br[251] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_252 bl[252] br[252] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_253 bl[253] br[253] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_254 bl[254] br[254] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_255 bl[255] br[255] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_256 bl[256] br[256] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_257 bl[257] br[257] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_258 bl[258] br[258] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_259 bl[259] br[259] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_260 bl[260] br[260] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_261 bl[261] br[261] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_262 bl[262] br[262] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_263 bl[263] br[263] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_264 bl[264] br[264] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_265 bl[265] br[265] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_266 bl[266] br[266] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_267 bl[267] br[267] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_268 bl[268] br[268] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_269 bl[269] br[269] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_270 bl[270] br[270] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_271 bl[271] br[271] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_272 bl[272] br[272] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_273 bl[273] br[273] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_274 bl[274] br[274] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_275 bl[275] br[275] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_276 bl[276] br[276] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_277 bl[277] br[277] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_278 bl[278] br[278] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_279 bl[279] br[279] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_280 bl[280] br[280] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_281 bl[281] br[281] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_282 bl[282] br[282] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_283 bl[283] br[283] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_284 bl[284] br[284] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_285 bl[285] br[285] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_286 bl[286] br[286] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_287 bl[287] br[287] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_288 bl[288] br[288] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_289 bl[289] br[289] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_290 bl[290] br[290] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_291 bl[291] br[291] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_292 bl[292] br[292] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_293 bl[293] br[293] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_294 bl[294] br[294] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_295 bl[295] br[295] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_296 bl[296] br[296] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_297 bl[297] br[297] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_298 bl[298] br[298] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_299 bl[299] br[299] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_300 bl[300] br[300] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_301 bl[301] br[301] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_302 bl[302] br[302] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_303 bl[303] br[303] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_304 bl[304] br[304] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_305 bl[305] br[305] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_306 bl[306] br[306] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_307 bl[307] br[307] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_308 bl[308] br[308] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_309 bl[309] br[309] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_310 bl[310] br[310] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_311 bl[311] br[311] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_312 bl[312] br[312] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_313 bl[313] br[313] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_314 bl[314] br[314] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_315 bl[315] br[315] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_316 bl[316] br[316] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_317 bl[317] br[317] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_318 bl[318] br[318] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_319 bl[319] br[319] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_320 bl[320] br[320] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_321 bl[321] br[321] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_322 bl[322] br[322] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_323 bl[323] br[323] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_324 bl[324] br[324] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_325 bl[325] br[325] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_326 bl[326] br[326] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_327 bl[327] br[327] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_328 bl[328] br[328] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_329 bl[329] br[329] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_330 bl[330] br[330] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_331 bl[331] br[331] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_332 bl[332] br[332] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_333 bl[333] br[333] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_334 bl[334] br[334] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_335 bl[335] br[335] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_336 bl[336] br[336] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_337 bl[337] br[337] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_338 bl[338] br[338] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_339 bl[339] br[339] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_340 bl[340] br[340] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_341 bl[341] br[341] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_342 bl[342] br[342] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_343 bl[343] br[343] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_344 bl[344] br[344] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_345 bl[345] br[345] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_346 bl[346] br[346] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_347 bl[347] br[347] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_348 bl[348] br[348] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_349 bl[349] br[349] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_350 bl[350] br[350] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_351 bl[351] br[351] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_352 bl[352] br[352] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_353 bl[353] br[353] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_354 bl[354] br[354] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_355 bl[355] br[355] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_356 bl[356] br[356] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_357 bl[357] br[357] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_358 bl[358] br[358] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_359 bl[359] br[359] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_360 bl[360] br[360] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_361 bl[361] br[361] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_362 bl[362] br[362] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_363 bl[363] br[363] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_364 bl[364] br[364] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_365 bl[365] br[365] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_366 bl[366] br[366] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_367 bl[367] br[367] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_368 bl[368] br[368] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_369 bl[369] br[369] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_370 bl[370] br[370] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_371 bl[371] br[371] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_372 bl[372] br[372] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_373 bl[373] br[373] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_374 bl[374] br[374] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_375 bl[375] br[375] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_376 bl[376] br[376] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_377 bl[377] br[377] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_378 bl[378] br[378] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_379 bl[379] br[379] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_380 bl[380] br[380] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_381 bl[381] br[381] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_382 bl[382] br[382] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_383 bl[383] br[383] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_384 bl[384] br[384] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_385 bl[385] br[385] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_386 bl[386] br[386] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_387 bl[387] br[387] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_388 bl[388] br[388] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_389 bl[389] br[389] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_390 bl[390] br[390] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_391 bl[391] br[391] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_392 bl[392] br[392] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_393 bl[393] br[393] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_394 bl[394] br[394] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_395 bl[395] br[395] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_396 bl[396] br[396] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_397 bl[397] br[397] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_398 bl[398] br[398] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_399 bl[399] br[399] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_400 bl[400] br[400] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_401 bl[401] br[401] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_402 bl[402] br[402] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_403 bl[403] br[403] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_404 bl[404] br[404] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_405 bl[405] br[405] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_406 bl[406] br[406] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_407 bl[407] br[407] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_408 bl[408] br[408] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_409 bl[409] br[409] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_410 bl[410] br[410] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_411 bl[411] br[411] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_412 bl[412] br[412] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_413 bl[413] br[413] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_414 bl[414] br[414] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_415 bl[415] br[415] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_416 bl[416] br[416] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_417 bl[417] br[417] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_418 bl[418] br[418] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_419 bl[419] br[419] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_420 bl[420] br[420] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_421 bl[421] br[421] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_422 bl[422] br[422] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_423 bl[423] br[423] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_424 bl[424] br[424] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_425 bl[425] br[425] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_426 bl[426] br[426] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_427 bl[427] br[427] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_428 bl[428] br[428] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_429 bl[429] br[429] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_430 bl[430] br[430] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_431 bl[431] br[431] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_432 bl[432] br[432] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_433 bl[433] br[433] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_434 bl[434] br[434] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_435 bl[435] br[435] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_436 bl[436] br[436] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_437 bl[437] br[437] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_438 bl[438] br[438] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_439 bl[439] br[439] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_440 bl[440] br[440] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_441 bl[441] br[441] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_442 bl[442] br[442] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_443 bl[443] br[443] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_444 bl[444] br[444] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_445 bl[445] br[445] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_446 bl[446] br[446] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_447 bl[447] br[447] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_448 bl[448] br[448] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_449 bl[449] br[449] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_450 bl[450] br[450] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_451 bl[451] br[451] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_452 bl[452] br[452] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_453 bl[453] br[453] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_454 bl[454] br[454] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_455 bl[455] br[455] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_456 bl[456] br[456] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_457 bl[457] br[457] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_458 bl[458] br[458] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_459 bl[459] br[459] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_460 bl[460] br[460] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_461 bl[461] br[461] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_462 bl[462] br[462] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_463 bl[463] br[463] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_464 bl[464] br[464] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_465 bl[465] br[465] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_466 bl[466] br[466] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_467 bl[467] br[467] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_468 bl[468] br[468] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_469 bl[469] br[469] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_470 bl[470] br[470] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_471 bl[471] br[471] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_472 bl[472] br[472] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_473 bl[473] br[473] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_474 bl[474] br[474] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_475 bl[475] br[475] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_476 bl[476] br[476] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_477 bl[477] br[477] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_478 bl[478] br[478] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_479 bl[479] br[479] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_480 bl[480] br[480] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_481 bl[481] br[481] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_482 bl[482] br[482] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_483 bl[483] br[483] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_484 bl[484] br[484] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_485 bl[485] br[485] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_486 bl[486] br[486] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_487 bl[487] br[487] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_488 bl[488] br[488] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_489 bl[489] br[489] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_490 bl[490] br[490] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_491 bl[491] br[491] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_492 bl[492] br[492] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_493 bl[493] br[493] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_494 bl[494] br[494] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_495 bl[495] br[495] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_496 bl[496] br[496] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_497 bl[497] br[497] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_498 bl[498] br[498] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_499 bl[499] br[499] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_500 bl[500] br[500] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_501 bl[501] br[501] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_502 bl[502] br[502] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_503 bl[503] br[503] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_504 bl[504] br[504] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_505 bl[505] br[505] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_506 bl[506] br[506] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_507 bl[507] br[507] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_508 bl[508] br[508] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_509 bl[509] br[509] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_510 bl[510] br[510] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_54_511 bl[511] br[511] vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xcell_55_0 bl[0] br[0] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_1 bl[1] br[1] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_2 bl[2] br[2] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_3 bl[3] br[3] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_4 bl[4] br[4] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_5 bl[5] br[5] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_6 bl[6] br[6] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_7 bl[7] br[7] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_8 bl[8] br[8] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_9 bl[9] br[9] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_10 bl[10] br[10] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_11 bl[11] br[11] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_12 bl[12] br[12] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_13 bl[13] br[13] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_14 bl[14] br[14] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_15 bl[15] br[15] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_16 bl[16] br[16] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_17 bl[17] br[17] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_18 bl[18] br[18] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_19 bl[19] br[19] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_20 bl[20] br[20] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_21 bl[21] br[21] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_22 bl[22] br[22] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_23 bl[23] br[23] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_24 bl[24] br[24] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_25 bl[25] br[25] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_26 bl[26] br[26] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_27 bl[27] br[27] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_28 bl[28] br[28] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_29 bl[29] br[29] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_30 bl[30] br[30] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_31 bl[31] br[31] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_32 bl[32] br[32] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_33 bl[33] br[33] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_34 bl[34] br[34] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_35 bl[35] br[35] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_36 bl[36] br[36] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_37 bl[37] br[37] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_38 bl[38] br[38] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_39 bl[39] br[39] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_40 bl[40] br[40] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_41 bl[41] br[41] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_42 bl[42] br[42] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_43 bl[43] br[43] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_44 bl[44] br[44] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_45 bl[45] br[45] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_46 bl[46] br[46] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_47 bl[47] br[47] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_48 bl[48] br[48] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_49 bl[49] br[49] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_50 bl[50] br[50] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_51 bl[51] br[51] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_52 bl[52] br[52] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_53 bl[53] br[53] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_54 bl[54] br[54] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_55 bl[55] br[55] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_56 bl[56] br[56] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_57 bl[57] br[57] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_58 bl[58] br[58] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_59 bl[59] br[59] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_60 bl[60] br[60] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_61 bl[61] br[61] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_62 bl[62] br[62] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_63 bl[63] br[63] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_64 bl[64] br[64] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_65 bl[65] br[65] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_66 bl[66] br[66] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_67 bl[67] br[67] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_68 bl[68] br[68] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_69 bl[69] br[69] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_70 bl[70] br[70] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_71 bl[71] br[71] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_72 bl[72] br[72] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_73 bl[73] br[73] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_74 bl[74] br[74] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_75 bl[75] br[75] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_76 bl[76] br[76] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_77 bl[77] br[77] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_78 bl[78] br[78] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_79 bl[79] br[79] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_80 bl[80] br[80] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_81 bl[81] br[81] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_82 bl[82] br[82] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_83 bl[83] br[83] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_84 bl[84] br[84] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_85 bl[85] br[85] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_86 bl[86] br[86] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_87 bl[87] br[87] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_88 bl[88] br[88] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_89 bl[89] br[89] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_90 bl[90] br[90] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_91 bl[91] br[91] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_92 bl[92] br[92] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_93 bl[93] br[93] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_94 bl[94] br[94] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_95 bl[95] br[95] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_96 bl[96] br[96] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_97 bl[97] br[97] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_98 bl[98] br[98] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_99 bl[99] br[99] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_100 bl[100] br[100] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_101 bl[101] br[101] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_102 bl[102] br[102] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_103 bl[103] br[103] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_104 bl[104] br[104] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_105 bl[105] br[105] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_106 bl[106] br[106] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_107 bl[107] br[107] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_108 bl[108] br[108] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_109 bl[109] br[109] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_110 bl[110] br[110] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_111 bl[111] br[111] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_112 bl[112] br[112] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_113 bl[113] br[113] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_114 bl[114] br[114] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_115 bl[115] br[115] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_116 bl[116] br[116] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_117 bl[117] br[117] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_118 bl[118] br[118] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_119 bl[119] br[119] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_120 bl[120] br[120] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_121 bl[121] br[121] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_122 bl[122] br[122] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_123 bl[123] br[123] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_124 bl[124] br[124] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_125 bl[125] br[125] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_126 bl[126] br[126] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_127 bl[127] br[127] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_128 bl[128] br[128] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_129 bl[129] br[129] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_130 bl[130] br[130] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_131 bl[131] br[131] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_132 bl[132] br[132] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_133 bl[133] br[133] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_134 bl[134] br[134] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_135 bl[135] br[135] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_136 bl[136] br[136] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_137 bl[137] br[137] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_138 bl[138] br[138] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_139 bl[139] br[139] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_140 bl[140] br[140] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_141 bl[141] br[141] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_142 bl[142] br[142] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_143 bl[143] br[143] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_144 bl[144] br[144] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_145 bl[145] br[145] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_146 bl[146] br[146] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_147 bl[147] br[147] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_148 bl[148] br[148] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_149 bl[149] br[149] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_150 bl[150] br[150] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_151 bl[151] br[151] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_152 bl[152] br[152] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_153 bl[153] br[153] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_154 bl[154] br[154] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_155 bl[155] br[155] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_156 bl[156] br[156] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_157 bl[157] br[157] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_158 bl[158] br[158] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_159 bl[159] br[159] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_160 bl[160] br[160] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_161 bl[161] br[161] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_162 bl[162] br[162] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_163 bl[163] br[163] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_164 bl[164] br[164] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_165 bl[165] br[165] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_166 bl[166] br[166] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_167 bl[167] br[167] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_168 bl[168] br[168] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_169 bl[169] br[169] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_170 bl[170] br[170] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_171 bl[171] br[171] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_172 bl[172] br[172] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_173 bl[173] br[173] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_174 bl[174] br[174] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_175 bl[175] br[175] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_176 bl[176] br[176] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_177 bl[177] br[177] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_178 bl[178] br[178] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_179 bl[179] br[179] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_180 bl[180] br[180] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_181 bl[181] br[181] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_182 bl[182] br[182] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_183 bl[183] br[183] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_184 bl[184] br[184] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_185 bl[185] br[185] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_186 bl[186] br[186] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_187 bl[187] br[187] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_188 bl[188] br[188] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_189 bl[189] br[189] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_190 bl[190] br[190] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_191 bl[191] br[191] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_192 bl[192] br[192] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_193 bl[193] br[193] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_194 bl[194] br[194] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_195 bl[195] br[195] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_196 bl[196] br[196] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_197 bl[197] br[197] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_198 bl[198] br[198] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_199 bl[199] br[199] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_200 bl[200] br[200] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_201 bl[201] br[201] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_202 bl[202] br[202] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_203 bl[203] br[203] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_204 bl[204] br[204] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_205 bl[205] br[205] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_206 bl[206] br[206] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_207 bl[207] br[207] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_208 bl[208] br[208] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_209 bl[209] br[209] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_210 bl[210] br[210] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_211 bl[211] br[211] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_212 bl[212] br[212] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_213 bl[213] br[213] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_214 bl[214] br[214] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_215 bl[215] br[215] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_216 bl[216] br[216] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_217 bl[217] br[217] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_218 bl[218] br[218] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_219 bl[219] br[219] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_220 bl[220] br[220] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_221 bl[221] br[221] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_222 bl[222] br[222] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_223 bl[223] br[223] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_224 bl[224] br[224] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_225 bl[225] br[225] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_226 bl[226] br[226] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_227 bl[227] br[227] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_228 bl[228] br[228] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_229 bl[229] br[229] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_230 bl[230] br[230] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_231 bl[231] br[231] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_232 bl[232] br[232] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_233 bl[233] br[233] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_234 bl[234] br[234] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_235 bl[235] br[235] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_236 bl[236] br[236] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_237 bl[237] br[237] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_238 bl[238] br[238] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_239 bl[239] br[239] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_240 bl[240] br[240] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_241 bl[241] br[241] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_242 bl[242] br[242] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_243 bl[243] br[243] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_244 bl[244] br[244] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_245 bl[245] br[245] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_246 bl[246] br[246] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_247 bl[247] br[247] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_248 bl[248] br[248] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_249 bl[249] br[249] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_250 bl[250] br[250] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_251 bl[251] br[251] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_252 bl[252] br[252] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_253 bl[253] br[253] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_254 bl[254] br[254] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_255 bl[255] br[255] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_256 bl[256] br[256] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_257 bl[257] br[257] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_258 bl[258] br[258] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_259 bl[259] br[259] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_260 bl[260] br[260] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_261 bl[261] br[261] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_262 bl[262] br[262] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_263 bl[263] br[263] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_264 bl[264] br[264] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_265 bl[265] br[265] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_266 bl[266] br[266] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_267 bl[267] br[267] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_268 bl[268] br[268] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_269 bl[269] br[269] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_270 bl[270] br[270] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_271 bl[271] br[271] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_272 bl[272] br[272] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_273 bl[273] br[273] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_274 bl[274] br[274] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_275 bl[275] br[275] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_276 bl[276] br[276] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_277 bl[277] br[277] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_278 bl[278] br[278] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_279 bl[279] br[279] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_280 bl[280] br[280] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_281 bl[281] br[281] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_282 bl[282] br[282] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_283 bl[283] br[283] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_284 bl[284] br[284] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_285 bl[285] br[285] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_286 bl[286] br[286] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_287 bl[287] br[287] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_288 bl[288] br[288] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_289 bl[289] br[289] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_290 bl[290] br[290] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_291 bl[291] br[291] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_292 bl[292] br[292] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_293 bl[293] br[293] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_294 bl[294] br[294] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_295 bl[295] br[295] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_296 bl[296] br[296] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_297 bl[297] br[297] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_298 bl[298] br[298] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_299 bl[299] br[299] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_300 bl[300] br[300] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_301 bl[301] br[301] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_302 bl[302] br[302] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_303 bl[303] br[303] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_304 bl[304] br[304] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_305 bl[305] br[305] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_306 bl[306] br[306] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_307 bl[307] br[307] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_308 bl[308] br[308] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_309 bl[309] br[309] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_310 bl[310] br[310] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_311 bl[311] br[311] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_312 bl[312] br[312] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_313 bl[313] br[313] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_314 bl[314] br[314] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_315 bl[315] br[315] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_316 bl[316] br[316] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_317 bl[317] br[317] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_318 bl[318] br[318] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_319 bl[319] br[319] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_320 bl[320] br[320] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_321 bl[321] br[321] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_322 bl[322] br[322] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_323 bl[323] br[323] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_324 bl[324] br[324] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_325 bl[325] br[325] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_326 bl[326] br[326] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_327 bl[327] br[327] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_328 bl[328] br[328] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_329 bl[329] br[329] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_330 bl[330] br[330] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_331 bl[331] br[331] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_332 bl[332] br[332] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_333 bl[333] br[333] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_334 bl[334] br[334] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_335 bl[335] br[335] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_336 bl[336] br[336] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_337 bl[337] br[337] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_338 bl[338] br[338] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_339 bl[339] br[339] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_340 bl[340] br[340] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_341 bl[341] br[341] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_342 bl[342] br[342] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_343 bl[343] br[343] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_344 bl[344] br[344] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_345 bl[345] br[345] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_346 bl[346] br[346] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_347 bl[347] br[347] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_348 bl[348] br[348] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_349 bl[349] br[349] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_350 bl[350] br[350] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_351 bl[351] br[351] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_352 bl[352] br[352] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_353 bl[353] br[353] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_354 bl[354] br[354] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_355 bl[355] br[355] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_356 bl[356] br[356] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_357 bl[357] br[357] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_358 bl[358] br[358] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_359 bl[359] br[359] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_360 bl[360] br[360] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_361 bl[361] br[361] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_362 bl[362] br[362] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_363 bl[363] br[363] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_364 bl[364] br[364] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_365 bl[365] br[365] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_366 bl[366] br[366] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_367 bl[367] br[367] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_368 bl[368] br[368] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_369 bl[369] br[369] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_370 bl[370] br[370] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_371 bl[371] br[371] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_372 bl[372] br[372] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_373 bl[373] br[373] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_374 bl[374] br[374] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_375 bl[375] br[375] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_376 bl[376] br[376] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_377 bl[377] br[377] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_378 bl[378] br[378] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_379 bl[379] br[379] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_380 bl[380] br[380] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_381 bl[381] br[381] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_382 bl[382] br[382] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_383 bl[383] br[383] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_384 bl[384] br[384] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_385 bl[385] br[385] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_386 bl[386] br[386] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_387 bl[387] br[387] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_388 bl[388] br[388] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_389 bl[389] br[389] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_390 bl[390] br[390] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_391 bl[391] br[391] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_392 bl[392] br[392] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_393 bl[393] br[393] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_394 bl[394] br[394] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_395 bl[395] br[395] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_396 bl[396] br[396] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_397 bl[397] br[397] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_398 bl[398] br[398] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_399 bl[399] br[399] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_400 bl[400] br[400] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_401 bl[401] br[401] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_402 bl[402] br[402] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_403 bl[403] br[403] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_404 bl[404] br[404] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_405 bl[405] br[405] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_406 bl[406] br[406] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_407 bl[407] br[407] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_408 bl[408] br[408] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_409 bl[409] br[409] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_410 bl[410] br[410] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_411 bl[411] br[411] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_412 bl[412] br[412] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_413 bl[413] br[413] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_414 bl[414] br[414] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_415 bl[415] br[415] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_416 bl[416] br[416] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_417 bl[417] br[417] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_418 bl[418] br[418] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_419 bl[419] br[419] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_420 bl[420] br[420] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_421 bl[421] br[421] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_422 bl[422] br[422] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_423 bl[423] br[423] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_424 bl[424] br[424] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_425 bl[425] br[425] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_426 bl[426] br[426] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_427 bl[427] br[427] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_428 bl[428] br[428] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_429 bl[429] br[429] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_430 bl[430] br[430] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_431 bl[431] br[431] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_432 bl[432] br[432] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_433 bl[433] br[433] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_434 bl[434] br[434] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_435 bl[435] br[435] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_436 bl[436] br[436] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_437 bl[437] br[437] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_438 bl[438] br[438] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_439 bl[439] br[439] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_440 bl[440] br[440] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_441 bl[441] br[441] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_442 bl[442] br[442] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_443 bl[443] br[443] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_444 bl[444] br[444] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_445 bl[445] br[445] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_446 bl[446] br[446] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_447 bl[447] br[447] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_448 bl[448] br[448] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_449 bl[449] br[449] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_450 bl[450] br[450] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_451 bl[451] br[451] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_452 bl[452] br[452] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_453 bl[453] br[453] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_454 bl[454] br[454] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_455 bl[455] br[455] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_456 bl[456] br[456] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_457 bl[457] br[457] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_458 bl[458] br[458] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_459 bl[459] br[459] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_460 bl[460] br[460] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_461 bl[461] br[461] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_462 bl[462] br[462] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_463 bl[463] br[463] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_464 bl[464] br[464] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_465 bl[465] br[465] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_466 bl[466] br[466] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_467 bl[467] br[467] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_468 bl[468] br[468] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_469 bl[469] br[469] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_470 bl[470] br[470] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_471 bl[471] br[471] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_472 bl[472] br[472] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_473 bl[473] br[473] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_474 bl[474] br[474] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_475 bl[475] br[475] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_476 bl[476] br[476] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_477 bl[477] br[477] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_478 bl[478] br[478] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_479 bl[479] br[479] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_480 bl[480] br[480] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_481 bl[481] br[481] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_482 bl[482] br[482] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_483 bl[483] br[483] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_484 bl[484] br[484] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_485 bl[485] br[485] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_486 bl[486] br[486] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_487 bl[487] br[487] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_488 bl[488] br[488] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_489 bl[489] br[489] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_490 bl[490] br[490] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_491 bl[491] br[491] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_492 bl[492] br[492] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_493 bl[493] br[493] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_494 bl[494] br[494] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_495 bl[495] br[495] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_496 bl[496] br[496] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_497 bl[497] br[497] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_498 bl[498] br[498] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_499 bl[499] br[499] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_500 bl[500] br[500] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_501 bl[501] br[501] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_502 bl[502] br[502] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_503 bl[503] br[503] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_504 bl[504] br[504] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_505 bl[505] br[505] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_506 bl[506] br[506] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_507 bl[507] br[507] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_508 bl[508] br[508] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_509 bl[509] br[509] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_510 bl[510] br[510] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_55_511 bl[511] br[511] vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xcell_56_0 bl[0] br[0] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_1 bl[1] br[1] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_2 bl[2] br[2] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_3 bl[3] br[3] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_4 bl[4] br[4] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_5 bl[5] br[5] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_6 bl[6] br[6] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_7 bl[7] br[7] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_8 bl[8] br[8] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_9 bl[9] br[9] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_10 bl[10] br[10] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_11 bl[11] br[11] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_12 bl[12] br[12] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_13 bl[13] br[13] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_14 bl[14] br[14] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_15 bl[15] br[15] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_16 bl[16] br[16] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_17 bl[17] br[17] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_18 bl[18] br[18] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_19 bl[19] br[19] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_20 bl[20] br[20] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_21 bl[21] br[21] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_22 bl[22] br[22] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_23 bl[23] br[23] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_24 bl[24] br[24] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_25 bl[25] br[25] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_26 bl[26] br[26] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_27 bl[27] br[27] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_28 bl[28] br[28] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_29 bl[29] br[29] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_30 bl[30] br[30] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_31 bl[31] br[31] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_32 bl[32] br[32] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_33 bl[33] br[33] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_34 bl[34] br[34] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_35 bl[35] br[35] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_36 bl[36] br[36] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_37 bl[37] br[37] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_38 bl[38] br[38] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_39 bl[39] br[39] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_40 bl[40] br[40] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_41 bl[41] br[41] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_42 bl[42] br[42] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_43 bl[43] br[43] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_44 bl[44] br[44] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_45 bl[45] br[45] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_46 bl[46] br[46] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_47 bl[47] br[47] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_48 bl[48] br[48] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_49 bl[49] br[49] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_50 bl[50] br[50] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_51 bl[51] br[51] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_52 bl[52] br[52] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_53 bl[53] br[53] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_54 bl[54] br[54] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_55 bl[55] br[55] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_56 bl[56] br[56] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_57 bl[57] br[57] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_58 bl[58] br[58] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_59 bl[59] br[59] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_60 bl[60] br[60] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_61 bl[61] br[61] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_62 bl[62] br[62] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_63 bl[63] br[63] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_64 bl[64] br[64] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_65 bl[65] br[65] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_66 bl[66] br[66] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_67 bl[67] br[67] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_68 bl[68] br[68] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_69 bl[69] br[69] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_70 bl[70] br[70] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_71 bl[71] br[71] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_72 bl[72] br[72] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_73 bl[73] br[73] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_74 bl[74] br[74] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_75 bl[75] br[75] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_76 bl[76] br[76] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_77 bl[77] br[77] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_78 bl[78] br[78] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_79 bl[79] br[79] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_80 bl[80] br[80] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_81 bl[81] br[81] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_82 bl[82] br[82] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_83 bl[83] br[83] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_84 bl[84] br[84] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_85 bl[85] br[85] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_86 bl[86] br[86] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_87 bl[87] br[87] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_88 bl[88] br[88] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_89 bl[89] br[89] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_90 bl[90] br[90] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_91 bl[91] br[91] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_92 bl[92] br[92] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_93 bl[93] br[93] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_94 bl[94] br[94] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_95 bl[95] br[95] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_96 bl[96] br[96] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_97 bl[97] br[97] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_98 bl[98] br[98] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_99 bl[99] br[99] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_100 bl[100] br[100] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_101 bl[101] br[101] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_102 bl[102] br[102] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_103 bl[103] br[103] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_104 bl[104] br[104] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_105 bl[105] br[105] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_106 bl[106] br[106] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_107 bl[107] br[107] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_108 bl[108] br[108] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_109 bl[109] br[109] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_110 bl[110] br[110] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_111 bl[111] br[111] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_112 bl[112] br[112] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_113 bl[113] br[113] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_114 bl[114] br[114] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_115 bl[115] br[115] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_116 bl[116] br[116] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_117 bl[117] br[117] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_118 bl[118] br[118] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_119 bl[119] br[119] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_120 bl[120] br[120] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_121 bl[121] br[121] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_122 bl[122] br[122] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_123 bl[123] br[123] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_124 bl[124] br[124] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_125 bl[125] br[125] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_126 bl[126] br[126] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_127 bl[127] br[127] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_128 bl[128] br[128] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_129 bl[129] br[129] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_130 bl[130] br[130] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_131 bl[131] br[131] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_132 bl[132] br[132] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_133 bl[133] br[133] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_134 bl[134] br[134] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_135 bl[135] br[135] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_136 bl[136] br[136] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_137 bl[137] br[137] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_138 bl[138] br[138] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_139 bl[139] br[139] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_140 bl[140] br[140] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_141 bl[141] br[141] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_142 bl[142] br[142] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_143 bl[143] br[143] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_144 bl[144] br[144] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_145 bl[145] br[145] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_146 bl[146] br[146] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_147 bl[147] br[147] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_148 bl[148] br[148] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_149 bl[149] br[149] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_150 bl[150] br[150] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_151 bl[151] br[151] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_152 bl[152] br[152] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_153 bl[153] br[153] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_154 bl[154] br[154] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_155 bl[155] br[155] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_156 bl[156] br[156] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_157 bl[157] br[157] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_158 bl[158] br[158] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_159 bl[159] br[159] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_160 bl[160] br[160] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_161 bl[161] br[161] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_162 bl[162] br[162] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_163 bl[163] br[163] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_164 bl[164] br[164] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_165 bl[165] br[165] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_166 bl[166] br[166] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_167 bl[167] br[167] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_168 bl[168] br[168] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_169 bl[169] br[169] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_170 bl[170] br[170] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_171 bl[171] br[171] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_172 bl[172] br[172] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_173 bl[173] br[173] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_174 bl[174] br[174] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_175 bl[175] br[175] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_176 bl[176] br[176] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_177 bl[177] br[177] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_178 bl[178] br[178] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_179 bl[179] br[179] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_180 bl[180] br[180] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_181 bl[181] br[181] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_182 bl[182] br[182] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_183 bl[183] br[183] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_184 bl[184] br[184] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_185 bl[185] br[185] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_186 bl[186] br[186] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_187 bl[187] br[187] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_188 bl[188] br[188] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_189 bl[189] br[189] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_190 bl[190] br[190] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_191 bl[191] br[191] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_192 bl[192] br[192] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_193 bl[193] br[193] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_194 bl[194] br[194] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_195 bl[195] br[195] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_196 bl[196] br[196] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_197 bl[197] br[197] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_198 bl[198] br[198] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_199 bl[199] br[199] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_200 bl[200] br[200] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_201 bl[201] br[201] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_202 bl[202] br[202] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_203 bl[203] br[203] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_204 bl[204] br[204] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_205 bl[205] br[205] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_206 bl[206] br[206] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_207 bl[207] br[207] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_208 bl[208] br[208] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_209 bl[209] br[209] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_210 bl[210] br[210] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_211 bl[211] br[211] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_212 bl[212] br[212] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_213 bl[213] br[213] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_214 bl[214] br[214] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_215 bl[215] br[215] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_216 bl[216] br[216] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_217 bl[217] br[217] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_218 bl[218] br[218] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_219 bl[219] br[219] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_220 bl[220] br[220] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_221 bl[221] br[221] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_222 bl[222] br[222] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_223 bl[223] br[223] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_224 bl[224] br[224] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_225 bl[225] br[225] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_226 bl[226] br[226] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_227 bl[227] br[227] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_228 bl[228] br[228] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_229 bl[229] br[229] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_230 bl[230] br[230] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_231 bl[231] br[231] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_232 bl[232] br[232] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_233 bl[233] br[233] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_234 bl[234] br[234] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_235 bl[235] br[235] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_236 bl[236] br[236] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_237 bl[237] br[237] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_238 bl[238] br[238] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_239 bl[239] br[239] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_240 bl[240] br[240] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_241 bl[241] br[241] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_242 bl[242] br[242] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_243 bl[243] br[243] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_244 bl[244] br[244] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_245 bl[245] br[245] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_246 bl[246] br[246] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_247 bl[247] br[247] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_248 bl[248] br[248] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_249 bl[249] br[249] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_250 bl[250] br[250] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_251 bl[251] br[251] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_252 bl[252] br[252] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_253 bl[253] br[253] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_254 bl[254] br[254] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_255 bl[255] br[255] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_256 bl[256] br[256] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_257 bl[257] br[257] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_258 bl[258] br[258] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_259 bl[259] br[259] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_260 bl[260] br[260] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_261 bl[261] br[261] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_262 bl[262] br[262] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_263 bl[263] br[263] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_264 bl[264] br[264] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_265 bl[265] br[265] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_266 bl[266] br[266] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_267 bl[267] br[267] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_268 bl[268] br[268] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_269 bl[269] br[269] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_270 bl[270] br[270] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_271 bl[271] br[271] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_272 bl[272] br[272] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_273 bl[273] br[273] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_274 bl[274] br[274] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_275 bl[275] br[275] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_276 bl[276] br[276] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_277 bl[277] br[277] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_278 bl[278] br[278] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_279 bl[279] br[279] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_280 bl[280] br[280] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_281 bl[281] br[281] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_282 bl[282] br[282] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_283 bl[283] br[283] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_284 bl[284] br[284] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_285 bl[285] br[285] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_286 bl[286] br[286] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_287 bl[287] br[287] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_288 bl[288] br[288] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_289 bl[289] br[289] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_290 bl[290] br[290] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_291 bl[291] br[291] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_292 bl[292] br[292] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_293 bl[293] br[293] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_294 bl[294] br[294] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_295 bl[295] br[295] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_296 bl[296] br[296] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_297 bl[297] br[297] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_298 bl[298] br[298] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_299 bl[299] br[299] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_300 bl[300] br[300] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_301 bl[301] br[301] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_302 bl[302] br[302] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_303 bl[303] br[303] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_304 bl[304] br[304] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_305 bl[305] br[305] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_306 bl[306] br[306] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_307 bl[307] br[307] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_308 bl[308] br[308] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_309 bl[309] br[309] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_310 bl[310] br[310] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_311 bl[311] br[311] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_312 bl[312] br[312] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_313 bl[313] br[313] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_314 bl[314] br[314] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_315 bl[315] br[315] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_316 bl[316] br[316] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_317 bl[317] br[317] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_318 bl[318] br[318] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_319 bl[319] br[319] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_320 bl[320] br[320] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_321 bl[321] br[321] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_322 bl[322] br[322] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_323 bl[323] br[323] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_324 bl[324] br[324] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_325 bl[325] br[325] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_326 bl[326] br[326] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_327 bl[327] br[327] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_328 bl[328] br[328] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_329 bl[329] br[329] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_330 bl[330] br[330] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_331 bl[331] br[331] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_332 bl[332] br[332] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_333 bl[333] br[333] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_334 bl[334] br[334] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_335 bl[335] br[335] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_336 bl[336] br[336] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_337 bl[337] br[337] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_338 bl[338] br[338] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_339 bl[339] br[339] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_340 bl[340] br[340] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_341 bl[341] br[341] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_342 bl[342] br[342] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_343 bl[343] br[343] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_344 bl[344] br[344] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_345 bl[345] br[345] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_346 bl[346] br[346] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_347 bl[347] br[347] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_348 bl[348] br[348] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_349 bl[349] br[349] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_350 bl[350] br[350] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_351 bl[351] br[351] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_352 bl[352] br[352] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_353 bl[353] br[353] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_354 bl[354] br[354] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_355 bl[355] br[355] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_356 bl[356] br[356] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_357 bl[357] br[357] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_358 bl[358] br[358] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_359 bl[359] br[359] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_360 bl[360] br[360] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_361 bl[361] br[361] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_362 bl[362] br[362] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_363 bl[363] br[363] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_364 bl[364] br[364] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_365 bl[365] br[365] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_366 bl[366] br[366] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_367 bl[367] br[367] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_368 bl[368] br[368] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_369 bl[369] br[369] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_370 bl[370] br[370] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_371 bl[371] br[371] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_372 bl[372] br[372] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_373 bl[373] br[373] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_374 bl[374] br[374] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_375 bl[375] br[375] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_376 bl[376] br[376] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_377 bl[377] br[377] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_378 bl[378] br[378] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_379 bl[379] br[379] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_380 bl[380] br[380] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_381 bl[381] br[381] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_382 bl[382] br[382] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_383 bl[383] br[383] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_384 bl[384] br[384] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_385 bl[385] br[385] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_386 bl[386] br[386] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_387 bl[387] br[387] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_388 bl[388] br[388] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_389 bl[389] br[389] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_390 bl[390] br[390] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_391 bl[391] br[391] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_392 bl[392] br[392] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_393 bl[393] br[393] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_394 bl[394] br[394] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_395 bl[395] br[395] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_396 bl[396] br[396] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_397 bl[397] br[397] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_398 bl[398] br[398] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_399 bl[399] br[399] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_400 bl[400] br[400] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_401 bl[401] br[401] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_402 bl[402] br[402] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_403 bl[403] br[403] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_404 bl[404] br[404] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_405 bl[405] br[405] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_406 bl[406] br[406] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_407 bl[407] br[407] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_408 bl[408] br[408] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_409 bl[409] br[409] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_410 bl[410] br[410] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_411 bl[411] br[411] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_412 bl[412] br[412] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_413 bl[413] br[413] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_414 bl[414] br[414] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_415 bl[415] br[415] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_416 bl[416] br[416] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_417 bl[417] br[417] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_418 bl[418] br[418] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_419 bl[419] br[419] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_420 bl[420] br[420] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_421 bl[421] br[421] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_422 bl[422] br[422] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_423 bl[423] br[423] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_424 bl[424] br[424] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_425 bl[425] br[425] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_426 bl[426] br[426] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_427 bl[427] br[427] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_428 bl[428] br[428] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_429 bl[429] br[429] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_430 bl[430] br[430] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_431 bl[431] br[431] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_432 bl[432] br[432] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_433 bl[433] br[433] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_434 bl[434] br[434] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_435 bl[435] br[435] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_436 bl[436] br[436] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_437 bl[437] br[437] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_438 bl[438] br[438] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_439 bl[439] br[439] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_440 bl[440] br[440] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_441 bl[441] br[441] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_442 bl[442] br[442] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_443 bl[443] br[443] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_444 bl[444] br[444] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_445 bl[445] br[445] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_446 bl[446] br[446] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_447 bl[447] br[447] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_448 bl[448] br[448] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_449 bl[449] br[449] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_450 bl[450] br[450] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_451 bl[451] br[451] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_452 bl[452] br[452] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_453 bl[453] br[453] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_454 bl[454] br[454] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_455 bl[455] br[455] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_456 bl[456] br[456] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_457 bl[457] br[457] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_458 bl[458] br[458] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_459 bl[459] br[459] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_460 bl[460] br[460] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_461 bl[461] br[461] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_462 bl[462] br[462] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_463 bl[463] br[463] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_464 bl[464] br[464] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_465 bl[465] br[465] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_466 bl[466] br[466] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_467 bl[467] br[467] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_468 bl[468] br[468] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_469 bl[469] br[469] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_470 bl[470] br[470] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_471 bl[471] br[471] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_472 bl[472] br[472] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_473 bl[473] br[473] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_474 bl[474] br[474] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_475 bl[475] br[475] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_476 bl[476] br[476] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_477 bl[477] br[477] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_478 bl[478] br[478] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_479 bl[479] br[479] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_480 bl[480] br[480] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_481 bl[481] br[481] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_482 bl[482] br[482] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_483 bl[483] br[483] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_484 bl[484] br[484] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_485 bl[485] br[485] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_486 bl[486] br[486] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_487 bl[487] br[487] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_488 bl[488] br[488] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_489 bl[489] br[489] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_490 bl[490] br[490] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_491 bl[491] br[491] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_492 bl[492] br[492] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_493 bl[493] br[493] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_494 bl[494] br[494] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_495 bl[495] br[495] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_496 bl[496] br[496] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_497 bl[497] br[497] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_498 bl[498] br[498] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_499 bl[499] br[499] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_500 bl[500] br[500] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_501 bl[501] br[501] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_502 bl[502] br[502] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_503 bl[503] br[503] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_504 bl[504] br[504] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_505 bl[505] br[505] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_506 bl[506] br[506] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_507 bl[507] br[507] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_508 bl[508] br[508] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_509 bl[509] br[509] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_510 bl[510] br[510] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_56_511 bl[511] br[511] vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xcell_57_0 bl[0] br[0] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_1 bl[1] br[1] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_2 bl[2] br[2] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_3 bl[3] br[3] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_4 bl[4] br[4] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_5 bl[5] br[5] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_6 bl[6] br[6] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_7 bl[7] br[7] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_8 bl[8] br[8] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_9 bl[9] br[9] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_10 bl[10] br[10] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_11 bl[11] br[11] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_12 bl[12] br[12] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_13 bl[13] br[13] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_14 bl[14] br[14] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_15 bl[15] br[15] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_16 bl[16] br[16] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_17 bl[17] br[17] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_18 bl[18] br[18] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_19 bl[19] br[19] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_20 bl[20] br[20] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_21 bl[21] br[21] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_22 bl[22] br[22] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_23 bl[23] br[23] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_24 bl[24] br[24] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_25 bl[25] br[25] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_26 bl[26] br[26] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_27 bl[27] br[27] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_28 bl[28] br[28] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_29 bl[29] br[29] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_30 bl[30] br[30] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_31 bl[31] br[31] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_32 bl[32] br[32] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_33 bl[33] br[33] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_34 bl[34] br[34] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_35 bl[35] br[35] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_36 bl[36] br[36] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_37 bl[37] br[37] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_38 bl[38] br[38] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_39 bl[39] br[39] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_40 bl[40] br[40] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_41 bl[41] br[41] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_42 bl[42] br[42] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_43 bl[43] br[43] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_44 bl[44] br[44] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_45 bl[45] br[45] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_46 bl[46] br[46] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_47 bl[47] br[47] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_48 bl[48] br[48] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_49 bl[49] br[49] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_50 bl[50] br[50] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_51 bl[51] br[51] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_52 bl[52] br[52] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_53 bl[53] br[53] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_54 bl[54] br[54] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_55 bl[55] br[55] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_56 bl[56] br[56] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_57 bl[57] br[57] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_58 bl[58] br[58] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_59 bl[59] br[59] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_60 bl[60] br[60] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_61 bl[61] br[61] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_62 bl[62] br[62] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_63 bl[63] br[63] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_64 bl[64] br[64] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_65 bl[65] br[65] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_66 bl[66] br[66] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_67 bl[67] br[67] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_68 bl[68] br[68] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_69 bl[69] br[69] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_70 bl[70] br[70] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_71 bl[71] br[71] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_72 bl[72] br[72] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_73 bl[73] br[73] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_74 bl[74] br[74] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_75 bl[75] br[75] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_76 bl[76] br[76] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_77 bl[77] br[77] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_78 bl[78] br[78] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_79 bl[79] br[79] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_80 bl[80] br[80] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_81 bl[81] br[81] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_82 bl[82] br[82] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_83 bl[83] br[83] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_84 bl[84] br[84] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_85 bl[85] br[85] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_86 bl[86] br[86] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_87 bl[87] br[87] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_88 bl[88] br[88] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_89 bl[89] br[89] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_90 bl[90] br[90] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_91 bl[91] br[91] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_92 bl[92] br[92] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_93 bl[93] br[93] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_94 bl[94] br[94] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_95 bl[95] br[95] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_96 bl[96] br[96] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_97 bl[97] br[97] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_98 bl[98] br[98] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_99 bl[99] br[99] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_100 bl[100] br[100] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_101 bl[101] br[101] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_102 bl[102] br[102] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_103 bl[103] br[103] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_104 bl[104] br[104] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_105 bl[105] br[105] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_106 bl[106] br[106] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_107 bl[107] br[107] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_108 bl[108] br[108] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_109 bl[109] br[109] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_110 bl[110] br[110] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_111 bl[111] br[111] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_112 bl[112] br[112] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_113 bl[113] br[113] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_114 bl[114] br[114] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_115 bl[115] br[115] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_116 bl[116] br[116] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_117 bl[117] br[117] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_118 bl[118] br[118] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_119 bl[119] br[119] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_120 bl[120] br[120] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_121 bl[121] br[121] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_122 bl[122] br[122] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_123 bl[123] br[123] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_124 bl[124] br[124] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_125 bl[125] br[125] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_126 bl[126] br[126] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_127 bl[127] br[127] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_128 bl[128] br[128] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_129 bl[129] br[129] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_130 bl[130] br[130] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_131 bl[131] br[131] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_132 bl[132] br[132] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_133 bl[133] br[133] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_134 bl[134] br[134] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_135 bl[135] br[135] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_136 bl[136] br[136] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_137 bl[137] br[137] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_138 bl[138] br[138] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_139 bl[139] br[139] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_140 bl[140] br[140] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_141 bl[141] br[141] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_142 bl[142] br[142] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_143 bl[143] br[143] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_144 bl[144] br[144] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_145 bl[145] br[145] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_146 bl[146] br[146] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_147 bl[147] br[147] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_148 bl[148] br[148] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_149 bl[149] br[149] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_150 bl[150] br[150] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_151 bl[151] br[151] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_152 bl[152] br[152] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_153 bl[153] br[153] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_154 bl[154] br[154] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_155 bl[155] br[155] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_156 bl[156] br[156] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_157 bl[157] br[157] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_158 bl[158] br[158] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_159 bl[159] br[159] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_160 bl[160] br[160] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_161 bl[161] br[161] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_162 bl[162] br[162] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_163 bl[163] br[163] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_164 bl[164] br[164] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_165 bl[165] br[165] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_166 bl[166] br[166] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_167 bl[167] br[167] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_168 bl[168] br[168] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_169 bl[169] br[169] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_170 bl[170] br[170] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_171 bl[171] br[171] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_172 bl[172] br[172] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_173 bl[173] br[173] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_174 bl[174] br[174] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_175 bl[175] br[175] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_176 bl[176] br[176] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_177 bl[177] br[177] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_178 bl[178] br[178] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_179 bl[179] br[179] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_180 bl[180] br[180] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_181 bl[181] br[181] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_182 bl[182] br[182] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_183 bl[183] br[183] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_184 bl[184] br[184] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_185 bl[185] br[185] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_186 bl[186] br[186] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_187 bl[187] br[187] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_188 bl[188] br[188] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_189 bl[189] br[189] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_190 bl[190] br[190] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_191 bl[191] br[191] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_192 bl[192] br[192] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_193 bl[193] br[193] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_194 bl[194] br[194] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_195 bl[195] br[195] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_196 bl[196] br[196] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_197 bl[197] br[197] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_198 bl[198] br[198] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_199 bl[199] br[199] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_200 bl[200] br[200] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_201 bl[201] br[201] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_202 bl[202] br[202] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_203 bl[203] br[203] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_204 bl[204] br[204] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_205 bl[205] br[205] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_206 bl[206] br[206] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_207 bl[207] br[207] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_208 bl[208] br[208] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_209 bl[209] br[209] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_210 bl[210] br[210] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_211 bl[211] br[211] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_212 bl[212] br[212] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_213 bl[213] br[213] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_214 bl[214] br[214] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_215 bl[215] br[215] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_216 bl[216] br[216] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_217 bl[217] br[217] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_218 bl[218] br[218] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_219 bl[219] br[219] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_220 bl[220] br[220] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_221 bl[221] br[221] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_222 bl[222] br[222] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_223 bl[223] br[223] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_224 bl[224] br[224] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_225 bl[225] br[225] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_226 bl[226] br[226] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_227 bl[227] br[227] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_228 bl[228] br[228] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_229 bl[229] br[229] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_230 bl[230] br[230] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_231 bl[231] br[231] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_232 bl[232] br[232] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_233 bl[233] br[233] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_234 bl[234] br[234] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_235 bl[235] br[235] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_236 bl[236] br[236] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_237 bl[237] br[237] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_238 bl[238] br[238] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_239 bl[239] br[239] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_240 bl[240] br[240] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_241 bl[241] br[241] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_242 bl[242] br[242] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_243 bl[243] br[243] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_244 bl[244] br[244] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_245 bl[245] br[245] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_246 bl[246] br[246] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_247 bl[247] br[247] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_248 bl[248] br[248] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_249 bl[249] br[249] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_250 bl[250] br[250] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_251 bl[251] br[251] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_252 bl[252] br[252] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_253 bl[253] br[253] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_254 bl[254] br[254] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_255 bl[255] br[255] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_256 bl[256] br[256] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_257 bl[257] br[257] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_258 bl[258] br[258] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_259 bl[259] br[259] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_260 bl[260] br[260] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_261 bl[261] br[261] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_262 bl[262] br[262] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_263 bl[263] br[263] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_264 bl[264] br[264] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_265 bl[265] br[265] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_266 bl[266] br[266] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_267 bl[267] br[267] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_268 bl[268] br[268] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_269 bl[269] br[269] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_270 bl[270] br[270] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_271 bl[271] br[271] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_272 bl[272] br[272] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_273 bl[273] br[273] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_274 bl[274] br[274] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_275 bl[275] br[275] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_276 bl[276] br[276] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_277 bl[277] br[277] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_278 bl[278] br[278] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_279 bl[279] br[279] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_280 bl[280] br[280] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_281 bl[281] br[281] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_282 bl[282] br[282] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_283 bl[283] br[283] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_284 bl[284] br[284] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_285 bl[285] br[285] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_286 bl[286] br[286] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_287 bl[287] br[287] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_288 bl[288] br[288] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_289 bl[289] br[289] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_290 bl[290] br[290] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_291 bl[291] br[291] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_292 bl[292] br[292] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_293 bl[293] br[293] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_294 bl[294] br[294] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_295 bl[295] br[295] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_296 bl[296] br[296] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_297 bl[297] br[297] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_298 bl[298] br[298] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_299 bl[299] br[299] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_300 bl[300] br[300] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_301 bl[301] br[301] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_302 bl[302] br[302] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_303 bl[303] br[303] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_304 bl[304] br[304] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_305 bl[305] br[305] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_306 bl[306] br[306] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_307 bl[307] br[307] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_308 bl[308] br[308] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_309 bl[309] br[309] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_310 bl[310] br[310] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_311 bl[311] br[311] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_312 bl[312] br[312] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_313 bl[313] br[313] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_314 bl[314] br[314] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_315 bl[315] br[315] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_316 bl[316] br[316] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_317 bl[317] br[317] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_318 bl[318] br[318] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_319 bl[319] br[319] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_320 bl[320] br[320] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_321 bl[321] br[321] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_322 bl[322] br[322] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_323 bl[323] br[323] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_324 bl[324] br[324] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_325 bl[325] br[325] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_326 bl[326] br[326] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_327 bl[327] br[327] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_328 bl[328] br[328] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_329 bl[329] br[329] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_330 bl[330] br[330] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_331 bl[331] br[331] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_332 bl[332] br[332] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_333 bl[333] br[333] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_334 bl[334] br[334] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_335 bl[335] br[335] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_336 bl[336] br[336] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_337 bl[337] br[337] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_338 bl[338] br[338] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_339 bl[339] br[339] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_340 bl[340] br[340] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_341 bl[341] br[341] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_342 bl[342] br[342] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_343 bl[343] br[343] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_344 bl[344] br[344] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_345 bl[345] br[345] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_346 bl[346] br[346] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_347 bl[347] br[347] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_348 bl[348] br[348] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_349 bl[349] br[349] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_350 bl[350] br[350] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_351 bl[351] br[351] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_352 bl[352] br[352] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_353 bl[353] br[353] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_354 bl[354] br[354] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_355 bl[355] br[355] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_356 bl[356] br[356] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_357 bl[357] br[357] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_358 bl[358] br[358] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_359 bl[359] br[359] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_360 bl[360] br[360] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_361 bl[361] br[361] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_362 bl[362] br[362] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_363 bl[363] br[363] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_364 bl[364] br[364] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_365 bl[365] br[365] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_366 bl[366] br[366] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_367 bl[367] br[367] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_368 bl[368] br[368] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_369 bl[369] br[369] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_370 bl[370] br[370] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_371 bl[371] br[371] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_372 bl[372] br[372] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_373 bl[373] br[373] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_374 bl[374] br[374] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_375 bl[375] br[375] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_376 bl[376] br[376] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_377 bl[377] br[377] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_378 bl[378] br[378] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_379 bl[379] br[379] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_380 bl[380] br[380] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_381 bl[381] br[381] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_382 bl[382] br[382] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_383 bl[383] br[383] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_384 bl[384] br[384] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_385 bl[385] br[385] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_386 bl[386] br[386] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_387 bl[387] br[387] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_388 bl[388] br[388] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_389 bl[389] br[389] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_390 bl[390] br[390] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_391 bl[391] br[391] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_392 bl[392] br[392] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_393 bl[393] br[393] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_394 bl[394] br[394] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_395 bl[395] br[395] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_396 bl[396] br[396] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_397 bl[397] br[397] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_398 bl[398] br[398] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_399 bl[399] br[399] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_400 bl[400] br[400] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_401 bl[401] br[401] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_402 bl[402] br[402] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_403 bl[403] br[403] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_404 bl[404] br[404] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_405 bl[405] br[405] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_406 bl[406] br[406] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_407 bl[407] br[407] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_408 bl[408] br[408] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_409 bl[409] br[409] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_410 bl[410] br[410] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_411 bl[411] br[411] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_412 bl[412] br[412] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_413 bl[413] br[413] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_414 bl[414] br[414] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_415 bl[415] br[415] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_416 bl[416] br[416] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_417 bl[417] br[417] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_418 bl[418] br[418] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_419 bl[419] br[419] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_420 bl[420] br[420] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_421 bl[421] br[421] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_422 bl[422] br[422] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_423 bl[423] br[423] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_424 bl[424] br[424] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_425 bl[425] br[425] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_426 bl[426] br[426] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_427 bl[427] br[427] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_428 bl[428] br[428] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_429 bl[429] br[429] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_430 bl[430] br[430] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_431 bl[431] br[431] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_432 bl[432] br[432] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_433 bl[433] br[433] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_434 bl[434] br[434] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_435 bl[435] br[435] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_436 bl[436] br[436] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_437 bl[437] br[437] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_438 bl[438] br[438] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_439 bl[439] br[439] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_440 bl[440] br[440] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_441 bl[441] br[441] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_442 bl[442] br[442] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_443 bl[443] br[443] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_444 bl[444] br[444] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_445 bl[445] br[445] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_446 bl[446] br[446] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_447 bl[447] br[447] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_448 bl[448] br[448] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_449 bl[449] br[449] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_450 bl[450] br[450] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_451 bl[451] br[451] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_452 bl[452] br[452] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_453 bl[453] br[453] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_454 bl[454] br[454] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_455 bl[455] br[455] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_456 bl[456] br[456] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_457 bl[457] br[457] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_458 bl[458] br[458] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_459 bl[459] br[459] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_460 bl[460] br[460] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_461 bl[461] br[461] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_462 bl[462] br[462] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_463 bl[463] br[463] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_464 bl[464] br[464] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_465 bl[465] br[465] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_466 bl[466] br[466] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_467 bl[467] br[467] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_468 bl[468] br[468] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_469 bl[469] br[469] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_470 bl[470] br[470] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_471 bl[471] br[471] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_472 bl[472] br[472] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_473 bl[473] br[473] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_474 bl[474] br[474] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_475 bl[475] br[475] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_476 bl[476] br[476] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_477 bl[477] br[477] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_478 bl[478] br[478] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_479 bl[479] br[479] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_480 bl[480] br[480] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_481 bl[481] br[481] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_482 bl[482] br[482] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_483 bl[483] br[483] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_484 bl[484] br[484] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_485 bl[485] br[485] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_486 bl[486] br[486] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_487 bl[487] br[487] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_488 bl[488] br[488] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_489 bl[489] br[489] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_490 bl[490] br[490] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_491 bl[491] br[491] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_492 bl[492] br[492] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_493 bl[493] br[493] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_494 bl[494] br[494] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_495 bl[495] br[495] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_496 bl[496] br[496] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_497 bl[497] br[497] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_498 bl[498] br[498] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_499 bl[499] br[499] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_500 bl[500] br[500] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_501 bl[501] br[501] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_502 bl[502] br[502] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_503 bl[503] br[503] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_504 bl[504] br[504] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_505 bl[505] br[505] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_506 bl[506] br[506] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_507 bl[507] br[507] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_508 bl[508] br[508] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_509 bl[509] br[509] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_510 bl[510] br[510] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_57_511 bl[511] br[511] vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xcell_58_0 bl[0] br[0] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_1 bl[1] br[1] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_2 bl[2] br[2] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_3 bl[3] br[3] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_4 bl[4] br[4] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_5 bl[5] br[5] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_6 bl[6] br[6] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_7 bl[7] br[7] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_8 bl[8] br[8] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_9 bl[9] br[9] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_10 bl[10] br[10] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_11 bl[11] br[11] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_12 bl[12] br[12] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_13 bl[13] br[13] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_14 bl[14] br[14] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_15 bl[15] br[15] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_16 bl[16] br[16] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_17 bl[17] br[17] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_18 bl[18] br[18] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_19 bl[19] br[19] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_20 bl[20] br[20] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_21 bl[21] br[21] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_22 bl[22] br[22] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_23 bl[23] br[23] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_24 bl[24] br[24] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_25 bl[25] br[25] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_26 bl[26] br[26] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_27 bl[27] br[27] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_28 bl[28] br[28] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_29 bl[29] br[29] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_30 bl[30] br[30] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_31 bl[31] br[31] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_32 bl[32] br[32] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_33 bl[33] br[33] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_34 bl[34] br[34] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_35 bl[35] br[35] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_36 bl[36] br[36] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_37 bl[37] br[37] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_38 bl[38] br[38] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_39 bl[39] br[39] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_40 bl[40] br[40] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_41 bl[41] br[41] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_42 bl[42] br[42] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_43 bl[43] br[43] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_44 bl[44] br[44] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_45 bl[45] br[45] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_46 bl[46] br[46] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_47 bl[47] br[47] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_48 bl[48] br[48] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_49 bl[49] br[49] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_50 bl[50] br[50] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_51 bl[51] br[51] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_52 bl[52] br[52] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_53 bl[53] br[53] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_54 bl[54] br[54] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_55 bl[55] br[55] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_56 bl[56] br[56] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_57 bl[57] br[57] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_58 bl[58] br[58] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_59 bl[59] br[59] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_60 bl[60] br[60] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_61 bl[61] br[61] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_62 bl[62] br[62] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_63 bl[63] br[63] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_64 bl[64] br[64] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_65 bl[65] br[65] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_66 bl[66] br[66] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_67 bl[67] br[67] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_68 bl[68] br[68] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_69 bl[69] br[69] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_70 bl[70] br[70] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_71 bl[71] br[71] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_72 bl[72] br[72] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_73 bl[73] br[73] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_74 bl[74] br[74] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_75 bl[75] br[75] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_76 bl[76] br[76] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_77 bl[77] br[77] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_78 bl[78] br[78] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_79 bl[79] br[79] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_80 bl[80] br[80] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_81 bl[81] br[81] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_82 bl[82] br[82] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_83 bl[83] br[83] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_84 bl[84] br[84] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_85 bl[85] br[85] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_86 bl[86] br[86] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_87 bl[87] br[87] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_88 bl[88] br[88] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_89 bl[89] br[89] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_90 bl[90] br[90] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_91 bl[91] br[91] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_92 bl[92] br[92] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_93 bl[93] br[93] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_94 bl[94] br[94] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_95 bl[95] br[95] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_96 bl[96] br[96] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_97 bl[97] br[97] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_98 bl[98] br[98] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_99 bl[99] br[99] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_100 bl[100] br[100] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_101 bl[101] br[101] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_102 bl[102] br[102] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_103 bl[103] br[103] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_104 bl[104] br[104] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_105 bl[105] br[105] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_106 bl[106] br[106] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_107 bl[107] br[107] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_108 bl[108] br[108] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_109 bl[109] br[109] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_110 bl[110] br[110] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_111 bl[111] br[111] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_112 bl[112] br[112] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_113 bl[113] br[113] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_114 bl[114] br[114] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_115 bl[115] br[115] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_116 bl[116] br[116] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_117 bl[117] br[117] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_118 bl[118] br[118] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_119 bl[119] br[119] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_120 bl[120] br[120] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_121 bl[121] br[121] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_122 bl[122] br[122] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_123 bl[123] br[123] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_124 bl[124] br[124] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_125 bl[125] br[125] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_126 bl[126] br[126] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_127 bl[127] br[127] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_128 bl[128] br[128] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_129 bl[129] br[129] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_130 bl[130] br[130] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_131 bl[131] br[131] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_132 bl[132] br[132] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_133 bl[133] br[133] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_134 bl[134] br[134] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_135 bl[135] br[135] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_136 bl[136] br[136] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_137 bl[137] br[137] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_138 bl[138] br[138] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_139 bl[139] br[139] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_140 bl[140] br[140] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_141 bl[141] br[141] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_142 bl[142] br[142] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_143 bl[143] br[143] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_144 bl[144] br[144] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_145 bl[145] br[145] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_146 bl[146] br[146] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_147 bl[147] br[147] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_148 bl[148] br[148] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_149 bl[149] br[149] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_150 bl[150] br[150] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_151 bl[151] br[151] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_152 bl[152] br[152] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_153 bl[153] br[153] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_154 bl[154] br[154] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_155 bl[155] br[155] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_156 bl[156] br[156] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_157 bl[157] br[157] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_158 bl[158] br[158] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_159 bl[159] br[159] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_160 bl[160] br[160] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_161 bl[161] br[161] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_162 bl[162] br[162] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_163 bl[163] br[163] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_164 bl[164] br[164] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_165 bl[165] br[165] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_166 bl[166] br[166] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_167 bl[167] br[167] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_168 bl[168] br[168] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_169 bl[169] br[169] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_170 bl[170] br[170] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_171 bl[171] br[171] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_172 bl[172] br[172] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_173 bl[173] br[173] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_174 bl[174] br[174] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_175 bl[175] br[175] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_176 bl[176] br[176] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_177 bl[177] br[177] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_178 bl[178] br[178] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_179 bl[179] br[179] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_180 bl[180] br[180] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_181 bl[181] br[181] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_182 bl[182] br[182] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_183 bl[183] br[183] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_184 bl[184] br[184] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_185 bl[185] br[185] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_186 bl[186] br[186] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_187 bl[187] br[187] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_188 bl[188] br[188] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_189 bl[189] br[189] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_190 bl[190] br[190] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_191 bl[191] br[191] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_192 bl[192] br[192] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_193 bl[193] br[193] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_194 bl[194] br[194] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_195 bl[195] br[195] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_196 bl[196] br[196] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_197 bl[197] br[197] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_198 bl[198] br[198] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_199 bl[199] br[199] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_200 bl[200] br[200] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_201 bl[201] br[201] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_202 bl[202] br[202] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_203 bl[203] br[203] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_204 bl[204] br[204] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_205 bl[205] br[205] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_206 bl[206] br[206] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_207 bl[207] br[207] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_208 bl[208] br[208] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_209 bl[209] br[209] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_210 bl[210] br[210] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_211 bl[211] br[211] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_212 bl[212] br[212] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_213 bl[213] br[213] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_214 bl[214] br[214] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_215 bl[215] br[215] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_216 bl[216] br[216] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_217 bl[217] br[217] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_218 bl[218] br[218] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_219 bl[219] br[219] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_220 bl[220] br[220] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_221 bl[221] br[221] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_222 bl[222] br[222] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_223 bl[223] br[223] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_224 bl[224] br[224] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_225 bl[225] br[225] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_226 bl[226] br[226] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_227 bl[227] br[227] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_228 bl[228] br[228] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_229 bl[229] br[229] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_230 bl[230] br[230] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_231 bl[231] br[231] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_232 bl[232] br[232] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_233 bl[233] br[233] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_234 bl[234] br[234] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_235 bl[235] br[235] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_236 bl[236] br[236] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_237 bl[237] br[237] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_238 bl[238] br[238] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_239 bl[239] br[239] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_240 bl[240] br[240] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_241 bl[241] br[241] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_242 bl[242] br[242] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_243 bl[243] br[243] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_244 bl[244] br[244] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_245 bl[245] br[245] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_246 bl[246] br[246] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_247 bl[247] br[247] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_248 bl[248] br[248] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_249 bl[249] br[249] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_250 bl[250] br[250] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_251 bl[251] br[251] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_252 bl[252] br[252] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_253 bl[253] br[253] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_254 bl[254] br[254] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_255 bl[255] br[255] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_256 bl[256] br[256] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_257 bl[257] br[257] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_258 bl[258] br[258] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_259 bl[259] br[259] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_260 bl[260] br[260] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_261 bl[261] br[261] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_262 bl[262] br[262] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_263 bl[263] br[263] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_264 bl[264] br[264] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_265 bl[265] br[265] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_266 bl[266] br[266] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_267 bl[267] br[267] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_268 bl[268] br[268] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_269 bl[269] br[269] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_270 bl[270] br[270] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_271 bl[271] br[271] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_272 bl[272] br[272] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_273 bl[273] br[273] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_274 bl[274] br[274] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_275 bl[275] br[275] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_276 bl[276] br[276] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_277 bl[277] br[277] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_278 bl[278] br[278] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_279 bl[279] br[279] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_280 bl[280] br[280] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_281 bl[281] br[281] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_282 bl[282] br[282] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_283 bl[283] br[283] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_284 bl[284] br[284] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_285 bl[285] br[285] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_286 bl[286] br[286] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_287 bl[287] br[287] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_288 bl[288] br[288] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_289 bl[289] br[289] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_290 bl[290] br[290] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_291 bl[291] br[291] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_292 bl[292] br[292] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_293 bl[293] br[293] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_294 bl[294] br[294] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_295 bl[295] br[295] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_296 bl[296] br[296] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_297 bl[297] br[297] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_298 bl[298] br[298] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_299 bl[299] br[299] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_300 bl[300] br[300] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_301 bl[301] br[301] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_302 bl[302] br[302] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_303 bl[303] br[303] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_304 bl[304] br[304] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_305 bl[305] br[305] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_306 bl[306] br[306] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_307 bl[307] br[307] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_308 bl[308] br[308] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_309 bl[309] br[309] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_310 bl[310] br[310] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_311 bl[311] br[311] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_312 bl[312] br[312] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_313 bl[313] br[313] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_314 bl[314] br[314] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_315 bl[315] br[315] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_316 bl[316] br[316] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_317 bl[317] br[317] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_318 bl[318] br[318] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_319 bl[319] br[319] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_320 bl[320] br[320] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_321 bl[321] br[321] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_322 bl[322] br[322] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_323 bl[323] br[323] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_324 bl[324] br[324] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_325 bl[325] br[325] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_326 bl[326] br[326] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_327 bl[327] br[327] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_328 bl[328] br[328] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_329 bl[329] br[329] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_330 bl[330] br[330] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_331 bl[331] br[331] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_332 bl[332] br[332] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_333 bl[333] br[333] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_334 bl[334] br[334] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_335 bl[335] br[335] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_336 bl[336] br[336] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_337 bl[337] br[337] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_338 bl[338] br[338] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_339 bl[339] br[339] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_340 bl[340] br[340] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_341 bl[341] br[341] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_342 bl[342] br[342] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_343 bl[343] br[343] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_344 bl[344] br[344] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_345 bl[345] br[345] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_346 bl[346] br[346] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_347 bl[347] br[347] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_348 bl[348] br[348] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_349 bl[349] br[349] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_350 bl[350] br[350] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_351 bl[351] br[351] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_352 bl[352] br[352] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_353 bl[353] br[353] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_354 bl[354] br[354] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_355 bl[355] br[355] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_356 bl[356] br[356] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_357 bl[357] br[357] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_358 bl[358] br[358] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_359 bl[359] br[359] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_360 bl[360] br[360] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_361 bl[361] br[361] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_362 bl[362] br[362] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_363 bl[363] br[363] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_364 bl[364] br[364] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_365 bl[365] br[365] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_366 bl[366] br[366] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_367 bl[367] br[367] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_368 bl[368] br[368] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_369 bl[369] br[369] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_370 bl[370] br[370] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_371 bl[371] br[371] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_372 bl[372] br[372] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_373 bl[373] br[373] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_374 bl[374] br[374] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_375 bl[375] br[375] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_376 bl[376] br[376] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_377 bl[377] br[377] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_378 bl[378] br[378] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_379 bl[379] br[379] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_380 bl[380] br[380] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_381 bl[381] br[381] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_382 bl[382] br[382] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_383 bl[383] br[383] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_384 bl[384] br[384] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_385 bl[385] br[385] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_386 bl[386] br[386] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_387 bl[387] br[387] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_388 bl[388] br[388] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_389 bl[389] br[389] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_390 bl[390] br[390] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_391 bl[391] br[391] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_392 bl[392] br[392] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_393 bl[393] br[393] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_394 bl[394] br[394] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_395 bl[395] br[395] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_396 bl[396] br[396] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_397 bl[397] br[397] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_398 bl[398] br[398] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_399 bl[399] br[399] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_400 bl[400] br[400] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_401 bl[401] br[401] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_402 bl[402] br[402] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_403 bl[403] br[403] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_404 bl[404] br[404] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_405 bl[405] br[405] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_406 bl[406] br[406] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_407 bl[407] br[407] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_408 bl[408] br[408] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_409 bl[409] br[409] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_410 bl[410] br[410] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_411 bl[411] br[411] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_412 bl[412] br[412] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_413 bl[413] br[413] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_414 bl[414] br[414] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_415 bl[415] br[415] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_416 bl[416] br[416] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_417 bl[417] br[417] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_418 bl[418] br[418] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_419 bl[419] br[419] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_420 bl[420] br[420] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_421 bl[421] br[421] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_422 bl[422] br[422] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_423 bl[423] br[423] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_424 bl[424] br[424] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_425 bl[425] br[425] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_426 bl[426] br[426] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_427 bl[427] br[427] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_428 bl[428] br[428] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_429 bl[429] br[429] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_430 bl[430] br[430] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_431 bl[431] br[431] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_432 bl[432] br[432] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_433 bl[433] br[433] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_434 bl[434] br[434] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_435 bl[435] br[435] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_436 bl[436] br[436] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_437 bl[437] br[437] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_438 bl[438] br[438] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_439 bl[439] br[439] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_440 bl[440] br[440] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_441 bl[441] br[441] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_442 bl[442] br[442] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_443 bl[443] br[443] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_444 bl[444] br[444] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_445 bl[445] br[445] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_446 bl[446] br[446] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_447 bl[447] br[447] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_448 bl[448] br[448] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_449 bl[449] br[449] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_450 bl[450] br[450] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_451 bl[451] br[451] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_452 bl[452] br[452] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_453 bl[453] br[453] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_454 bl[454] br[454] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_455 bl[455] br[455] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_456 bl[456] br[456] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_457 bl[457] br[457] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_458 bl[458] br[458] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_459 bl[459] br[459] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_460 bl[460] br[460] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_461 bl[461] br[461] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_462 bl[462] br[462] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_463 bl[463] br[463] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_464 bl[464] br[464] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_465 bl[465] br[465] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_466 bl[466] br[466] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_467 bl[467] br[467] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_468 bl[468] br[468] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_469 bl[469] br[469] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_470 bl[470] br[470] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_471 bl[471] br[471] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_472 bl[472] br[472] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_473 bl[473] br[473] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_474 bl[474] br[474] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_475 bl[475] br[475] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_476 bl[476] br[476] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_477 bl[477] br[477] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_478 bl[478] br[478] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_479 bl[479] br[479] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_480 bl[480] br[480] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_481 bl[481] br[481] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_482 bl[482] br[482] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_483 bl[483] br[483] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_484 bl[484] br[484] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_485 bl[485] br[485] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_486 bl[486] br[486] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_487 bl[487] br[487] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_488 bl[488] br[488] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_489 bl[489] br[489] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_490 bl[490] br[490] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_491 bl[491] br[491] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_492 bl[492] br[492] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_493 bl[493] br[493] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_494 bl[494] br[494] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_495 bl[495] br[495] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_496 bl[496] br[496] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_497 bl[497] br[497] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_498 bl[498] br[498] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_499 bl[499] br[499] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_500 bl[500] br[500] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_501 bl[501] br[501] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_502 bl[502] br[502] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_503 bl[503] br[503] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_504 bl[504] br[504] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_505 bl[505] br[505] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_506 bl[506] br[506] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_507 bl[507] br[507] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_508 bl[508] br[508] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_509 bl[509] br[509] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_510 bl[510] br[510] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_58_511 bl[511] br[511] vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xcell_59_0 bl[0] br[0] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_1 bl[1] br[1] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_2 bl[2] br[2] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_3 bl[3] br[3] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_4 bl[4] br[4] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_5 bl[5] br[5] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_6 bl[6] br[6] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_7 bl[7] br[7] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_8 bl[8] br[8] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_9 bl[9] br[9] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_10 bl[10] br[10] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_11 bl[11] br[11] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_12 bl[12] br[12] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_13 bl[13] br[13] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_14 bl[14] br[14] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_15 bl[15] br[15] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_16 bl[16] br[16] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_17 bl[17] br[17] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_18 bl[18] br[18] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_19 bl[19] br[19] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_20 bl[20] br[20] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_21 bl[21] br[21] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_22 bl[22] br[22] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_23 bl[23] br[23] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_24 bl[24] br[24] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_25 bl[25] br[25] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_26 bl[26] br[26] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_27 bl[27] br[27] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_28 bl[28] br[28] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_29 bl[29] br[29] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_30 bl[30] br[30] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_31 bl[31] br[31] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_32 bl[32] br[32] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_33 bl[33] br[33] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_34 bl[34] br[34] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_35 bl[35] br[35] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_36 bl[36] br[36] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_37 bl[37] br[37] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_38 bl[38] br[38] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_39 bl[39] br[39] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_40 bl[40] br[40] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_41 bl[41] br[41] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_42 bl[42] br[42] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_43 bl[43] br[43] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_44 bl[44] br[44] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_45 bl[45] br[45] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_46 bl[46] br[46] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_47 bl[47] br[47] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_48 bl[48] br[48] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_49 bl[49] br[49] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_50 bl[50] br[50] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_51 bl[51] br[51] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_52 bl[52] br[52] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_53 bl[53] br[53] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_54 bl[54] br[54] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_55 bl[55] br[55] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_56 bl[56] br[56] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_57 bl[57] br[57] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_58 bl[58] br[58] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_59 bl[59] br[59] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_60 bl[60] br[60] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_61 bl[61] br[61] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_62 bl[62] br[62] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_63 bl[63] br[63] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_64 bl[64] br[64] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_65 bl[65] br[65] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_66 bl[66] br[66] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_67 bl[67] br[67] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_68 bl[68] br[68] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_69 bl[69] br[69] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_70 bl[70] br[70] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_71 bl[71] br[71] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_72 bl[72] br[72] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_73 bl[73] br[73] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_74 bl[74] br[74] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_75 bl[75] br[75] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_76 bl[76] br[76] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_77 bl[77] br[77] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_78 bl[78] br[78] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_79 bl[79] br[79] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_80 bl[80] br[80] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_81 bl[81] br[81] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_82 bl[82] br[82] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_83 bl[83] br[83] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_84 bl[84] br[84] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_85 bl[85] br[85] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_86 bl[86] br[86] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_87 bl[87] br[87] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_88 bl[88] br[88] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_89 bl[89] br[89] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_90 bl[90] br[90] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_91 bl[91] br[91] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_92 bl[92] br[92] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_93 bl[93] br[93] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_94 bl[94] br[94] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_95 bl[95] br[95] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_96 bl[96] br[96] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_97 bl[97] br[97] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_98 bl[98] br[98] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_99 bl[99] br[99] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_100 bl[100] br[100] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_101 bl[101] br[101] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_102 bl[102] br[102] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_103 bl[103] br[103] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_104 bl[104] br[104] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_105 bl[105] br[105] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_106 bl[106] br[106] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_107 bl[107] br[107] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_108 bl[108] br[108] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_109 bl[109] br[109] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_110 bl[110] br[110] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_111 bl[111] br[111] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_112 bl[112] br[112] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_113 bl[113] br[113] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_114 bl[114] br[114] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_115 bl[115] br[115] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_116 bl[116] br[116] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_117 bl[117] br[117] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_118 bl[118] br[118] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_119 bl[119] br[119] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_120 bl[120] br[120] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_121 bl[121] br[121] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_122 bl[122] br[122] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_123 bl[123] br[123] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_124 bl[124] br[124] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_125 bl[125] br[125] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_126 bl[126] br[126] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_127 bl[127] br[127] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_128 bl[128] br[128] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_129 bl[129] br[129] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_130 bl[130] br[130] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_131 bl[131] br[131] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_132 bl[132] br[132] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_133 bl[133] br[133] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_134 bl[134] br[134] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_135 bl[135] br[135] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_136 bl[136] br[136] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_137 bl[137] br[137] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_138 bl[138] br[138] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_139 bl[139] br[139] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_140 bl[140] br[140] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_141 bl[141] br[141] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_142 bl[142] br[142] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_143 bl[143] br[143] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_144 bl[144] br[144] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_145 bl[145] br[145] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_146 bl[146] br[146] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_147 bl[147] br[147] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_148 bl[148] br[148] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_149 bl[149] br[149] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_150 bl[150] br[150] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_151 bl[151] br[151] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_152 bl[152] br[152] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_153 bl[153] br[153] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_154 bl[154] br[154] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_155 bl[155] br[155] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_156 bl[156] br[156] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_157 bl[157] br[157] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_158 bl[158] br[158] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_159 bl[159] br[159] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_160 bl[160] br[160] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_161 bl[161] br[161] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_162 bl[162] br[162] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_163 bl[163] br[163] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_164 bl[164] br[164] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_165 bl[165] br[165] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_166 bl[166] br[166] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_167 bl[167] br[167] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_168 bl[168] br[168] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_169 bl[169] br[169] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_170 bl[170] br[170] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_171 bl[171] br[171] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_172 bl[172] br[172] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_173 bl[173] br[173] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_174 bl[174] br[174] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_175 bl[175] br[175] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_176 bl[176] br[176] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_177 bl[177] br[177] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_178 bl[178] br[178] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_179 bl[179] br[179] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_180 bl[180] br[180] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_181 bl[181] br[181] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_182 bl[182] br[182] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_183 bl[183] br[183] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_184 bl[184] br[184] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_185 bl[185] br[185] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_186 bl[186] br[186] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_187 bl[187] br[187] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_188 bl[188] br[188] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_189 bl[189] br[189] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_190 bl[190] br[190] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_191 bl[191] br[191] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_192 bl[192] br[192] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_193 bl[193] br[193] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_194 bl[194] br[194] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_195 bl[195] br[195] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_196 bl[196] br[196] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_197 bl[197] br[197] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_198 bl[198] br[198] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_199 bl[199] br[199] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_200 bl[200] br[200] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_201 bl[201] br[201] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_202 bl[202] br[202] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_203 bl[203] br[203] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_204 bl[204] br[204] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_205 bl[205] br[205] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_206 bl[206] br[206] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_207 bl[207] br[207] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_208 bl[208] br[208] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_209 bl[209] br[209] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_210 bl[210] br[210] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_211 bl[211] br[211] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_212 bl[212] br[212] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_213 bl[213] br[213] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_214 bl[214] br[214] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_215 bl[215] br[215] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_216 bl[216] br[216] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_217 bl[217] br[217] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_218 bl[218] br[218] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_219 bl[219] br[219] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_220 bl[220] br[220] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_221 bl[221] br[221] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_222 bl[222] br[222] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_223 bl[223] br[223] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_224 bl[224] br[224] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_225 bl[225] br[225] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_226 bl[226] br[226] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_227 bl[227] br[227] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_228 bl[228] br[228] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_229 bl[229] br[229] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_230 bl[230] br[230] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_231 bl[231] br[231] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_232 bl[232] br[232] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_233 bl[233] br[233] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_234 bl[234] br[234] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_235 bl[235] br[235] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_236 bl[236] br[236] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_237 bl[237] br[237] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_238 bl[238] br[238] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_239 bl[239] br[239] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_240 bl[240] br[240] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_241 bl[241] br[241] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_242 bl[242] br[242] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_243 bl[243] br[243] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_244 bl[244] br[244] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_245 bl[245] br[245] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_246 bl[246] br[246] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_247 bl[247] br[247] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_248 bl[248] br[248] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_249 bl[249] br[249] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_250 bl[250] br[250] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_251 bl[251] br[251] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_252 bl[252] br[252] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_253 bl[253] br[253] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_254 bl[254] br[254] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_255 bl[255] br[255] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_256 bl[256] br[256] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_257 bl[257] br[257] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_258 bl[258] br[258] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_259 bl[259] br[259] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_260 bl[260] br[260] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_261 bl[261] br[261] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_262 bl[262] br[262] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_263 bl[263] br[263] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_264 bl[264] br[264] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_265 bl[265] br[265] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_266 bl[266] br[266] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_267 bl[267] br[267] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_268 bl[268] br[268] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_269 bl[269] br[269] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_270 bl[270] br[270] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_271 bl[271] br[271] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_272 bl[272] br[272] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_273 bl[273] br[273] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_274 bl[274] br[274] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_275 bl[275] br[275] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_276 bl[276] br[276] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_277 bl[277] br[277] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_278 bl[278] br[278] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_279 bl[279] br[279] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_280 bl[280] br[280] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_281 bl[281] br[281] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_282 bl[282] br[282] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_283 bl[283] br[283] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_284 bl[284] br[284] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_285 bl[285] br[285] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_286 bl[286] br[286] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_287 bl[287] br[287] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_288 bl[288] br[288] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_289 bl[289] br[289] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_290 bl[290] br[290] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_291 bl[291] br[291] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_292 bl[292] br[292] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_293 bl[293] br[293] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_294 bl[294] br[294] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_295 bl[295] br[295] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_296 bl[296] br[296] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_297 bl[297] br[297] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_298 bl[298] br[298] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_299 bl[299] br[299] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_300 bl[300] br[300] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_301 bl[301] br[301] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_302 bl[302] br[302] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_303 bl[303] br[303] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_304 bl[304] br[304] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_305 bl[305] br[305] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_306 bl[306] br[306] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_307 bl[307] br[307] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_308 bl[308] br[308] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_309 bl[309] br[309] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_310 bl[310] br[310] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_311 bl[311] br[311] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_312 bl[312] br[312] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_313 bl[313] br[313] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_314 bl[314] br[314] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_315 bl[315] br[315] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_316 bl[316] br[316] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_317 bl[317] br[317] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_318 bl[318] br[318] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_319 bl[319] br[319] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_320 bl[320] br[320] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_321 bl[321] br[321] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_322 bl[322] br[322] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_323 bl[323] br[323] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_324 bl[324] br[324] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_325 bl[325] br[325] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_326 bl[326] br[326] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_327 bl[327] br[327] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_328 bl[328] br[328] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_329 bl[329] br[329] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_330 bl[330] br[330] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_331 bl[331] br[331] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_332 bl[332] br[332] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_333 bl[333] br[333] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_334 bl[334] br[334] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_335 bl[335] br[335] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_336 bl[336] br[336] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_337 bl[337] br[337] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_338 bl[338] br[338] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_339 bl[339] br[339] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_340 bl[340] br[340] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_341 bl[341] br[341] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_342 bl[342] br[342] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_343 bl[343] br[343] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_344 bl[344] br[344] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_345 bl[345] br[345] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_346 bl[346] br[346] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_347 bl[347] br[347] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_348 bl[348] br[348] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_349 bl[349] br[349] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_350 bl[350] br[350] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_351 bl[351] br[351] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_352 bl[352] br[352] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_353 bl[353] br[353] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_354 bl[354] br[354] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_355 bl[355] br[355] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_356 bl[356] br[356] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_357 bl[357] br[357] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_358 bl[358] br[358] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_359 bl[359] br[359] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_360 bl[360] br[360] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_361 bl[361] br[361] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_362 bl[362] br[362] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_363 bl[363] br[363] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_364 bl[364] br[364] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_365 bl[365] br[365] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_366 bl[366] br[366] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_367 bl[367] br[367] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_368 bl[368] br[368] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_369 bl[369] br[369] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_370 bl[370] br[370] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_371 bl[371] br[371] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_372 bl[372] br[372] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_373 bl[373] br[373] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_374 bl[374] br[374] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_375 bl[375] br[375] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_376 bl[376] br[376] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_377 bl[377] br[377] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_378 bl[378] br[378] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_379 bl[379] br[379] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_380 bl[380] br[380] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_381 bl[381] br[381] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_382 bl[382] br[382] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_383 bl[383] br[383] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_384 bl[384] br[384] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_385 bl[385] br[385] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_386 bl[386] br[386] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_387 bl[387] br[387] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_388 bl[388] br[388] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_389 bl[389] br[389] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_390 bl[390] br[390] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_391 bl[391] br[391] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_392 bl[392] br[392] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_393 bl[393] br[393] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_394 bl[394] br[394] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_395 bl[395] br[395] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_396 bl[396] br[396] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_397 bl[397] br[397] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_398 bl[398] br[398] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_399 bl[399] br[399] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_400 bl[400] br[400] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_401 bl[401] br[401] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_402 bl[402] br[402] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_403 bl[403] br[403] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_404 bl[404] br[404] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_405 bl[405] br[405] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_406 bl[406] br[406] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_407 bl[407] br[407] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_408 bl[408] br[408] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_409 bl[409] br[409] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_410 bl[410] br[410] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_411 bl[411] br[411] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_412 bl[412] br[412] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_413 bl[413] br[413] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_414 bl[414] br[414] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_415 bl[415] br[415] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_416 bl[416] br[416] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_417 bl[417] br[417] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_418 bl[418] br[418] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_419 bl[419] br[419] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_420 bl[420] br[420] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_421 bl[421] br[421] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_422 bl[422] br[422] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_423 bl[423] br[423] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_424 bl[424] br[424] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_425 bl[425] br[425] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_426 bl[426] br[426] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_427 bl[427] br[427] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_428 bl[428] br[428] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_429 bl[429] br[429] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_430 bl[430] br[430] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_431 bl[431] br[431] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_432 bl[432] br[432] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_433 bl[433] br[433] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_434 bl[434] br[434] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_435 bl[435] br[435] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_436 bl[436] br[436] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_437 bl[437] br[437] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_438 bl[438] br[438] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_439 bl[439] br[439] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_440 bl[440] br[440] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_441 bl[441] br[441] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_442 bl[442] br[442] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_443 bl[443] br[443] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_444 bl[444] br[444] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_445 bl[445] br[445] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_446 bl[446] br[446] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_447 bl[447] br[447] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_448 bl[448] br[448] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_449 bl[449] br[449] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_450 bl[450] br[450] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_451 bl[451] br[451] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_452 bl[452] br[452] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_453 bl[453] br[453] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_454 bl[454] br[454] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_455 bl[455] br[455] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_456 bl[456] br[456] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_457 bl[457] br[457] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_458 bl[458] br[458] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_459 bl[459] br[459] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_460 bl[460] br[460] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_461 bl[461] br[461] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_462 bl[462] br[462] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_463 bl[463] br[463] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_464 bl[464] br[464] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_465 bl[465] br[465] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_466 bl[466] br[466] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_467 bl[467] br[467] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_468 bl[468] br[468] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_469 bl[469] br[469] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_470 bl[470] br[470] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_471 bl[471] br[471] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_472 bl[472] br[472] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_473 bl[473] br[473] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_474 bl[474] br[474] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_475 bl[475] br[475] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_476 bl[476] br[476] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_477 bl[477] br[477] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_478 bl[478] br[478] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_479 bl[479] br[479] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_480 bl[480] br[480] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_481 bl[481] br[481] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_482 bl[482] br[482] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_483 bl[483] br[483] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_484 bl[484] br[484] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_485 bl[485] br[485] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_486 bl[486] br[486] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_487 bl[487] br[487] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_488 bl[488] br[488] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_489 bl[489] br[489] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_490 bl[490] br[490] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_491 bl[491] br[491] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_492 bl[492] br[492] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_493 bl[493] br[493] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_494 bl[494] br[494] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_495 bl[495] br[495] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_496 bl[496] br[496] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_497 bl[497] br[497] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_498 bl[498] br[498] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_499 bl[499] br[499] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_500 bl[500] br[500] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_501 bl[501] br[501] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_502 bl[502] br[502] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_503 bl[503] br[503] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_504 bl[504] br[504] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_505 bl[505] br[505] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_506 bl[506] br[506] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_507 bl[507] br[507] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_508 bl[508] br[508] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_509 bl[509] br[509] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_510 bl[510] br[510] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_59_511 bl[511] br[511] vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xcell_60_0 bl[0] br[0] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_1 bl[1] br[1] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_2 bl[2] br[2] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_3 bl[3] br[3] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_4 bl[4] br[4] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_5 bl[5] br[5] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_6 bl[6] br[6] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_7 bl[7] br[7] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_8 bl[8] br[8] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_9 bl[9] br[9] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_10 bl[10] br[10] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_11 bl[11] br[11] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_12 bl[12] br[12] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_13 bl[13] br[13] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_14 bl[14] br[14] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_15 bl[15] br[15] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_16 bl[16] br[16] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_17 bl[17] br[17] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_18 bl[18] br[18] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_19 bl[19] br[19] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_20 bl[20] br[20] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_21 bl[21] br[21] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_22 bl[22] br[22] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_23 bl[23] br[23] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_24 bl[24] br[24] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_25 bl[25] br[25] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_26 bl[26] br[26] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_27 bl[27] br[27] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_28 bl[28] br[28] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_29 bl[29] br[29] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_30 bl[30] br[30] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_31 bl[31] br[31] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_32 bl[32] br[32] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_33 bl[33] br[33] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_34 bl[34] br[34] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_35 bl[35] br[35] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_36 bl[36] br[36] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_37 bl[37] br[37] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_38 bl[38] br[38] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_39 bl[39] br[39] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_40 bl[40] br[40] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_41 bl[41] br[41] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_42 bl[42] br[42] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_43 bl[43] br[43] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_44 bl[44] br[44] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_45 bl[45] br[45] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_46 bl[46] br[46] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_47 bl[47] br[47] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_48 bl[48] br[48] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_49 bl[49] br[49] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_50 bl[50] br[50] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_51 bl[51] br[51] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_52 bl[52] br[52] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_53 bl[53] br[53] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_54 bl[54] br[54] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_55 bl[55] br[55] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_56 bl[56] br[56] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_57 bl[57] br[57] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_58 bl[58] br[58] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_59 bl[59] br[59] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_60 bl[60] br[60] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_61 bl[61] br[61] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_62 bl[62] br[62] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_63 bl[63] br[63] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_64 bl[64] br[64] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_65 bl[65] br[65] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_66 bl[66] br[66] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_67 bl[67] br[67] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_68 bl[68] br[68] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_69 bl[69] br[69] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_70 bl[70] br[70] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_71 bl[71] br[71] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_72 bl[72] br[72] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_73 bl[73] br[73] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_74 bl[74] br[74] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_75 bl[75] br[75] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_76 bl[76] br[76] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_77 bl[77] br[77] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_78 bl[78] br[78] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_79 bl[79] br[79] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_80 bl[80] br[80] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_81 bl[81] br[81] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_82 bl[82] br[82] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_83 bl[83] br[83] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_84 bl[84] br[84] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_85 bl[85] br[85] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_86 bl[86] br[86] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_87 bl[87] br[87] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_88 bl[88] br[88] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_89 bl[89] br[89] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_90 bl[90] br[90] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_91 bl[91] br[91] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_92 bl[92] br[92] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_93 bl[93] br[93] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_94 bl[94] br[94] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_95 bl[95] br[95] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_96 bl[96] br[96] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_97 bl[97] br[97] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_98 bl[98] br[98] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_99 bl[99] br[99] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_100 bl[100] br[100] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_101 bl[101] br[101] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_102 bl[102] br[102] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_103 bl[103] br[103] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_104 bl[104] br[104] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_105 bl[105] br[105] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_106 bl[106] br[106] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_107 bl[107] br[107] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_108 bl[108] br[108] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_109 bl[109] br[109] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_110 bl[110] br[110] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_111 bl[111] br[111] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_112 bl[112] br[112] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_113 bl[113] br[113] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_114 bl[114] br[114] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_115 bl[115] br[115] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_116 bl[116] br[116] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_117 bl[117] br[117] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_118 bl[118] br[118] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_119 bl[119] br[119] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_120 bl[120] br[120] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_121 bl[121] br[121] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_122 bl[122] br[122] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_123 bl[123] br[123] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_124 bl[124] br[124] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_125 bl[125] br[125] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_126 bl[126] br[126] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_127 bl[127] br[127] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_128 bl[128] br[128] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_129 bl[129] br[129] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_130 bl[130] br[130] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_131 bl[131] br[131] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_132 bl[132] br[132] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_133 bl[133] br[133] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_134 bl[134] br[134] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_135 bl[135] br[135] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_136 bl[136] br[136] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_137 bl[137] br[137] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_138 bl[138] br[138] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_139 bl[139] br[139] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_140 bl[140] br[140] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_141 bl[141] br[141] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_142 bl[142] br[142] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_143 bl[143] br[143] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_144 bl[144] br[144] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_145 bl[145] br[145] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_146 bl[146] br[146] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_147 bl[147] br[147] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_148 bl[148] br[148] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_149 bl[149] br[149] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_150 bl[150] br[150] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_151 bl[151] br[151] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_152 bl[152] br[152] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_153 bl[153] br[153] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_154 bl[154] br[154] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_155 bl[155] br[155] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_156 bl[156] br[156] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_157 bl[157] br[157] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_158 bl[158] br[158] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_159 bl[159] br[159] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_160 bl[160] br[160] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_161 bl[161] br[161] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_162 bl[162] br[162] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_163 bl[163] br[163] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_164 bl[164] br[164] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_165 bl[165] br[165] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_166 bl[166] br[166] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_167 bl[167] br[167] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_168 bl[168] br[168] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_169 bl[169] br[169] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_170 bl[170] br[170] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_171 bl[171] br[171] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_172 bl[172] br[172] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_173 bl[173] br[173] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_174 bl[174] br[174] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_175 bl[175] br[175] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_176 bl[176] br[176] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_177 bl[177] br[177] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_178 bl[178] br[178] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_179 bl[179] br[179] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_180 bl[180] br[180] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_181 bl[181] br[181] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_182 bl[182] br[182] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_183 bl[183] br[183] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_184 bl[184] br[184] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_185 bl[185] br[185] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_186 bl[186] br[186] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_187 bl[187] br[187] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_188 bl[188] br[188] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_189 bl[189] br[189] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_190 bl[190] br[190] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_191 bl[191] br[191] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_192 bl[192] br[192] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_193 bl[193] br[193] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_194 bl[194] br[194] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_195 bl[195] br[195] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_196 bl[196] br[196] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_197 bl[197] br[197] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_198 bl[198] br[198] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_199 bl[199] br[199] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_200 bl[200] br[200] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_201 bl[201] br[201] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_202 bl[202] br[202] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_203 bl[203] br[203] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_204 bl[204] br[204] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_205 bl[205] br[205] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_206 bl[206] br[206] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_207 bl[207] br[207] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_208 bl[208] br[208] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_209 bl[209] br[209] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_210 bl[210] br[210] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_211 bl[211] br[211] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_212 bl[212] br[212] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_213 bl[213] br[213] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_214 bl[214] br[214] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_215 bl[215] br[215] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_216 bl[216] br[216] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_217 bl[217] br[217] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_218 bl[218] br[218] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_219 bl[219] br[219] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_220 bl[220] br[220] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_221 bl[221] br[221] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_222 bl[222] br[222] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_223 bl[223] br[223] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_224 bl[224] br[224] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_225 bl[225] br[225] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_226 bl[226] br[226] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_227 bl[227] br[227] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_228 bl[228] br[228] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_229 bl[229] br[229] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_230 bl[230] br[230] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_231 bl[231] br[231] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_232 bl[232] br[232] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_233 bl[233] br[233] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_234 bl[234] br[234] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_235 bl[235] br[235] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_236 bl[236] br[236] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_237 bl[237] br[237] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_238 bl[238] br[238] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_239 bl[239] br[239] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_240 bl[240] br[240] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_241 bl[241] br[241] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_242 bl[242] br[242] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_243 bl[243] br[243] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_244 bl[244] br[244] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_245 bl[245] br[245] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_246 bl[246] br[246] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_247 bl[247] br[247] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_248 bl[248] br[248] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_249 bl[249] br[249] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_250 bl[250] br[250] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_251 bl[251] br[251] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_252 bl[252] br[252] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_253 bl[253] br[253] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_254 bl[254] br[254] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_255 bl[255] br[255] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_256 bl[256] br[256] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_257 bl[257] br[257] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_258 bl[258] br[258] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_259 bl[259] br[259] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_260 bl[260] br[260] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_261 bl[261] br[261] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_262 bl[262] br[262] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_263 bl[263] br[263] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_264 bl[264] br[264] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_265 bl[265] br[265] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_266 bl[266] br[266] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_267 bl[267] br[267] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_268 bl[268] br[268] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_269 bl[269] br[269] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_270 bl[270] br[270] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_271 bl[271] br[271] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_272 bl[272] br[272] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_273 bl[273] br[273] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_274 bl[274] br[274] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_275 bl[275] br[275] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_276 bl[276] br[276] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_277 bl[277] br[277] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_278 bl[278] br[278] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_279 bl[279] br[279] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_280 bl[280] br[280] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_281 bl[281] br[281] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_282 bl[282] br[282] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_283 bl[283] br[283] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_284 bl[284] br[284] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_285 bl[285] br[285] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_286 bl[286] br[286] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_287 bl[287] br[287] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_288 bl[288] br[288] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_289 bl[289] br[289] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_290 bl[290] br[290] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_291 bl[291] br[291] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_292 bl[292] br[292] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_293 bl[293] br[293] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_294 bl[294] br[294] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_295 bl[295] br[295] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_296 bl[296] br[296] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_297 bl[297] br[297] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_298 bl[298] br[298] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_299 bl[299] br[299] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_300 bl[300] br[300] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_301 bl[301] br[301] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_302 bl[302] br[302] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_303 bl[303] br[303] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_304 bl[304] br[304] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_305 bl[305] br[305] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_306 bl[306] br[306] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_307 bl[307] br[307] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_308 bl[308] br[308] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_309 bl[309] br[309] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_310 bl[310] br[310] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_311 bl[311] br[311] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_312 bl[312] br[312] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_313 bl[313] br[313] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_314 bl[314] br[314] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_315 bl[315] br[315] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_316 bl[316] br[316] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_317 bl[317] br[317] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_318 bl[318] br[318] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_319 bl[319] br[319] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_320 bl[320] br[320] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_321 bl[321] br[321] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_322 bl[322] br[322] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_323 bl[323] br[323] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_324 bl[324] br[324] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_325 bl[325] br[325] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_326 bl[326] br[326] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_327 bl[327] br[327] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_328 bl[328] br[328] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_329 bl[329] br[329] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_330 bl[330] br[330] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_331 bl[331] br[331] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_332 bl[332] br[332] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_333 bl[333] br[333] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_334 bl[334] br[334] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_335 bl[335] br[335] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_336 bl[336] br[336] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_337 bl[337] br[337] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_338 bl[338] br[338] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_339 bl[339] br[339] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_340 bl[340] br[340] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_341 bl[341] br[341] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_342 bl[342] br[342] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_343 bl[343] br[343] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_344 bl[344] br[344] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_345 bl[345] br[345] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_346 bl[346] br[346] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_347 bl[347] br[347] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_348 bl[348] br[348] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_349 bl[349] br[349] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_350 bl[350] br[350] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_351 bl[351] br[351] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_352 bl[352] br[352] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_353 bl[353] br[353] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_354 bl[354] br[354] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_355 bl[355] br[355] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_356 bl[356] br[356] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_357 bl[357] br[357] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_358 bl[358] br[358] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_359 bl[359] br[359] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_360 bl[360] br[360] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_361 bl[361] br[361] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_362 bl[362] br[362] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_363 bl[363] br[363] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_364 bl[364] br[364] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_365 bl[365] br[365] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_366 bl[366] br[366] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_367 bl[367] br[367] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_368 bl[368] br[368] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_369 bl[369] br[369] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_370 bl[370] br[370] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_371 bl[371] br[371] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_372 bl[372] br[372] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_373 bl[373] br[373] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_374 bl[374] br[374] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_375 bl[375] br[375] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_376 bl[376] br[376] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_377 bl[377] br[377] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_378 bl[378] br[378] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_379 bl[379] br[379] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_380 bl[380] br[380] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_381 bl[381] br[381] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_382 bl[382] br[382] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_383 bl[383] br[383] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_384 bl[384] br[384] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_385 bl[385] br[385] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_386 bl[386] br[386] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_387 bl[387] br[387] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_388 bl[388] br[388] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_389 bl[389] br[389] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_390 bl[390] br[390] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_391 bl[391] br[391] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_392 bl[392] br[392] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_393 bl[393] br[393] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_394 bl[394] br[394] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_395 bl[395] br[395] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_396 bl[396] br[396] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_397 bl[397] br[397] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_398 bl[398] br[398] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_399 bl[399] br[399] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_400 bl[400] br[400] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_401 bl[401] br[401] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_402 bl[402] br[402] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_403 bl[403] br[403] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_404 bl[404] br[404] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_405 bl[405] br[405] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_406 bl[406] br[406] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_407 bl[407] br[407] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_408 bl[408] br[408] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_409 bl[409] br[409] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_410 bl[410] br[410] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_411 bl[411] br[411] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_412 bl[412] br[412] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_413 bl[413] br[413] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_414 bl[414] br[414] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_415 bl[415] br[415] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_416 bl[416] br[416] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_417 bl[417] br[417] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_418 bl[418] br[418] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_419 bl[419] br[419] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_420 bl[420] br[420] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_421 bl[421] br[421] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_422 bl[422] br[422] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_423 bl[423] br[423] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_424 bl[424] br[424] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_425 bl[425] br[425] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_426 bl[426] br[426] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_427 bl[427] br[427] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_428 bl[428] br[428] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_429 bl[429] br[429] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_430 bl[430] br[430] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_431 bl[431] br[431] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_432 bl[432] br[432] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_433 bl[433] br[433] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_434 bl[434] br[434] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_435 bl[435] br[435] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_436 bl[436] br[436] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_437 bl[437] br[437] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_438 bl[438] br[438] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_439 bl[439] br[439] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_440 bl[440] br[440] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_441 bl[441] br[441] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_442 bl[442] br[442] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_443 bl[443] br[443] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_444 bl[444] br[444] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_445 bl[445] br[445] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_446 bl[446] br[446] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_447 bl[447] br[447] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_448 bl[448] br[448] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_449 bl[449] br[449] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_450 bl[450] br[450] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_451 bl[451] br[451] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_452 bl[452] br[452] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_453 bl[453] br[453] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_454 bl[454] br[454] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_455 bl[455] br[455] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_456 bl[456] br[456] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_457 bl[457] br[457] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_458 bl[458] br[458] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_459 bl[459] br[459] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_460 bl[460] br[460] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_461 bl[461] br[461] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_462 bl[462] br[462] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_463 bl[463] br[463] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_464 bl[464] br[464] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_465 bl[465] br[465] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_466 bl[466] br[466] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_467 bl[467] br[467] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_468 bl[468] br[468] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_469 bl[469] br[469] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_470 bl[470] br[470] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_471 bl[471] br[471] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_472 bl[472] br[472] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_473 bl[473] br[473] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_474 bl[474] br[474] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_475 bl[475] br[475] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_476 bl[476] br[476] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_477 bl[477] br[477] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_478 bl[478] br[478] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_479 bl[479] br[479] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_480 bl[480] br[480] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_481 bl[481] br[481] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_482 bl[482] br[482] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_483 bl[483] br[483] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_484 bl[484] br[484] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_485 bl[485] br[485] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_486 bl[486] br[486] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_487 bl[487] br[487] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_488 bl[488] br[488] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_489 bl[489] br[489] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_490 bl[490] br[490] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_491 bl[491] br[491] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_492 bl[492] br[492] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_493 bl[493] br[493] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_494 bl[494] br[494] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_495 bl[495] br[495] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_496 bl[496] br[496] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_497 bl[497] br[497] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_498 bl[498] br[498] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_499 bl[499] br[499] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_500 bl[500] br[500] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_501 bl[501] br[501] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_502 bl[502] br[502] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_503 bl[503] br[503] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_504 bl[504] br[504] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_505 bl[505] br[505] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_506 bl[506] br[506] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_507 bl[507] br[507] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_508 bl[508] br[508] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_509 bl[509] br[509] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_510 bl[510] br[510] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_60_511 bl[511] br[511] vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xcell_61_0 bl[0] br[0] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_1 bl[1] br[1] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_2 bl[2] br[2] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_3 bl[3] br[3] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_4 bl[4] br[4] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_5 bl[5] br[5] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_6 bl[6] br[6] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_7 bl[7] br[7] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_8 bl[8] br[8] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_9 bl[9] br[9] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_10 bl[10] br[10] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_11 bl[11] br[11] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_12 bl[12] br[12] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_13 bl[13] br[13] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_14 bl[14] br[14] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_15 bl[15] br[15] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_16 bl[16] br[16] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_17 bl[17] br[17] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_18 bl[18] br[18] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_19 bl[19] br[19] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_20 bl[20] br[20] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_21 bl[21] br[21] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_22 bl[22] br[22] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_23 bl[23] br[23] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_24 bl[24] br[24] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_25 bl[25] br[25] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_26 bl[26] br[26] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_27 bl[27] br[27] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_28 bl[28] br[28] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_29 bl[29] br[29] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_30 bl[30] br[30] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_31 bl[31] br[31] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_32 bl[32] br[32] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_33 bl[33] br[33] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_34 bl[34] br[34] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_35 bl[35] br[35] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_36 bl[36] br[36] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_37 bl[37] br[37] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_38 bl[38] br[38] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_39 bl[39] br[39] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_40 bl[40] br[40] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_41 bl[41] br[41] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_42 bl[42] br[42] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_43 bl[43] br[43] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_44 bl[44] br[44] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_45 bl[45] br[45] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_46 bl[46] br[46] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_47 bl[47] br[47] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_48 bl[48] br[48] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_49 bl[49] br[49] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_50 bl[50] br[50] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_51 bl[51] br[51] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_52 bl[52] br[52] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_53 bl[53] br[53] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_54 bl[54] br[54] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_55 bl[55] br[55] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_56 bl[56] br[56] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_57 bl[57] br[57] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_58 bl[58] br[58] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_59 bl[59] br[59] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_60 bl[60] br[60] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_61 bl[61] br[61] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_62 bl[62] br[62] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_63 bl[63] br[63] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_64 bl[64] br[64] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_65 bl[65] br[65] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_66 bl[66] br[66] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_67 bl[67] br[67] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_68 bl[68] br[68] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_69 bl[69] br[69] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_70 bl[70] br[70] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_71 bl[71] br[71] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_72 bl[72] br[72] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_73 bl[73] br[73] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_74 bl[74] br[74] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_75 bl[75] br[75] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_76 bl[76] br[76] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_77 bl[77] br[77] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_78 bl[78] br[78] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_79 bl[79] br[79] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_80 bl[80] br[80] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_81 bl[81] br[81] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_82 bl[82] br[82] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_83 bl[83] br[83] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_84 bl[84] br[84] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_85 bl[85] br[85] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_86 bl[86] br[86] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_87 bl[87] br[87] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_88 bl[88] br[88] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_89 bl[89] br[89] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_90 bl[90] br[90] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_91 bl[91] br[91] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_92 bl[92] br[92] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_93 bl[93] br[93] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_94 bl[94] br[94] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_95 bl[95] br[95] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_96 bl[96] br[96] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_97 bl[97] br[97] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_98 bl[98] br[98] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_99 bl[99] br[99] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_100 bl[100] br[100] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_101 bl[101] br[101] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_102 bl[102] br[102] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_103 bl[103] br[103] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_104 bl[104] br[104] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_105 bl[105] br[105] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_106 bl[106] br[106] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_107 bl[107] br[107] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_108 bl[108] br[108] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_109 bl[109] br[109] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_110 bl[110] br[110] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_111 bl[111] br[111] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_112 bl[112] br[112] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_113 bl[113] br[113] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_114 bl[114] br[114] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_115 bl[115] br[115] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_116 bl[116] br[116] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_117 bl[117] br[117] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_118 bl[118] br[118] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_119 bl[119] br[119] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_120 bl[120] br[120] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_121 bl[121] br[121] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_122 bl[122] br[122] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_123 bl[123] br[123] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_124 bl[124] br[124] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_125 bl[125] br[125] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_126 bl[126] br[126] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_127 bl[127] br[127] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_128 bl[128] br[128] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_129 bl[129] br[129] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_130 bl[130] br[130] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_131 bl[131] br[131] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_132 bl[132] br[132] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_133 bl[133] br[133] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_134 bl[134] br[134] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_135 bl[135] br[135] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_136 bl[136] br[136] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_137 bl[137] br[137] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_138 bl[138] br[138] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_139 bl[139] br[139] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_140 bl[140] br[140] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_141 bl[141] br[141] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_142 bl[142] br[142] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_143 bl[143] br[143] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_144 bl[144] br[144] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_145 bl[145] br[145] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_146 bl[146] br[146] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_147 bl[147] br[147] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_148 bl[148] br[148] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_149 bl[149] br[149] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_150 bl[150] br[150] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_151 bl[151] br[151] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_152 bl[152] br[152] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_153 bl[153] br[153] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_154 bl[154] br[154] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_155 bl[155] br[155] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_156 bl[156] br[156] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_157 bl[157] br[157] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_158 bl[158] br[158] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_159 bl[159] br[159] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_160 bl[160] br[160] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_161 bl[161] br[161] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_162 bl[162] br[162] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_163 bl[163] br[163] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_164 bl[164] br[164] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_165 bl[165] br[165] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_166 bl[166] br[166] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_167 bl[167] br[167] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_168 bl[168] br[168] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_169 bl[169] br[169] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_170 bl[170] br[170] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_171 bl[171] br[171] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_172 bl[172] br[172] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_173 bl[173] br[173] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_174 bl[174] br[174] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_175 bl[175] br[175] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_176 bl[176] br[176] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_177 bl[177] br[177] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_178 bl[178] br[178] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_179 bl[179] br[179] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_180 bl[180] br[180] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_181 bl[181] br[181] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_182 bl[182] br[182] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_183 bl[183] br[183] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_184 bl[184] br[184] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_185 bl[185] br[185] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_186 bl[186] br[186] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_187 bl[187] br[187] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_188 bl[188] br[188] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_189 bl[189] br[189] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_190 bl[190] br[190] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_191 bl[191] br[191] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_192 bl[192] br[192] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_193 bl[193] br[193] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_194 bl[194] br[194] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_195 bl[195] br[195] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_196 bl[196] br[196] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_197 bl[197] br[197] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_198 bl[198] br[198] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_199 bl[199] br[199] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_200 bl[200] br[200] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_201 bl[201] br[201] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_202 bl[202] br[202] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_203 bl[203] br[203] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_204 bl[204] br[204] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_205 bl[205] br[205] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_206 bl[206] br[206] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_207 bl[207] br[207] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_208 bl[208] br[208] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_209 bl[209] br[209] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_210 bl[210] br[210] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_211 bl[211] br[211] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_212 bl[212] br[212] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_213 bl[213] br[213] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_214 bl[214] br[214] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_215 bl[215] br[215] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_216 bl[216] br[216] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_217 bl[217] br[217] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_218 bl[218] br[218] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_219 bl[219] br[219] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_220 bl[220] br[220] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_221 bl[221] br[221] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_222 bl[222] br[222] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_223 bl[223] br[223] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_224 bl[224] br[224] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_225 bl[225] br[225] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_226 bl[226] br[226] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_227 bl[227] br[227] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_228 bl[228] br[228] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_229 bl[229] br[229] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_230 bl[230] br[230] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_231 bl[231] br[231] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_232 bl[232] br[232] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_233 bl[233] br[233] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_234 bl[234] br[234] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_235 bl[235] br[235] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_236 bl[236] br[236] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_237 bl[237] br[237] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_238 bl[238] br[238] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_239 bl[239] br[239] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_240 bl[240] br[240] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_241 bl[241] br[241] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_242 bl[242] br[242] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_243 bl[243] br[243] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_244 bl[244] br[244] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_245 bl[245] br[245] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_246 bl[246] br[246] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_247 bl[247] br[247] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_248 bl[248] br[248] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_249 bl[249] br[249] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_250 bl[250] br[250] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_251 bl[251] br[251] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_252 bl[252] br[252] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_253 bl[253] br[253] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_254 bl[254] br[254] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_255 bl[255] br[255] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_256 bl[256] br[256] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_257 bl[257] br[257] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_258 bl[258] br[258] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_259 bl[259] br[259] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_260 bl[260] br[260] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_261 bl[261] br[261] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_262 bl[262] br[262] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_263 bl[263] br[263] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_264 bl[264] br[264] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_265 bl[265] br[265] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_266 bl[266] br[266] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_267 bl[267] br[267] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_268 bl[268] br[268] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_269 bl[269] br[269] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_270 bl[270] br[270] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_271 bl[271] br[271] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_272 bl[272] br[272] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_273 bl[273] br[273] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_274 bl[274] br[274] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_275 bl[275] br[275] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_276 bl[276] br[276] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_277 bl[277] br[277] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_278 bl[278] br[278] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_279 bl[279] br[279] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_280 bl[280] br[280] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_281 bl[281] br[281] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_282 bl[282] br[282] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_283 bl[283] br[283] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_284 bl[284] br[284] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_285 bl[285] br[285] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_286 bl[286] br[286] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_287 bl[287] br[287] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_288 bl[288] br[288] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_289 bl[289] br[289] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_290 bl[290] br[290] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_291 bl[291] br[291] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_292 bl[292] br[292] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_293 bl[293] br[293] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_294 bl[294] br[294] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_295 bl[295] br[295] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_296 bl[296] br[296] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_297 bl[297] br[297] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_298 bl[298] br[298] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_299 bl[299] br[299] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_300 bl[300] br[300] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_301 bl[301] br[301] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_302 bl[302] br[302] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_303 bl[303] br[303] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_304 bl[304] br[304] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_305 bl[305] br[305] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_306 bl[306] br[306] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_307 bl[307] br[307] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_308 bl[308] br[308] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_309 bl[309] br[309] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_310 bl[310] br[310] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_311 bl[311] br[311] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_312 bl[312] br[312] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_313 bl[313] br[313] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_314 bl[314] br[314] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_315 bl[315] br[315] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_316 bl[316] br[316] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_317 bl[317] br[317] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_318 bl[318] br[318] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_319 bl[319] br[319] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_320 bl[320] br[320] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_321 bl[321] br[321] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_322 bl[322] br[322] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_323 bl[323] br[323] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_324 bl[324] br[324] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_325 bl[325] br[325] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_326 bl[326] br[326] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_327 bl[327] br[327] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_328 bl[328] br[328] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_329 bl[329] br[329] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_330 bl[330] br[330] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_331 bl[331] br[331] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_332 bl[332] br[332] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_333 bl[333] br[333] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_334 bl[334] br[334] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_335 bl[335] br[335] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_336 bl[336] br[336] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_337 bl[337] br[337] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_338 bl[338] br[338] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_339 bl[339] br[339] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_340 bl[340] br[340] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_341 bl[341] br[341] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_342 bl[342] br[342] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_343 bl[343] br[343] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_344 bl[344] br[344] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_345 bl[345] br[345] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_346 bl[346] br[346] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_347 bl[347] br[347] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_348 bl[348] br[348] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_349 bl[349] br[349] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_350 bl[350] br[350] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_351 bl[351] br[351] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_352 bl[352] br[352] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_353 bl[353] br[353] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_354 bl[354] br[354] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_355 bl[355] br[355] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_356 bl[356] br[356] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_357 bl[357] br[357] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_358 bl[358] br[358] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_359 bl[359] br[359] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_360 bl[360] br[360] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_361 bl[361] br[361] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_362 bl[362] br[362] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_363 bl[363] br[363] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_364 bl[364] br[364] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_365 bl[365] br[365] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_366 bl[366] br[366] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_367 bl[367] br[367] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_368 bl[368] br[368] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_369 bl[369] br[369] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_370 bl[370] br[370] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_371 bl[371] br[371] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_372 bl[372] br[372] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_373 bl[373] br[373] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_374 bl[374] br[374] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_375 bl[375] br[375] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_376 bl[376] br[376] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_377 bl[377] br[377] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_378 bl[378] br[378] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_379 bl[379] br[379] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_380 bl[380] br[380] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_381 bl[381] br[381] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_382 bl[382] br[382] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_383 bl[383] br[383] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_384 bl[384] br[384] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_385 bl[385] br[385] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_386 bl[386] br[386] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_387 bl[387] br[387] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_388 bl[388] br[388] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_389 bl[389] br[389] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_390 bl[390] br[390] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_391 bl[391] br[391] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_392 bl[392] br[392] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_393 bl[393] br[393] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_394 bl[394] br[394] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_395 bl[395] br[395] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_396 bl[396] br[396] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_397 bl[397] br[397] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_398 bl[398] br[398] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_399 bl[399] br[399] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_400 bl[400] br[400] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_401 bl[401] br[401] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_402 bl[402] br[402] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_403 bl[403] br[403] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_404 bl[404] br[404] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_405 bl[405] br[405] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_406 bl[406] br[406] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_407 bl[407] br[407] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_408 bl[408] br[408] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_409 bl[409] br[409] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_410 bl[410] br[410] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_411 bl[411] br[411] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_412 bl[412] br[412] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_413 bl[413] br[413] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_414 bl[414] br[414] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_415 bl[415] br[415] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_416 bl[416] br[416] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_417 bl[417] br[417] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_418 bl[418] br[418] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_419 bl[419] br[419] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_420 bl[420] br[420] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_421 bl[421] br[421] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_422 bl[422] br[422] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_423 bl[423] br[423] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_424 bl[424] br[424] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_425 bl[425] br[425] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_426 bl[426] br[426] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_427 bl[427] br[427] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_428 bl[428] br[428] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_429 bl[429] br[429] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_430 bl[430] br[430] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_431 bl[431] br[431] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_432 bl[432] br[432] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_433 bl[433] br[433] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_434 bl[434] br[434] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_435 bl[435] br[435] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_436 bl[436] br[436] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_437 bl[437] br[437] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_438 bl[438] br[438] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_439 bl[439] br[439] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_440 bl[440] br[440] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_441 bl[441] br[441] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_442 bl[442] br[442] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_443 bl[443] br[443] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_444 bl[444] br[444] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_445 bl[445] br[445] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_446 bl[446] br[446] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_447 bl[447] br[447] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_448 bl[448] br[448] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_449 bl[449] br[449] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_450 bl[450] br[450] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_451 bl[451] br[451] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_452 bl[452] br[452] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_453 bl[453] br[453] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_454 bl[454] br[454] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_455 bl[455] br[455] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_456 bl[456] br[456] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_457 bl[457] br[457] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_458 bl[458] br[458] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_459 bl[459] br[459] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_460 bl[460] br[460] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_461 bl[461] br[461] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_462 bl[462] br[462] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_463 bl[463] br[463] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_464 bl[464] br[464] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_465 bl[465] br[465] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_466 bl[466] br[466] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_467 bl[467] br[467] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_468 bl[468] br[468] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_469 bl[469] br[469] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_470 bl[470] br[470] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_471 bl[471] br[471] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_472 bl[472] br[472] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_473 bl[473] br[473] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_474 bl[474] br[474] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_475 bl[475] br[475] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_476 bl[476] br[476] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_477 bl[477] br[477] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_478 bl[478] br[478] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_479 bl[479] br[479] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_480 bl[480] br[480] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_481 bl[481] br[481] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_482 bl[482] br[482] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_483 bl[483] br[483] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_484 bl[484] br[484] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_485 bl[485] br[485] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_486 bl[486] br[486] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_487 bl[487] br[487] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_488 bl[488] br[488] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_489 bl[489] br[489] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_490 bl[490] br[490] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_491 bl[491] br[491] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_492 bl[492] br[492] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_493 bl[493] br[493] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_494 bl[494] br[494] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_495 bl[495] br[495] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_496 bl[496] br[496] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_497 bl[497] br[497] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_498 bl[498] br[498] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_499 bl[499] br[499] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_500 bl[500] br[500] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_501 bl[501] br[501] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_502 bl[502] br[502] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_503 bl[503] br[503] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_504 bl[504] br[504] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_505 bl[505] br[505] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_506 bl[506] br[506] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_507 bl[507] br[507] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_508 bl[508] br[508] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_509 bl[509] br[509] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_510 bl[510] br[510] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_61_511 bl[511] br[511] vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xcell_62_0 bl[0] br[0] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_1 bl[1] br[1] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_2 bl[2] br[2] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_3 bl[3] br[3] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_4 bl[4] br[4] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_5 bl[5] br[5] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_6 bl[6] br[6] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_7 bl[7] br[7] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_8 bl[8] br[8] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_9 bl[9] br[9] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_10 bl[10] br[10] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_11 bl[11] br[11] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_12 bl[12] br[12] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_13 bl[13] br[13] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_14 bl[14] br[14] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_15 bl[15] br[15] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_16 bl[16] br[16] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_17 bl[17] br[17] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_18 bl[18] br[18] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_19 bl[19] br[19] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_20 bl[20] br[20] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_21 bl[21] br[21] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_22 bl[22] br[22] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_23 bl[23] br[23] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_24 bl[24] br[24] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_25 bl[25] br[25] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_26 bl[26] br[26] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_27 bl[27] br[27] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_28 bl[28] br[28] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_29 bl[29] br[29] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_30 bl[30] br[30] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_31 bl[31] br[31] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_32 bl[32] br[32] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_33 bl[33] br[33] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_34 bl[34] br[34] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_35 bl[35] br[35] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_36 bl[36] br[36] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_37 bl[37] br[37] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_38 bl[38] br[38] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_39 bl[39] br[39] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_40 bl[40] br[40] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_41 bl[41] br[41] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_42 bl[42] br[42] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_43 bl[43] br[43] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_44 bl[44] br[44] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_45 bl[45] br[45] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_46 bl[46] br[46] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_47 bl[47] br[47] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_48 bl[48] br[48] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_49 bl[49] br[49] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_50 bl[50] br[50] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_51 bl[51] br[51] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_52 bl[52] br[52] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_53 bl[53] br[53] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_54 bl[54] br[54] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_55 bl[55] br[55] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_56 bl[56] br[56] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_57 bl[57] br[57] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_58 bl[58] br[58] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_59 bl[59] br[59] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_60 bl[60] br[60] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_61 bl[61] br[61] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_62 bl[62] br[62] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_63 bl[63] br[63] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_64 bl[64] br[64] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_65 bl[65] br[65] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_66 bl[66] br[66] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_67 bl[67] br[67] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_68 bl[68] br[68] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_69 bl[69] br[69] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_70 bl[70] br[70] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_71 bl[71] br[71] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_72 bl[72] br[72] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_73 bl[73] br[73] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_74 bl[74] br[74] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_75 bl[75] br[75] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_76 bl[76] br[76] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_77 bl[77] br[77] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_78 bl[78] br[78] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_79 bl[79] br[79] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_80 bl[80] br[80] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_81 bl[81] br[81] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_82 bl[82] br[82] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_83 bl[83] br[83] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_84 bl[84] br[84] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_85 bl[85] br[85] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_86 bl[86] br[86] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_87 bl[87] br[87] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_88 bl[88] br[88] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_89 bl[89] br[89] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_90 bl[90] br[90] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_91 bl[91] br[91] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_92 bl[92] br[92] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_93 bl[93] br[93] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_94 bl[94] br[94] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_95 bl[95] br[95] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_96 bl[96] br[96] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_97 bl[97] br[97] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_98 bl[98] br[98] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_99 bl[99] br[99] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_100 bl[100] br[100] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_101 bl[101] br[101] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_102 bl[102] br[102] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_103 bl[103] br[103] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_104 bl[104] br[104] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_105 bl[105] br[105] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_106 bl[106] br[106] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_107 bl[107] br[107] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_108 bl[108] br[108] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_109 bl[109] br[109] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_110 bl[110] br[110] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_111 bl[111] br[111] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_112 bl[112] br[112] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_113 bl[113] br[113] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_114 bl[114] br[114] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_115 bl[115] br[115] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_116 bl[116] br[116] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_117 bl[117] br[117] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_118 bl[118] br[118] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_119 bl[119] br[119] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_120 bl[120] br[120] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_121 bl[121] br[121] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_122 bl[122] br[122] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_123 bl[123] br[123] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_124 bl[124] br[124] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_125 bl[125] br[125] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_126 bl[126] br[126] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_127 bl[127] br[127] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_128 bl[128] br[128] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_129 bl[129] br[129] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_130 bl[130] br[130] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_131 bl[131] br[131] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_132 bl[132] br[132] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_133 bl[133] br[133] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_134 bl[134] br[134] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_135 bl[135] br[135] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_136 bl[136] br[136] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_137 bl[137] br[137] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_138 bl[138] br[138] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_139 bl[139] br[139] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_140 bl[140] br[140] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_141 bl[141] br[141] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_142 bl[142] br[142] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_143 bl[143] br[143] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_144 bl[144] br[144] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_145 bl[145] br[145] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_146 bl[146] br[146] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_147 bl[147] br[147] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_148 bl[148] br[148] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_149 bl[149] br[149] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_150 bl[150] br[150] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_151 bl[151] br[151] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_152 bl[152] br[152] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_153 bl[153] br[153] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_154 bl[154] br[154] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_155 bl[155] br[155] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_156 bl[156] br[156] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_157 bl[157] br[157] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_158 bl[158] br[158] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_159 bl[159] br[159] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_160 bl[160] br[160] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_161 bl[161] br[161] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_162 bl[162] br[162] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_163 bl[163] br[163] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_164 bl[164] br[164] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_165 bl[165] br[165] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_166 bl[166] br[166] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_167 bl[167] br[167] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_168 bl[168] br[168] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_169 bl[169] br[169] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_170 bl[170] br[170] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_171 bl[171] br[171] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_172 bl[172] br[172] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_173 bl[173] br[173] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_174 bl[174] br[174] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_175 bl[175] br[175] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_176 bl[176] br[176] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_177 bl[177] br[177] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_178 bl[178] br[178] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_179 bl[179] br[179] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_180 bl[180] br[180] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_181 bl[181] br[181] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_182 bl[182] br[182] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_183 bl[183] br[183] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_184 bl[184] br[184] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_185 bl[185] br[185] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_186 bl[186] br[186] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_187 bl[187] br[187] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_188 bl[188] br[188] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_189 bl[189] br[189] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_190 bl[190] br[190] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_191 bl[191] br[191] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_192 bl[192] br[192] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_193 bl[193] br[193] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_194 bl[194] br[194] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_195 bl[195] br[195] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_196 bl[196] br[196] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_197 bl[197] br[197] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_198 bl[198] br[198] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_199 bl[199] br[199] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_200 bl[200] br[200] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_201 bl[201] br[201] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_202 bl[202] br[202] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_203 bl[203] br[203] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_204 bl[204] br[204] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_205 bl[205] br[205] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_206 bl[206] br[206] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_207 bl[207] br[207] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_208 bl[208] br[208] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_209 bl[209] br[209] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_210 bl[210] br[210] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_211 bl[211] br[211] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_212 bl[212] br[212] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_213 bl[213] br[213] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_214 bl[214] br[214] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_215 bl[215] br[215] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_216 bl[216] br[216] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_217 bl[217] br[217] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_218 bl[218] br[218] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_219 bl[219] br[219] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_220 bl[220] br[220] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_221 bl[221] br[221] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_222 bl[222] br[222] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_223 bl[223] br[223] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_224 bl[224] br[224] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_225 bl[225] br[225] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_226 bl[226] br[226] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_227 bl[227] br[227] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_228 bl[228] br[228] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_229 bl[229] br[229] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_230 bl[230] br[230] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_231 bl[231] br[231] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_232 bl[232] br[232] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_233 bl[233] br[233] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_234 bl[234] br[234] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_235 bl[235] br[235] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_236 bl[236] br[236] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_237 bl[237] br[237] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_238 bl[238] br[238] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_239 bl[239] br[239] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_240 bl[240] br[240] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_241 bl[241] br[241] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_242 bl[242] br[242] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_243 bl[243] br[243] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_244 bl[244] br[244] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_245 bl[245] br[245] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_246 bl[246] br[246] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_247 bl[247] br[247] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_248 bl[248] br[248] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_249 bl[249] br[249] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_250 bl[250] br[250] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_251 bl[251] br[251] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_252 bl[252] br[252] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_253 bl[253] br[253] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_254 bl[254] br[254] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_255 bl[255] br[255] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_256 bl[256] br[256] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_257 bl[257] br[257] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_258 bl[258] br[258] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_259 bl[259] br[259] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_260 bl[260] br[260] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_261 bl[261] br[261] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_262 bl[262] br[262] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_263 bl[263] br[263] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_264 bl[264] br[264] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_265 bl[265] br[265] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_266 bl[266] br[266] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_267 bl[267] br[267] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_268 bl[268] br[268] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_269 bl[269] br[269] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_270 bl[270] br[270] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_271 bl[271] br[271] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_272 bl[272] br[272] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_273 bl[273] br[273] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_274 bl[274] br[274] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_275 bl[275] br[275] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_276 bl[276] br[276] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_277 bl[277] br[277] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_278 bl[278] br[278] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_279 bl[279] br[279] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_280 bl[280] br[280] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_281 bl[281] br[281] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_282 bl[282] br[282] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_283 bl[283] br[283] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_284 bl[284] br[284] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_285 bl[285] br[285] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_286 bl[286] br[286] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_287 bl[287] br[287] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_288 bl[288] br[288] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_289 bl[289] br[289] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_290 bl[290] br[290] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_291 bl[291] br[291] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_292 bl[292] br[292] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_293 bl[293] br[293] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_294 bl[294] br[294] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_295 bl[295] br[295] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_296 bl[296] br[296] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_297 bl[297] br[297] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_298 bl[298] br[298] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_299 bl[299] br[299] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_300 bl[300] br[300] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_301 bl[301] br[301] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_302 bl[302] br[302] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_303 bl[303] br[303] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_304 bl[304] br[304] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_305 bl[305] br[305] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_306 bl[306] br[306] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_307 bl[307] br[307] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_308 bl[308] br[308] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_309 bl[309] br[309] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_310 bl[310] br[310] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_311 bl[311] br[311] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_312 bl[312] br[312] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_313 bl[313] br[313] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_314 bl[314] br[314] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_315 bl[315] br[315] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_316 bl[316] br[316] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_317 bl[317] br[317] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_318 bl[318] br[318] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_319 bl[319] br[319] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_320 bl[320] br[320] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_321 bl[321] br[321] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_322 bl[322] br[322] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_323 bl[323] br[323] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_324 bl[324] br[324] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_325 bl[325] br[325] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_326 bl[326] br[326] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_327 bl[327] br[327] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_328 bl[328] br[328] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_329 bl[329] br[329] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_330 bl[330] br[330] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_331 bl[331] br[331] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_332 bl[332] br[332] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_333 bl[333] br[333] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_334 bl[334] br[334] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_335 bl[335] br[335] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_336 bl[336] br[336] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_337 bl[337] br[337] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_338 bl[338] br[338] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_339 bl[339] br[339] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_340 bl[340] br[340] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_341 bl[341] br[341] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_342 bl[342] br[342] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_343 bl[343] br[343] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_344 bl[344] br[344] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_345 bl[345] br[345] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_346 bl[346] br[346] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_347 bl[347] br[347] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_348 bl[348] br[348] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_349 bl[349] br[349] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_350 bl[350] br[350] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_351 bl[351] br[351] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_352 bl[352] br[352] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_353 bl[353] br[353] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_354 bl[354] br[354] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_355 bl[355] br[355] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_356 bl[356] br[356] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_357 bl[357] br[357] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_358 bl[358] br[358] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_359 bl[359] br[359] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_360 bl[360] br[360] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_361 bl[361] br[361] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_362 bl[362] br[362] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_363 bl[363] br[363] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_364 bl[364] br[364] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_365 bl[365] br[365] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_366 bl[366] br[366] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_367 bl[367] br[367] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_368 bl[368] br[368] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_369 bl[369] br[369] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_370 bl[370] br[370] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_371 bl[371] br[371] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_372 bl[372] br[372] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_373 bl[373] br[373] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_374 bl[374] br[374] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_375 bl[375] br[375] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_376 bl[376] br[376] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_377 bl[377] br[377] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_378 bl[378] br[378] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_379 bl[379] br[379] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_380 bl[380] br[380] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_381 bl[381] br[381] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_382 bl[382] br[382] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_383 bl[383] br[383] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_384 bl[384] br[384] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_385 bl[385] br[385] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_386 bl[386] br[386] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_387 bl[387] br[387] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_388 bl[388] br[388] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_389 bl[389] br[389] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_390 bl[390] br[390] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_391 bl[391] br[391] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_392 bl[392] br[392] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_393 bl[393] br[393] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_394 bl[394] br[394] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_395 bl[395] br[395] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_396 bl[396] br[396] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_397 bl[397] br[397] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_398 bl[398] br[398] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_399 bl[399] br[399] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_400 bl[400] br[400] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_401 bl[401] br[401] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_402 bl[402] br[402] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_403 bl[403] br[403] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_404 bl[404] br[404] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_405 bl[405] br[405] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_406 bl[406] br[406] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_407 bl[407] br[407] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_408 bl[408] br[408] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_409 bl[409] br[409] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_410 bl[410] br[410] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_411 bl[411] br[411] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_412 bl[412] br[412] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_413 bl[413] br[413] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_414 bl[414] br[414] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_415 bl[415] br[415] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_416 bl[416] br[416] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_417 bl[417] br[417] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_418 bl[418] br[418] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_419 bl[419] br[419] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_420 bl[420] br[420] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_421 bl[421] br[421] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_422 bl[422] br[422] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_423 bl[423] br[423] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_424 bl[424] br[424] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_425 bl[425] br[425] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_426 bl[426] br[426] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_427 bl[427] br[427] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_428 bl[428] br[428] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_429 bl[429] br[429] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_430 bl[430] br[430] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_431 bl[431] br[431] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_432 bl[432] br[432] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_433 bl[433] br[433] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_434 bl[434] br[434] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_435 bl[435] br[435] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_436 bl[436] br[436] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_437 bl[437] br[437] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_438 bl[438] br[438] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_439 bl[439] br[439] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_440 bl[440] br[440] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_441 bl[441] br[441] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_442 bl[442] br[442] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_443 bl[443] br[443] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_444 bl[444] br[444] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_445 bl[445] br[445] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_446 bl[446] br[446] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_447 bl[447] br[447] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_448 bl[448] br[448] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_449 bl[449] br[449] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_450 bl[450] br[450] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_451 bl[451] br[451] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_452 bl[452] br[452] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_453 bl[453] br[453] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_454 bl[454] br[454] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_455 bl[455] br[455] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_456 bl[456] br[456] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_457 bl[457] br[457] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_458 bl[458] br[458] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_459 bl[459] br[459] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_460 bl[460] br[460] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_461 bl[461] br[461] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_462 bl[462] br[462] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_463 bl[463] br[463] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_464 bl[464] br[464] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_465 bl[465] br[465] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_466 bl[466] br[466] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_467 bl[467] br[467] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_468 bl[468] br[468] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_469 bl[469] br[469] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_470 bl[470] br[470] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_471 bl[471] br[471] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_472 bl[472] br[472] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_473 bl[473] br[473] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_474 bl[474] br[474] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_475 bl[475] br[475] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_476 bl[476] br[476] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_477 bl[477] br[477] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_478 bl[478] br[478] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_479 bl[479] br[479] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_480 bl[480] br[480] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_481 bl[481] br[481] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_482 bl[482] br[482] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_483 bl[483] br[483] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_484 bl[484] br[484] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_485 bl[485] br[485] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_486 bl[486] br[486] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_487 bl[487] br[487] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_488 bl[488] br[488] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_489 bl[489] br[489] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_490 bl[490] br[490] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_491 bl[491] br[491] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_492 bl[492] br[492] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_493 bl[493] br[493] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_494 bl[494] br[494] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_495 bl[495] br[495] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_496 bl[496] br[496] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_497 bl[497] br[497] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_498 bl[498] br[498] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_499 bl[499] br[499] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_500 bl[500] br[500] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_501 bl[501] br[501] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_502 bl[502] br[502] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_503 bl[503] br[503] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_504 bl[504] br[504] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_505 bl[505] br[505] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_506 bl[506] br[506] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_507 bl[507] br[507] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_508 bl[508] br[508] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_509 bl[509] br[509] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_510 bl[510] br[510] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_62_511 bl[511] br[511] vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xcell_63_0 bl[0] br[0] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_1 bl[1] br[1] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_2 bl[2] br[2] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_3 bl[3] br[3] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_4 bl[4] br[4] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_5 bl[5] br[5] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_6 bl[6] br[6] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_7 bl[7] br[7] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_8 bl[8] br[8] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_9 bl[9] br[9] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_10 bl[10] br[10] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_11 bl[11] br[11] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_12 bl[12] br[12] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_13 bl[13] br[13] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_14 bl[14] br[14] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_15 bl[15] br[15] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_16 bl[16] br[16] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_17 bl[17] br[17] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_18 bl[18] br[18] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_19 bl[19] br[19] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_20 bl[20] br[20] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_21 bl[21] br[21] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_22 bl[22] br[22] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_23 bl[23] br[23] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_24 bl[24] br[24] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_25 bl[25] br[25] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_26 bl[26] br[26] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_27 bl[27] br[27] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_28 bl[28] br[28] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_29 bl[29] br[29] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_30 bl[30] br[30] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_31 bl[31] br[31] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_32 bl[32] br[32] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_33 bl[33] br[33] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_34 bl[34] br[34] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_35 bl[35] br[35] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_36 bl[36] br[36] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_37 bl[37] br[37] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_38 bl[38] br[38] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_39 bl[39] br[39] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_40 bl[40] br[40] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_41 bl[41] br[41] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_42 bl[42] br[42] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_43 bl[43] br[43] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_44 bl[44] br[44] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_45 bl[45] br[45] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_46 bl[46] br[46] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_47 bl[47] br[47] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_48 bl[48] br[48] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_49 bl[49] br[49] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_50 bl[50] br[50] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_51 bl[51] br[51] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_52 bl[52] br[52] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_53 bl[53] br[53] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_54 bl[54] br[54] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_55 bl[55] br[55] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_56 bl[56] br[56] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_57 bl[57] br[57] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_58 bl[58] br[58] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_59 bl[59] br[59] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_60 bl[60] br[60] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_61 bl[61] br[61] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_62 bl[62] br[62] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_63 bl[63] br[63] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_64 bl[64] br[64] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_65 bl[65] br[65] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_66 bl[66] br[66] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_67 bl[67] br[67] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_68 bl[68] br[68] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_69 bl[69] br[69] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_70 bl[70] br[70] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_71 bl[71] br[71] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_72 bl[72] br[72] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_73 bl[73] br[73] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_74 bl[74] br[74] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_75 bl[75] br[75] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_76 bl[76] br[76] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_77 bl[77] br[77] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_78 bl[78] br[78] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_79 bl[79] br[79] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_80 bl[80] br[80] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_81 bl[81] br[81] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_82 bl[82] br[82] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_83 bl[83] br[83] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_84 bl[84] br[84] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_85 bl[85] br[85] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_86 bl[86] br[86] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_87 bl[87] br[87] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_88 bl[88] br[88] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_89 bl[89] br[89] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_90 bl[90] br[90] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_91 bl[91] br[91] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_92 bl[92] br[92] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_93 bl[93] br[93] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_94 bl[94] br[94] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_95 bl[95] br[95] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_96 bl[96] br[96] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_97 bl[97] br[97] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_98 bl[98] br[98] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_99 bl[99] br[99] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_100 bl[100] br[100] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_101 bl[101] br[101] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_102 bl[102] br[102] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_103 bl[103] br[103] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_104 bl[104] br[104] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_105 bl[105] br[105] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_106 bl[106] br[106] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_107 bl[107] br[107] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_108 bl[108] br[108] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_109 bl[109] br[109] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_110 bl[110] br[110] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_111 bl[111] br[111] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_112 bl[112] br[112] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_113 bl[113] br[113] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_114 bl[114] br[114] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_115 bl[115] br[115] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_116 bl[116] br[116] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_117 bl[117] br[117] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_118 bl[118] br[118] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_119 bl[119] br[119] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_120 bl[120] br[120] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_121 bl[121] br[121] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_122 bl[122] br[122] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_123 bl[123] br[123] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_124 bl[124] br[124] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_125 bl[125] br[125] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_126 bl[126] br[126] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_127 bl[127] br[127] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_128 bl[128] br[128] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_129 bl[129] br[129] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_130 bl[130] br[130] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_131 bl[131] br[131] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_132 bl[132] br[132] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_133 bl[133] br[133] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_134 bl[134] br[134] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_135 bl[135] br[135] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_136 bl[136] br[136] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_137 bl[137] br[137] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_138 bl[138] br[138] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_139 bl[139] br[139] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_140 bl[140] br[140] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_141 bl[141] br[141] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_142 bl[142] br[142] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_143 bl[143] br[143] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_144 bl[144] br[144] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_145 bl[145] br[145] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_146 bl[146] br[146] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_147 bl[147] br[147] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_148 bl[148] br[148] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_149 bl[149] br[149] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_150 bl[150] br[150] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_151 bl[151] br[151] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_152 bl[152] br[152] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_153 bl[153] br[153] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_154 bl[154] br[154] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_155 bl[155] br[155] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_156 bl[156] br[156] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_157 bl[157] br[157] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_158 bl[158] br[158] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_159 bl[159] br[159] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_160 bl[160] br[160] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_161 bl[161] br[161] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_162 bl[162] br[162] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_163 bl[163] br[163] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_164 bl[164] br[164] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_165 bl[165] br[165] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_166 bl[166] br[166] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_167 bl[167] br[167] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_168 bl[168] br[168] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_169 bl[169] br[169] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_170 bl[170] br[170] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_171 bl[171] br[171] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_172 bl[172] br[172] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_173 bl[173] br[173] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_174 bl[174] br[174] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_175 bl[175] br[175] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_176 bl[176] br[176] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_177 bl[177] br[177] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_178 bl[178] br[178] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_179 bl[179] br[179] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_180 bl[180] br[180] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_181 bl[181] br[181] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_182 bl[182] br[182] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_183 bl[183] br[183] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_184 bl[184] br[184] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_185 bl[185] br[185] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_186 bl[186] br[186] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_187 bl[187] br[187] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_188 bl[188] br[188] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_189 bl[189] br[189] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_190 bl[190] br[190] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_191 bl[191] br[191] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_192 bl[192] br[192] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_193 bl[193] br[193] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_194 bl[194] br[194] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_195 bl[195] br[195] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_196 bl[196] br[196] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_197 bl[197] br[197] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_198 bl[198] br[198] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_199 bl[199] br[199] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_200 bl[200] br[200] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_201 bl[201] br[201] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_202 bl[202] br[202] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_203 bl[203] br[203] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_204 bl[204] br[204] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_205 bl[205] br[205] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_206 bl[206] br[206] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_207 bl[207] br[207] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_208 bl[208] br[208] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_209 bl[209] br[209] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_210 bl[210] br[210] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_211 bl[211] br[211] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_212 bl[212] br[212] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_213 bl[213] br[213] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_214 bl[214] br[214] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_215 bl[215] br[215] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_216 bl[216] br[216] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_217 bl[217] br[217] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_218 bl[218] br[218] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_219 bl[219] br[219] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_220 bl[220] br[220] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_221 bl[221] br[221] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_222 bl[222] br[222] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_223 bl[223] br[223] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_224 bl[224] br[224] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_225 bl[225] br[225] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_226 bl[226] br[226] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_227 bl[227] br[227] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_228 bl[228] br[228] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_229 bl[229] br[229] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_230 bl[230] br[230] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_231 bl[231] br[231] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_232 bl[232] br[232] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_233 bl[233] br[233] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_234 bl[234] br[234] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_235 bl[235] br[235] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_236 bl[236] br[236] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_237 bl[237] br[237] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_238 bl[238] br[238] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_239 bl[239] br[239] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_240 bl[240] br[240] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_241 bl[241] br[241] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_242 bl[242] br[242] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_243 bl[243] br[243] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_244 bl[244] br[244] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_245 bl[245] br[245] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_246 bl[246] br[246] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_247 bl[247] br[247] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_248 bl[248] br[248] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_249 bl[249] br[249] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_250 bl[250] br[250] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_251 bl[251] br[251] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_252 bl[252] br[252] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_253 bl[253] br[253] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_254 bl[254] br[254] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_255 bl[255] br[255] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_256 bl[256] br[256] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_257 bl[257] br[257] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_258 bl[258] br[258] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_259 bl[259] br[259] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_260 bl[260] br[260] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_261 bl[261] br[261] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_262 bl[262] br[262] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_263 bl[263] br[263] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_264 bl[264] br[264] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_265 bl[265] br[265] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_266 bl[266] br[266] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_267 bl[267] br[267] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_268 bl[268] br[268] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_269 bl[269] br[269] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_270 bl[270] br[270] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_271 bl[271] br[271] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_272 bl[272] br[272] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_273 bl[273] br[273] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_274 bl[274] br[274] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_275 bl[275] br[275] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_276 bl[276] br[276] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_277 bl[277] br[277] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_278 bl[278] br[278] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_279 bl[279] br[279] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_280 bl[280] br[280] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_281 bl[281] br[281] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_282 bl[282] br[282] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_283 bl[283] br[283] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_284 bl[284] br[284] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_285 bl[285] br[285] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_286 bl[286] br[286] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_287 bl[287] br[287] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_288 bl[288] br[288] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_289 bl[289] br[289] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_290 bl[290] br[290] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_291 bl[291] br[291] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_292 bl[292] br[292] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_293 bl[293] br[293] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_294 bl[294] br[294] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_295 bl[295] br[295] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_296 bl[296] br[296] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_297 bl[297] br[297] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_298 bl[298] br[298] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_299 bl[299] br[299] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_300 bl[300] br[300] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_301 bl[301] br[301] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_302 bl[302] br[302] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_303 bl[303] br[303] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_304 bl[304] br[304] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_305 bl[305] br[305] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_306 bl[306] br[306] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_307 bl[307] br[307] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_308 bl[308] br[308] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_309 bl[309] br[309] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_310 bl[310] br[310] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_311 bl[311] br[311] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_312 bl[312] br[312] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_313 bl[313] br[313] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_314 bl[314] br[314] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_315 bl[315] br[315] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_316 bl[316] br[316] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_317 bl[317] br[317] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_318 bl[318] br[318] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_319 bl[319] br[319] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_320 bl[320] br[320] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_321 bl[321] br[321] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_322 bl[322] br[322] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_323 bl[323] br[323] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_324 bl[324] br[324] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_325 bl[325] br[325] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_326 bl[326] br[326] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_327 bl[327] br[327] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_328 bl[328] br[328] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_329 bl[329] br[329] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_330 bl[330] br[330] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_331 bl[331] br[331] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_332 bl[332] br[332] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_333 bl[333] br[333] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_334 bl[334] br[334] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_335 bl[335] br[335] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_336 bl[336] br[336] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_337 bl[337] br[337] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_338 bl[338] br[338] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_339 bl[339] br[339] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_340 bl[340] br[340] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_341 bl[341] br[341] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_342 bl[342] br[342] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_343 bl[343] br[343] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_344 bl[344] br[344] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_345 bl[345] br[345] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_346 bl[346] br[346] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_347 bl[347] br[347] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_348 bl[348] br[348] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_349 bl[349] br[349] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_350 bl[350] br[350] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_351 bl[351] br[351] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_352 bl[352] br[352] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_353 bl[353] br[353] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_354 bl[354] br[354] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_355 bl[355] br[355] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_356 bl[356] br[356] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_357 bl[357] br[357] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_358 bl[358] br[358] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_359 bl[359] br[359] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_360 bl[360] br[360] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_361 bl[361] br[361] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_362 bl[362] br[362] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_363 bl[363] br[363] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_364 bl[364] br[364] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_365 bl[365] br[365] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_366 bl[366] br[366] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_367 bl[367] br[367] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_368 bl[368] br[368] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_369 bl[369] br[369] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_370 bl[370] br[370] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_371 bl[371] br[371] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_372 bl[372] br[372] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_373 bl[373] br[373] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_374 bl[374] br[374] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_375 bl[375] br[375] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_376 bl[376] br[376] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_377 bl[377] br[377] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_378 bl[378] br[378] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_379 bl[379] br[379] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_380 bl[380] br[380] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_381 bl[381] br[381] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_382 bl[382] br[382] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_383 bl[383] br[383] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_384 bl[384] br[384] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_385 bl[385] br[385] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_386 bl[386] br[386] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_387 bl[387] br[387] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_388 bl[388] br[388] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_389 bl[389] br[389] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_390 bl[390] br[390] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_391 bl[391] br[391] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_392 bl[392] br[392] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_393 bl[393] br[393] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_394 bl[394] br[394] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_395 bl[395] br[395] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_396 bl[396] br[396] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_397 bl[397] br[397] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_398 bl[398] br[398] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_399 bl[399] br[399] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_400 bl[400] br[400] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_401 bl[401] br[401] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_402 bl[402] br[402] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_403 bl[403] br[403] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_404 bl[404] br[404] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_405 bl[405] br[405] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_406 bl[406] br[406] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_407 bl[407] br[407] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_408 bl[408] br[408] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_409 bl[409] br[409] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_410 bl[410] br[410] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_411 bl[411] br[411] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_412 bl[412] br[412] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_413 bl[413] br[413] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_414 bl[414] br[414] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_415 bl[415] br[415] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_416 bl[416] br[416] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_417 bl[417] br[417] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_418 bl[418] br[418] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_419 bl[419] br[419] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_420 bl[420] br[420] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_421 bl[421] br[421] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_422 bl[422] br[422] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_423 bl[423] br[423] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_424 bl[424] br[424] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_425 bl[425] br[425] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_426 bl[426] br[426] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_427 bl[427] br[427] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_428 bl[428] br[428] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_429 bl[429] br[429] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_430 bl[430] br[430] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_431 bl[431] br[431] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_432 bl[432] br[432] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_433 bl[433] br[433] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_434 bl[434] br[434] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_435 bl[435] br[435] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_436 bl[436] br[436] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_437 bl[437] br[437] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_438 bl[438] br[438] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_439 bl[439] br[439] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_440 bl[440] br[440] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_441 bl[441] br[441] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_442 bl[442] br[442] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_443 bl[443] br[443] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_444 bl[444] br[444] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_445 bl[445] br[445] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_446 bl[446] br[446] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_447 bl[447] br[447] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_448 bl[448] br[448] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_449 bl[449] br[449] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_450 bl[450] br[450] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_451 bl[451] br[451] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_452 bl[452] br[452] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_453 bl[453] br[453] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_454 bl[454] br[454] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_455 bl[455] br[455] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_456 bl[456] br[456] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_457 bl[457] br[457] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_458 bl[458] br[458] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_459 bl[459] br[459] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_460 bl[460] br[460] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_461 bl[461] br[461] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_462 bl[462] br[462] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_463 bl[463] br[463] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_464 bl[464] br[464] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_465 bl[465] br[465] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_466 bl[466] br[466] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_467 bl[467] br[467] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_468 bl[468] br[468] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_469 bl[469] br[469] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_470 bl[470] br[470] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_471 bl[471] br[471] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_472 bl[472] br[472] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_473 bl[473] br[473] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_474 bl[474] br[474] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_475 bl[475] br[475] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_476 bl[476] br[476] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_477 bl[477] br[477] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_478 bl[478] br[478] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_479 bl[479] br[479] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_480 bl[480] br[480] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_481 bl[481] br[481] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_482 bl[482] br[482] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_483 bl[483] br[483] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_484 bl[484] br[484] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_485 bl[485] br[485] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_486 bl[486] br[486] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_487 bl[487] br[487] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_488 bl[488] br[488] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_489 bl[489] br[489] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_490 bl[490] br[490] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_491 bl[491] br[491] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_492 bl[492] br[492] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_493 bl[493] br[493] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_494 bl[494] br[494] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_495 bl[495] br[495] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_496 bl[496] br[496] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_497 bl[497] br[497] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_498 bl[498] br[498] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_499 bl[499] br[499] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_500 bl[500] br[500] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_501 bl[501] br[501] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_502 bl[502] br[502] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_503 bl[503] br[503] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_504 bl[504] br[504] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_505 bl[505] br[505] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_506 bl[506] br[506] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_507 bl[507] br[507] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_508 bl[508] br[508] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_509 bl[509] br[509] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_510 bl[510] br[510] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xcell_63_511 bl[511] br[511] vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_0 dummy_bl dummy_br vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_0 vdd vdd vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_1 dummy_bl dummy_br vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_1 vdd vdd vdd vss wl[0] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_2 dummy_bl dummy_br vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_2 vdd vdd vdd vss wl[1] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_3 dummy_bl dummy_br vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_3 vdd vdd vdd vss wl[2] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_4 dummy_bl dummy_br vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_4 vdd vdd vdd vss wl[3] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_5 dummy_bl dummy_br vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_5 vdd vdd vdd vss wl[4] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_6 dummy_bl dummy_br vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_6 vdd vdd vdd vss wl[5] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_7 dummy_bl dummy_br vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_7 vdd vdd vdd vss wl[6] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_8 dummy_bl dummy_br vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_8 vdd vdd vdd vss wl[7] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_9 dummy_bl dummy_br vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_9 vdd vdd vdd vss wl[8] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_10 dummy_bl dummy_br vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_10 vdd vdd vdd vss wl[9] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_11 dummy_bl dummy_br vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_11 vdd vdd vdd vss wl[10] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_12 dummy_bl dummy_br vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_12 vdd vdd vdd vss wl[11] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_13 dummy_bl dummy_br vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_13 vdd vdd vdd vss wl[12] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_14 dummy_bl dummy_br vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_14 vdd vdd vdd vss wl[13] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_15 dummy_bl dummy_br vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_15 vdd vdd vdd vss wl[14] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_16 dummy_bl dummy_br vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_16 vdd vdd vdd vss wl[15] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_17 dummy_bl dummy_br vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_17 vdd vdd vdd vss wl[16] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_18 dummy_bl dummy_br vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_18 vdd vdd vdd vss wl[17] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_19 dummy_bl dummy_br vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_19 vdd vdd vdd vss wl[18] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_20 dummy_bl dummy_br vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_20 vdd vdd vdd vss wl[19] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_21 dummy_bl dummy_br vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_21 vdd vdd vdd vss wl[20] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_22 dummy_bl dummy_br vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_22 vdd vdd vdd vss wl[21] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_23 dummy_bl dummy_br vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_23 vdd vdd vdd vss wl[22] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_24 dummy_bl dummy_br vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_24 vdd vdd vdd vss wl[23] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_25 dummy_bl dummy_br vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_25 vdd vdd vdd vss wl[24] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_26 dummy_bl dummy_br vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_26 vdd vdd vdd vss wl[25] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_27 dummy_bl dummy_br vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_27 vdd vdd vdd vss wl[26] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_28 dummy_bl dummy_br vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_28 vdd vdd vdd vss wl[27] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_29 dummy_bl dummy_br vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_29 vdd vdd vdd vss wl[28] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_30 dummy_bl dummy_br vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_30 vdd vdd vdd vss wl[29] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_31 dummy_bl dummy_br vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_31 vdd vdd vdd vss wl[30] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_32 dummy_bl dummy_br vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_32 vdd vdd vdd vss wl[31] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_33 dummy_bl dummy_br vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_33 vdd vdd vdd vss wl[32] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_34 dummy_bl dummy_br vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_34 vdd vdd vdd vss wl[33] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_35 dummy_bl dummy_br vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_35 vdd vdd vdd vss wl[34] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_36 dummy_bl dummy_br vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_36 vdd vdd vdd vss wl[35] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_37 dummy_bl dummy_br vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_37 vdd vdd vdd vss wl[36] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_38 dummy_bl dummy_br vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_38 vdd vdd vdd vss wl[37] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_39 dummy_bl dummy_br vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_39 vdd vdd vdd vss wl[38] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_40 dummy_bl dummy_br vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_40 vdd vdd vdd vss wl[39] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_41 dummy_bl dummy_br vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_41 vdd vdd vdd vss wl[40] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_42 dummy_bl dummy_br vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_42 vdd vdd vdd vss wl[41] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_43 dummy_bl dummy_br vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_43 vdd vdd vdd vss wl[42] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_44 dummy_bl dummy_br vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_44 vdd vdd vdd vss wl[43] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_45 dummy_bl dummy_br vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_45 vdd vdd vdd vss wl[44] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_46 dummy_bl dummy_br vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_46 vdd vdd vdd vss wl[45] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_47 dummy_bl dummy_br vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_47 vdd vdd vdd vss wl[46] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_48 dummy_bl dummy_br vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_48 vdd vdd vdd vss wl[47] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_49 dummy_bl dummy_br vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_49 vdd vdd vdd vss wl[48] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_50 dummy_bl dummy_br vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_50 vdd vdd vdd vss wl[49] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_51 dummy_bl dummy_br vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_51 vdd vdd vdd vss wl[50] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_52 dummy_bl dummy_br vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_52 vdd vdd vdd vss wl[51] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_53 dummy_bl dummy_br vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_53 vdd vdd vdd vss wl[52] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_54 dummy_bl dummy_br vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_54 vdd vdd vdd vss wl[53] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_55 dummy_bl dummy_br vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_55 vdd vdd vdd vss wl[54] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_56 dummy_bl dummy_br vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_56 vdd vdd vdd vss wl[55] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_57 dummy_bl dummy_br vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_57 vdd vdd vdd vss wl[56] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_58 dummy_bl dummy_br vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_58 vdd vdd vdd vss wl[57] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_59 dummy_bl dummy_br vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_59 vdd vdd vdd vss wl[58] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_60 dummy_bl dummy_br vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_60 vdd vdd vdd vss wl[59] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_61 dummy_bl dummy_br vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_61 vdd vdd vdd vss wl[60] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_62 dummy_bl dummy_br vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_62 vdd vdd vdd vss wl[61] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_63 dummy_bl dummy_br vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_63 vdd vdd vdd vss wl[62] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_64 dummy_bl dummy_br vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_64 vdd vdd vdd vss wl[63] vss vdd sram_sp_cell_wrapper
  Xdummy_col_left_65 dummy_bl dummy_br vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_col_right_65 vdd vdd vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_0 bl[0] br[0] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_0 bl[0] br[0] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_1 bl[1] br[1] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_1 bl[1] br[1] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_2 bl[2] br[2] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_2 bl[2] br[2] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_3 bl[3] br[3] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_3 bl[3] br[3] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_4 bl[4] br[4] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_4 bl[4] br[4] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_5 bl[5] br[5] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_5 bl[5] br[5] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_6 bl[6] br[6] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_6 bl[6] br[6] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_7 bl[7] br[7] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_7 bl[7] br[7] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_8 bl[8] br[8] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_8 bl[8] br[8] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_9 bl[9] br[9] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_9 bl[9] br[9] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_10 bl[10] br[10] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_10 bl[10] br[10] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_11 bl[11] br[11] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_11 bl[11] br[11] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_12 bl[12] br[12] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_12 bl[12] br[12] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_13 bl[13] br[13] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_13 bl[13] br[13] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_14 bl[14] br[14] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_14 bl[14] br[14] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_15 bl[15] br[15] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_15 bl[15] br[15] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_16 bl[16] br[16] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_16 bl[16] br[16] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_17 bl[17] br[17] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_17 bl[17] br[17] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_18 bl[18] br[18] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_18 bl[18] br[18] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_19 bl[19] br[19] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_19 bl[19] br[19] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_20 bl[20] br[20] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_20 bl[20] br[20] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_21 bl[21] br[21] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_21 bl[21] br[21] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_22 bl[22] br[22] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_22 bl[22] br[22] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_23 bl[23] br[23] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_23 bl[23] br[23] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_24 bl[24] br[24] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_24 bl[24] br[24] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_25 bl[25] br[25] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_25 bl[25] br[25] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_26 bl[26] br[26] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_26 bl[26] br[26] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_27 bl[27] br[27] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_27 bl[27] br[27] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_28 bl[28] br[28] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_28 bl[28] br[28] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_29 bl[29] br[29] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_29 bl[29] br[29] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_30 bl[30] br[30] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_30 bl[30] br[30] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_31 bl[31] br[31] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_31 bl[31] br[31] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_32 bl[32] br[32] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_32 bl[32] br[32] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_33 bl[33] br[33] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_33 bl[33] br[33] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_34 bl[34] br[34] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_34 bl[34] br[34] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_35 bl[35] br[35] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_35 bl[35] br[35] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_36 bl[36] br[36] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_36 bl[36] br[36] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_37 bl[37] br[37] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_37 bl[37] br[37] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_38 bl[38] br[38] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_38 bl[38] br[38] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_39 bl[39] br[39] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_39 bl[39] br[39] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_40 bl[40] br[40] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_40 bl[40] br[40] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_41 bl[41] br[41] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_41 bl[41] br[41] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_42 bl[42] br[42] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_42 bl[42] br[42] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_43 bl[43] br[43] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_43 bl[43] br[43] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_44 bl[44] br[44] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_44 bl[44] br[44] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_45 bl[45] br[45] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_45 bl[45] br[45] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_46 bl[46] br[46] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_46 bl[46] br[46] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_47 bl[47] br[47] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_47 bl[47] br[47] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_48 bl[48] br[48] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_48 bl[48] br[48] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_49 bl[49] br[49] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_49 bl[49] br[49] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_50 bl[50] br[50] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_50 bl[50] br[50] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_51 bl[51] br[51] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_51 bl[51] br[51] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_52 bl[52] br[52] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_52 bl[52] br[52] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_53 bl[53] br[53] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_53 bl[53] br[53] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_54 bl[54] br[54] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_54 bl[54] br[54] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_55 bl[55] br[55] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_55 bl[55] br[55] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_56 bl[56] br[56] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_56 bl[56] br[56] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_57 bl[57] br[57] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_57 bl[57] br[57] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_58 bl[58] br[58] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_58 bl[58] br[58] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_59 bl[59] br[59] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_59 bl[59] br[59] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_60 bl[60] br[60] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_60 bl[60] br[60] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_61 bl[61] br[61] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_61 bl[61] br[61] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_62 bl[62] br[62] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_62 bl[62] br[62] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_63 bl[63] br[63] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_63 bl[63] br[63] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_64 bl[64] br[64] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_64 bl[64] br[64] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_65 bl[65] br[65] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_65 bl[65] br[65] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_66 bl[66] br[66] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_66 bl[66] br[66] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_67 bl[67] br[67] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_67 bl[67] br[67] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_68 bl[68] br[68] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_68 bl[68] br[68] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_69 bl[69] br[69] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_69 bl[69] br[69] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_70 bl[70] br[70] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_70 bl[70] br[70] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_71 bl[71] br[71] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_71 bl[71] br[71] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_72 bl[72] br[72] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_72 bl[72] br[72] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_73 bl[73] br[73] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_73 bl[73] br[73] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_74 bl[74] br[74] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_74 bl[74] br[74] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_75 bl[75] br[75] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_75 bl[75] br[75] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_76 bl[76] br[76] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_76 bl[76] br[76] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_77 bl[77] br[77] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_77 bl[77] br[77] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_78 bl[78] br[78] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_78 bl[78] br[78] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_79 bl[79] br[79] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_79 bl[79] br[79] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_80 bl[80] br[80] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_80 bl[80] br[80] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_81 bl[81] br[81] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_81 bl[81] br[81] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_82 bl[82] br[82] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_82 bl[82] br[82] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_83 bl[83] br[83] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_83 bl[83] br[83] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_84 bl[84] br[84] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_84 bl[84] br[84] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_85 bl[85] br[85] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_85 bl[85] br[85] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_86 bl[86] br[86] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_86 bl[86] br[86] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_87 bl[87] br[87] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_87 bl[87] br[87] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_88 bl[88] br[88] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_88 bl[88] br[88] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_89 bl[89] br[89] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_89 bl[89] br[89] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_90 bl[90] br[90] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_90 bl[90] br[90] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_91 bl[91] br[91] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_91 bl[91] br[91] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_92 bl[92] br[92] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_92 bl[92] br[92] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_93 bl[93] br[93] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_93 bl[93] br[93] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_94 bl[94] br[94] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_94 bl[94] br[94] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_95 bl[95] br[95] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_95 bl[95] br[95] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_96 bl[96] br[96] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_96 bl[96] br[96] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_97 bl[97] br[97] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_97 bl[97] br[97] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_98 bl[98] br[98] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_98 bl[98] br[98] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_99 bl[99] br[99] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_99 bl[99] br[99] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_100 bl[100] br[100] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_100 bl[100] br[100] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_101 bl[101] br[101] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_101 bl[101] br[101] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_102 bl[102] br[102] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_102 bl[102] br[102] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_103 bl[103] br[103] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_103 bl[103] br[103] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_104 bl[104] br[104] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_104 bl[104] br[104] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_105 bl[105] br[105] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_105 bl[105] br[105] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_106 bl[106] br[106] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_106 bl[106] br[106] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_107 bl[107] br[107] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_107 bl[107] br[107] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_108 bl[108] br[108] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_108 bl[108] br[108] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_109 bl[109] br[109] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_109 bl[109] br[109] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_110 bl[110] br[110] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_110 bl[110] br[110] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_111 bl[111] br[111] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_111 bl[111] br[111] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_112 bl[112] br[112] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_112 bl[112] br[112] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_113 bl[113] br[113] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_113 bl[113] br[113] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_114 bl[114] br[114] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_114 bl[114] br[114] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_115 bl[115] br[115] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_115 bl[115] br[115] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_116 bl[116] br[116] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_116 bl[116] br[116] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_117 bl[117] br[117] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_117 bl[117] br[117] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_118 bl[118] br[118] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_118 bl[118] br[118] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_119 bl[119] br[119] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_119 bl[119] br[119] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_120 bl[120] br[120] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_120 bl[120] br[120] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_121 bl[121] br[121] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_121 bl[121] br[121] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_122 bl[122] br[122] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_122 bl[122] br[122] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_123 bl[123] br[123] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_123 bl[123] br[123] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_124 bl[124] br[124] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_124 bl[124] br[124] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_125 bl[125] br[125] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_125 bl[125] br[125] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_126 bl[126] br[126] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_126 bl[126] br[126] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_127 bl[127] br[127] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_127 bl[127] br[127] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_128 bl[128] br[128] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_128 bl[128] br[128] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_129 bl[129] br[129] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_129 bl[129] br[129] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_130 bl[130] br[130] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_130 bl[130] br[130] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_131 bl[131] br[131] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_131 bl[131] br[131] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_132 bl[132] br[132] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_132 bl[132] br[132] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_133 bl[133] br[133] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_133 bl[133] br[133] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_134 bl[134] br[134] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_134 bl[134] br[134] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_135 bl[135] br[135] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_135 bl[135] br[135] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_136 bl[136] br[136] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_136 bl[136] br[136] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_137 bl[137] br[137] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_137 bl[137] br[137] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_138 bl[138] br[138] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_138 bl[138] br[138] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_139 bl[139] br[139] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_139 bl[139] br[139] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_140 bl[140] br[140] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_140 bl[140] br[140] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_141 bl[141] br[141] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_141 bl[141] br[141] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_142 bl[142] br[142] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_142 bl[142] br[142] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_143 bl[143] br[143] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_143 bl[143] br[143] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_144 bl[144] br[144] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_144 bl[144] br[144] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_145 bl[145] br[145] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_145 bl[145] br[145] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_146 bl[146] br[146] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_146 bl[146] br[146] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_147 bl[147] br[147] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_147 bl[147] br[147] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_148 bl[148] br[148] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_148 bl[148] br[148] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_149 bl[149] br[149] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_149 bl[149] br[149] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_150 bl[150] br[150] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_150 bl[150] br[150] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_151 bl[151] br[151] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_151 bl[151] br[151] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_152 bl[152] br[152] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_152 bl[152] br[152] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_153 bl[153] br[153] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_153 bl[153] br[153] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_154 bl[154] br[154] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_154 bl[154] br[154] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_155 bl[155] br[155] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_155 bl[155] br[155] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_156 bl[156] br[156] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_156 bl[156] br[156] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_157 bl[157] br[157] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_157 bl[157] br[157] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_158 bl[158] br[158] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_158 bl[158] br[158] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_159 bl[159] br[159] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_159 bl[159] br[159] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_160 bl[160] br[160] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_160 bl[160] br[160] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_161 bl[161] br[161] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_161 bl[161] br[161] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_162 bl[162] br[162] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_162 bl[162] br[162] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_163 bl[163] br[163] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_163 bl[163] br[163] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_164 bl[164] br[164] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_164 bl[164] br[164] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_165 bl[165] br[165] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_165 bl[165] br[165] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_166 bl[166] br[166] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_166 bl[166] br[166] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_167 bl[167] br[167] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_167 bl[167] br[167] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_168 bl[168] br[168] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_168 bl[168] br[168] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_169 bl[169] br[169] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_169 bl[169] br[169] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_170 bl[170] br[170] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_170 bl[170] br[170] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_171 bl[171] br[171] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_171 bl[171] br[171] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_172 bl[172] br[172] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_172 bl[172] br[172] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_173 bl[173] br[173] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_173 bl[173] br[173] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_174 bl[174] br[174] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_174 bl[174] br[174] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_175 bl[175] br[175] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_175 bl[175] br[175] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_176 bl[176] br[176] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_176 bl[176] br[176] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_177 bl[177] br[177] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_177 bl[177] br[177] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_178 bl[178] br[178] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_178 bl[178] br[178] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_179 bl[179] br[179] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_179 bl[179] br[179] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_180 bl[180] br[180] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_180 bl[180] br[180] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_181 bl[181] br[181] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_181 bl[181] br[181] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_182 bl[182] br[182] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_182 bl[182] br[182] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_183 bl[183] br[183] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_183 bl[183] br[183] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_184 bl[184] br[184] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_184 bl[184] br[184] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_185 bl[185] br[185] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_185 bl[185] br[185] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_186 bl[186] br[186] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_186 bl[186] br[186] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_187 bl[187] br[187] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_187 bl[187] br[187] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_188 bl[188] br[188] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_188 bl[188] br[188] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_189 bl[189] br[189] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_189 bl[189] br[189] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_190 bl[190] br[190] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_190 bl[190] br[190] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_191 bl[191] br[191] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_191 bl[191] br[191] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_192 bl[192] br[192] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_192 bl[192] br[192] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_193 bl[193] br[193] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_193 bl[193] br[193] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_194 bl[194] br[194] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_194 bl[194] br[194] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_195 bl[195] br[195] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_195 bl[195] br[195] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_196 bl[196] br[196] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_196 bl[196] br[196] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_197 bl[197] br[197] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_197 bl[197] br[197] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_198 bl[198] br[198] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_198 bl[198] br[198] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_199 bl[199] br[199] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_199 bl[199] br[199] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_200 bl[200] br[200] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_200 bl[200] br[200] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_201 bl[201] br[201] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_201 bl[201] br[201] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_202 bl[202] br[202] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_202 bl[202] br[202] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_203 bl[203] br[203] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_203 bl[203] br[203] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_204 bl[204] br[204] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_204 bl[204] br[204] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_205 bl[205] br[205] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_205 bl[205] br[205] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_206 bl[206] br[206] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_206 bl[206] br[206] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_207 bl[207] br[207] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_207 bl[207] br[207] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_208 bl[208] br[208] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_208 bl[208] br[208] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_209 bl[209] br[209] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_209 bl[209] br[209] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_210 bl[210] br[210] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_210 bl[210] br[210] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_211 bl[211] br[211] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_211 bl[211] br[211] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_212 bl[212] br[212] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_212 bl[212] br[212] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_213 bl[213] br[213] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_213 bl[213] br[213] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_214 bl[214] br[214] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_214 bl[214] br[214] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_215 bl[215] br[215] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_215 bl[215] br[215] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_216 bl[216] br[216] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_216 bl[216] br[216] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_217 bl[217] br[217] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_217 bl[217] br[217] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_218 bl[218] br[218] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_218 bl[218] br[218] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_219 bl[219] br[219] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_219 bl[219] br[219] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_220 bl[220] br[220] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_220 bl[220] br[220] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_221 bl[221] br[221] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_221 bl[221] br[221] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_222 bl[222] br[222] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_222 bl[222] br[222] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_223 bl[223] br[223] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_223 bl[223] br[223] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_224 bl[224] br[224] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_224 bl[224] br[224] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_225 bl[225] br[225] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_225 bl[225] br[225] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_226 bl[226] br[226] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_226 bl[226] br[226] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_227 bl[227] br[227] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_227 bl[227] br[227] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_228 bl[228] br[228] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_228 bl[228] br[228] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_229 bl[229] br[229] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_229 bl[229] br[229] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_230 bl[230] br[230] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_230 bl[230] br[230] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_231 bl[231] br[231] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_231 bl[231] br[231] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_232 bl[232] br[232] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_232 bl[232] br[232] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_233 bl[233] br[233] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_233 bl[233] br[233] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_234 bl[234] br[234] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_234 bl[234] br[234] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_235 bl[235] br[235] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_235 bl[235] br[235] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_236 bl[236] br[236] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_236 bl[236] br[236] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_237 bl[237] br[237] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_237 bl[237] br[237] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_238 bl[238] br[238] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_238 bl[238] br[238] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_239 bl[239] br[239] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_239 bl[239] br[239] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_240 bl[240] br[240] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_240 bl[240] br[240] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_241 bl[241] br[241] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_241 bl[241] br[241] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_242 bl[242] br[242] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_242 bl[242] br[242] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_243 bl[243] br[243] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_243 bl[243] br[243] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_244 bl[244] br[244] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_244 bl[244] br[244] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_245 bl[245] br[245] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_245 bl[245] br[245] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_246 bl[246] br[246] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_246 bl[246] br[246] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_247 bl[247] br[247] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_247 bl[247] br[247] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_248 bl[248] br[248] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_248 bl[248] br[248] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_249 bl[249] br[249] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_249 bl[249] br[249] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_250 bl[250] br[250] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_250 bl[250] br[250] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_251 bl[251] br[251] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_251 bl[251] br[251] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_252 bl[252] br[252] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_252 bl[252] br[252] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_253 bl[253] br[253] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_253 bl[253] br[253] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_254 bl[254] br[254] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_254 bl[254] br[254] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_255 bl[255] br[255] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_255 bl[255] br[255] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_256 bl[256] br[256] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_256 bl[256] br[256] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_257 bl[257] br[257] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_257 bl[257] br[257] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_258 bl[258] br[258] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_258 bl[258] br[258] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_259 bl[259] br[259] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_259 bl[259] br[259] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_260 bl[260] br[260] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_260 bl[260] br[260] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_261 bl[261] br[261] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_261 bl[261] br[261] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_262 bl[262] br[262] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_262 bl[262] br[262] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_263 bl[263] br[263] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_263 bl[263] br[263] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_264 bl[264] br[264] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_264 bl[264] br[264] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_265 bl[265] br[265] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_265 bl[265] br[265] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_266 bl[266] br[266] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_266 bl[266] br[266] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_267 bl[267] br[267] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_267 bl[267] br[267] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_268 bl[268] br[268] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_268 bl[268] br[268] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_269 bl[269] br[269] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_269 bl[269] br[269] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_270 bl[270] br[270] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_270 bl[270] br[270] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_271 bl[271] br[271] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_271 bl[271] br[271] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_272 bl[272] br[272] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_272 bl[272] br[272] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_273 bl[273] br[273] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_273 bl[273] br[273] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_274 bl[274] br[274] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_274 bl[274] br[274] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_275 bl[275] br[275] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_275 bl[275] br[275] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_276 bl[276] br[276] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_276 bl[276] br[276] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_277 bl[277] br[277] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_277 bl[277] br[277] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_278 bl[278] br[278] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_278 bl[278] br[278] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_279 bl[279] br[279] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_279 bl[279] br[279] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_280 bl[280] br[280] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_280 bl[280] br[280] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_281 bl[281] br[281] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_281 bl[281] br[281] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_282 bl[282] br[282] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_282 bl[282] br[282] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_283 bl[283] br[283] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_283 bl[283] br[283] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_284 bl[284] br[284] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_284 bl[284] br[284] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_285 bl[285] br[285] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_285 bl[285] br[285] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_286 bl[286] br[286] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_286 bl[286] br[286] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_287 bl[287] br[287] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_287 bl[287] br[287] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_288 bl[288] br[288] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_288 bl[288] br[288] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_289 bl[289] br[289] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_289 bl[289] br[289] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_290 bl[290] br[290] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_290 bl[290] br[290] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_291 bl[291] br[291] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_291 bl[291] br[291] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_292 bl[292] br[292] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_292 bl[292] br[292] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_293 bl[293] br[293] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_293 bl[293] br[293] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_294 bl[294] br[294] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_294 bl[294] br[294] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_295 bl[295] br[295] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_295 bl[295] br[295] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_296 bl[296] br[296] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_296 bl[296] br[296] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_297 bl[297] br[297] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_297 bl[297] br[297] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_298 bl[298] br[298] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_298 bl[298] br[298] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_299 bl[299] br[299] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_299 bl[299] br[299] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_300 bl[300] br[300] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_300 bl[300] br[300] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_301 bl[301] br[301] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_301 bl[301] br[301] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_302 bl[302] br[302] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_302 bl[302] br[302] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_303 bl[303] br[303] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_303 bl[303] br[303] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_304 bl[304] br[304] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_304 bl[304] br[304] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_305 bl[305] br[305] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_305 bl[305] br[305] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_306 bl[306] br[306] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_306 bl[306] br[306] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_307 bl[307] br[307] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_307 bl[307] br[307] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_308 bl[308] br[308] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_308 bl[308] br[308] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_309 bl[309] br[309] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_309 bl[309] br[309] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_310 bl[310] br[310] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_310 bl[310] br[310] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_311 bl[311] br[311] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_311 bl[311] br[311] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_312 bl[312] br[312] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_312 bl[312] br[312] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_313 bl[313] br[313] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_313 bl[313] br[313] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_314 bl[314] br[314] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_314 bl[314] br[314] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_315 bl[315] br[315] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_315 bl[315] br[315] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_316 bl[316] br[316] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_316 bl[316] br[316] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_317 bl[317] br[317] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_317 bl[317] br[317] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_318 bl[318] br[318] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_318 bl[318] br[318] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_319 bl[319] br[319] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_319 bl[319] br[319] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_320 bl[320] br[320] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_320 bl[320] br[320] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_321 bl[321] br[321] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_321 bl[321] br[321] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_322 bl[322] br[322] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_322 bl[322] br[322] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_323 bl[323] br[323] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_323 bl[323] br[323] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_324 bl[324] br[324] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_324 bl[324] br[324] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_325 bl[325] br[325] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_325 bl[325] br[325] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_326 bl[326] br[326] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_326 bl[326] br[326] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_327 bl[327] br[327] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_327 bl[327] br[327] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_328 bl[328] br[328] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_328 bl[328] br[328] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_329 bl[329] br[329] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_329 bl[329] br[329] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_330 bl[330] br[330] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_330 bl[330] br[330] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_331 bl[331] br[331] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_331 bl[331] br[331] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_332 bl[332] br[332] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_332 bl[332] br[332] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_333 bl[333] br[333] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_333 bl[333] br[333] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_334 bl[334] br[334] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_334 bl[334] br[334] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_335 bl[335] br[335] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_335 bl[335] br[335] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_336 bl[336] br[336] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_336 bl[336] br[336] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_337 bl[337] br[337] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_337 bl[337] br[337] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_338 bl[338] br[338] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_338 bl[338] br[338] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_339 bl[339] br[339] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_339 bl[339] br[339] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_340 bl[340] br[340] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_340 bl[340] br[340] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_341 bl[341] br[341] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_341 bl[341] br[341] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_342 bl[342] br[342] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_342 bl[342] br[342] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_343 bl[343] br[343] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_343 bl[343] br[343] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_344 bl[344] br[344] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_344 bl[344] br[344] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_345 bl[345] br[345] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_345 bl[345] br[345] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_346 bl[346] br[346] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_346 bl[346] br[346] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_347 bl[347] br[347] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_347 bl[347] br[347] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_348 bl[348] br[348] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_348 bl[348] br[348] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_349 bl[349] br[349] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_349 bl[349] br[349] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_350 bl[350] br[350] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_350 bl[350] br[350] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_351 bl[351] br[351] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_351 bl[351] br[351] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_352 bl[352] br[352] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_352 bl[352] br[352] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_353 bl[353] br[353] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_353 bl[353] br[353] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_354 bl[354] br[354] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_354 bl[354] br[354] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_355 bl[355] br[355] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_355 bl[355] br[355] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_356 bl[356] br[356] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_356 bl[356] br[356] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_357 bl[357] br[357] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_357 bl[357] br[357] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_358 bl[358] br[358] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_358 bl[358] br[358] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_359 bl[359] br[359] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_359 bl[359] br[359] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_360 bl[360] br[360] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_360 bl[360] br[360] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_361 bl[361] br[361] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_361 bl[361] br[361] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_362 bl[362] br[362] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_362 bl[362] br[362] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_363 bl[363] br[363] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_363 bl[363] br[363] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_364 bl[364] br[364] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_364 bl[364] br[364] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_365 bl[365] br[365] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_365 bl[365] br[365] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_366 bl[366] br[366] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_366 bl[366] br[366] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_367 bl[367] br[367] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_367 bl[367] br[367] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_368 bl[368] br[368] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_368 bl[368] br[368] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_369 bl[369] br[369] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_369 bl[369] br[369] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_370 bl[370] br[370] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_370 bl[370] br[370] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_371 bl[371] br[371] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_371 bl[371] br[371] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_372 bl[372] br[372] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_372 bl[372] br[372] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_373 bl[373] br[373] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_373 bl[373] br[373] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_374 bl[374] br[374] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_374 bl[374] br[374] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_375 bl[375] br[375] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_375 bl[375] br[375] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_376 bl[376] br[376] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_376 bl[376] br[376] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_377 bl[377] br[377] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_377 bl[377] br[377] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_378 bl[378] br[378] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_378 bl[378] br[378] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_379 bl[379] br[379] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_379 bl[379] br[379] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_380 bl[380] br[380] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_380 bl[380] br[380] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_381 bl[381] br[381] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_381 bl[381] br[381] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_382 bl[382] br[382] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_382 bl[382] br[382] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_383 bl[383] br[383] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_383 bl[383] br[383] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_384 bl[384] br[384] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_384 bl[384] br[384] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_385 bl[385] br[385] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_385 bl[385] br[385] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_386 bl[386] br[386] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_386 bl[386] br[386] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_387 bl[387] br[387] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_387 bl[387] br[387] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_388 bl[388] br[388] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_388 bl[388] br[388] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_389 bl[389] br[389] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_389 bl[389] br[389] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_390 bl[390] br[390] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_390 bl[390] br[390] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_391 bl[391] br[391] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_391 bl[391] br[391] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_392 bl[392] br[392] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_392 bl[392] br[392] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_393 bl[393] br[393] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_393 bl[393] br[393] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_394 bl[394] br[394] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_394 bl[394] br[394] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_395 bl[395] br[395] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_395 bl[395] br[395] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_396 bl[396] br[396] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_396 bl[396] br[396] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_397 bl[397] br[397] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_397 bl[397] br[397] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_398 bl[398] br[398] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_398 bl[398] br[398] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_399 bl[399] br[399] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_399 bl[399] br[399] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_400 bl[400] br[400] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_400 bl[400] br[400] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_401 bl[401] br[401] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_401 bl[401] br[401] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_402 bl[402] br[402] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_402 bl[402] br[402] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_403 bl[403] br[403] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_403 bl[403] br[403] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_404 bl[404] br[404] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_404 bl[404] br[404] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_405 bl[405] br[405] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_405 bl[405] br[405] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_406 bl[406] br[406] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_406 bl[406] br[406] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_407 bl[407] br[407] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_407 bl[407] br[407] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_408 bl[408] br[408] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_408 bl[408] br[408] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_409 bl[409] br[409] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_409 bl[409] br[409] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_410 bl[410] br[410] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_410 bl[410] br[410] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_411 bl[411] br[411] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_411 bl[411] br[411] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_412 bl[412] br[412] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_412 bl[412] br[412] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_413 bl[413] br[413] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_413 bl[413] br[413] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_414 bl[414] br[414] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_414 bl[414] br[414] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_415 bl[415] br[415] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_415 bl[415] br[415] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_416 bl[416] br[416] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_416 bl[416] br[416] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_417 bl[417] br[417] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_417 bl[417] br[417] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_418 bl[418] br[418] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_418 bl[418] br[418] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_419 bl[419] br[419] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_419 bl[419] br[419] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_420 bl[420] br[420] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_420 bl[420] br[420] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_421 bl[421] br[421] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_421 bl[421] br[421] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_422 bl[422] br[422] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_422 bl[422] br[422] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_423 bl[423] br[423] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_423 bl[423] br[423] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_424 bl[424] br[424] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_424 bl[424] br[424] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_425 bl[425] br[425] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_425 bl[425] br[425] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_426 bl[426] br[426] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_426 bl[426] br[426] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_427 bl[427] br[427] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_427 bl[427] br[427] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_428 bl[428] br[428] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_428 bl[428] br[428] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_429 bl[429] br[429] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_429 bl[429] br[429] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_430 bl[430] br[430] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_430 bl[430] br[430] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_431 bl[431] br[431] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_431 bl[431] br[431] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_432 bl[432] br[432] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_432 bl[432] br[432] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_433 bl[433] br[433] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_433 bl[433] br[433] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_434 bl[434] br[434] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_434 bl[434] br[434] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_435 bl[435] br[435] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_435 bl[435] br[435] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_436 bl[436] br[436] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_436 bl[436] br[436] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_437 bl[437] br[437] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_437 bl[437] br[437] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_438 bl[438] br[438] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_438 bl[438] br[438] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_439 bl[439] br[439] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_439 bl[439] br[439] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_440 bl[440] br[440] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_440 bl[440] br[440] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_441 bl[441] br[441] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_441 bl[441] br[441] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_442 bl[442] br[442] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_442 bl[442] br[442] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_443 bl[443] br[443] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_443 bl[443] br[443] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_444 bl[444] br[444] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_444 bl[444] br[444] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_445 bl[445] br[445] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_445 bl[445] br[445] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_446 bl[446] br[446] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_446 bl[446] br[446] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_447 bl[447] br[447] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_447 bl[447] br[447] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_448 bl[448] br[448] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_448 bl[448] br[448] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_449 bl[449] br[449] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_449 bl[449] br[449] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_450 bl[450] br[450] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_450 bl[450] br[450] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_451 bl[451] br[451] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_451 bl[451] br[451] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_452 bl[452] br[452] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_452 bl[452] br[452] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_453 bl[453] br[453] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_453 bl[453] br[453] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_454 bl[454] br[454] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_454 bl[454] br[454] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_455 bl[455] br[455] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_455 bl[455] br[455] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_456 bl[456] br[456] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_456 bl[456] br[456] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_457 bl[457] br[457] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_457 bl[457] br[457] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_458 bl[458] br[458] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_458 bl[458] br[458] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_459 bl[459] br[459] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_459 bl[459] br[459] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_460 bl[460] br[460] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_460 bl[460] br[460] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_461 bl[461] br[461] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_461 bl[461] br[461] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_462 bl[462] br[462] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_462 bl[462] br[462] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_463 bl[463] br[463] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_463 bl[463] br[463] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_464 bl[464] br[464] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_464 bl[464] br[464] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_465 bl[465] br[465] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_465 bl[465] br[465] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_466 bl[466] br[466] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_466 bl[466] br[466] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_467 bl[467] br[467] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_467 bl[467] br[467] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_468 bl[468] br[468] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_468 bl[468] br[468] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_469 bl[469] br[469] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_469 bl[469] br[469] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_470 bl[470] br[470] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_470 bl[470] br[470] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_471 bl[471] br[471] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_471 bl[471] br[471] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_472 bl[472] br[472] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_472 bl[472] br[472] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_473 bl[473] br[473] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_473 bl[473] br[473] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_474 bl[474] br[474] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_474 bl[474] br[474] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_475 bl[475] br[475] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_475 bl[475] br[475] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_476 bl[476] br[476] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_476 bl[476] br[476] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_477 bl[477] br[477] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_477 bl[477] br[477] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_478 bl[478] br[478] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_478 bl[478] br[478] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_479 bl[479] br[479] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_479 bl[479] br[479] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_480 bl[480] br[480] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_480 bl[480] br[480] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_481 bl[481] br[481] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_481 bl[481] br[481] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_482 bl[482] br[482] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_482 bl[482] br[482] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_483 bl[483] br[483] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_483 bl[483] br[483] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_484 bl[484] br[484] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_484 bl[484] br[484] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_485 bl[485] br[485] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_485 bl[485] br[485] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_486 bl[486] br[486] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_486 bl[486] br[486] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_487 bl[487] br[487] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_487 bl[487] br[487] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_488 bl[488] br[488] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_488 bl[488] br[488] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_489 bl[489] br[489] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_489 bl[489] br[489] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_490 bl[490] br[490] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_490 bl[490] br[490] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_491 bl[491] br[491] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_491 bl[491] br[491] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_492 bl[492] br[492] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_492 bl[492] br[492] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_493 bl[493] br[493] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_493 bl[493] br[493] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_494 bl[494] br[494] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_494 bl[494] br[494] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_495 bl[495] br[495] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_495 bl[495] br[495] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_496 bl[496] br[496] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_496 bl[496] br[496] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_497 bl[497] br[497] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_497 bl[497] br[497] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_498 bl[498] br[498] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_498 bl[498] br[498] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_499 bl[499] br[499] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_499 bl[499] br[499] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_500 bl[500] br[500] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_500 bl[500] br[500] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_501 bl[501] br[501] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_501 bl[501] br[501] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_502 bl[502] br[502] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_502 bl[502] br[502] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_503 bl[503] br[503] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_503 bl[503] br[503] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_504 bl[504] br[504] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_504 bl[504] br[504] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_505 bl[505] br[505] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_505 bl[505] br[505] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_506 bl[506] br[506] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_506 bl[506] br[506] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_507 bl[507] br[507] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_507 bl[507] br[507] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_508 bl[508] br[508] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_508 bl[508] br[508] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_509 bl[509] br[509] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_509 bl[509] br[509] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_510 bl[510] br[510] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_510 bl[510] br[510] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_top_511 bl[511] br[511] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xdummy_row_bot_511 bl[511] br[511] vdd vss vss vss vdd sram_sp_cell_wrapper
  Xcolend_top_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_colend_wrapper
  Xcolend_bot_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_colend_wrapper
  Xhstrap_0_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_0 dummy_br vdd vss dummy_bl vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_1 br[0] vdd vss bl[0] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_1 br[0] vdd vss bl[0] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_1 br[0] vdd vss bl[0] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_2 br[1] vdd vss bl[1] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_2 br[1] vdd vss bl[1] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_2 br[1] vdd vss bl[1] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_3 br[2] vdd vss bl[2] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_3 br[2] vdd vss bl[2] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_3 br[2] vdd vss bl[2] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_4 br[3] vdd vss bl[3] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_4 br[3] vdd vss bl[3] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_4 br[3] vdd vss bl[3] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_5 br[4] vdd vss bl[4] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_5 br[4] vdd vss bl[4] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_5 br[4] vdd vss bl[4] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_6 br[5] vdd vss bl[5] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_6 br[5] vdd vss bl[5] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_6 br[5] vdd vss bl[5] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_7 br[6] vdd vss bl[6] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_7 br[6] vdd vss bl[6] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_7 br[6] vdd vss bl[6] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_8 br[7] vdd vss bl[7] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_8 br[7] vdd vss bl[7] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_8 br[7] vdd vss bl[7] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_9 br[8] vdd vss bl[8] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_9 br[8] vdd vss bl[8] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_9 br[8] vdd vss bl[8] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_10 br[9] vdd vss bl[9] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_10 br[9] vdd vss bl[9] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_10 br[9] vdd vss bl[9] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_11 br[10] vdd vss bl[10] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_11 br[10] vdd vss bl[10] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_11 br[10] vdd vss bl[10] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_12 br[11] vdd vss bl[11] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_12 br[11] vdd vss bl[11] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_12 br[11] vdd vss bl[11] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_13 br[12] vdd vss bl[12] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_13 br[12] vdd vss bl[12] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_13 br[12] vdd vss bl[12] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_14 br[13] vdd vss bl[13] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_14 br[13] vdd vss bl[13] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_14 br[13] vdd vss bl[13] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_15 br[14] vdd vss bl[14] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_15 br[14] vdd vss bl[14] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_15 br[14] vdd vss bl[14] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_16 br[15] vdd vss bl[15] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_16 br[15] vdd vss bl[15] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_16 br[15] vdd vss bl[15] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_17 br[16] vdd vss bl[16] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_17 br[16] vdd vss bl[16] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_17 br[16] vdd vss bl[16] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_18 br[17] vdd vss bl[17] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_18 br[17] vdd vss bl[17] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_18 br[17] vdd vss bl[17] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_19 br[18] vdd vss bl[18] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_19 br[18] vdd vss bl[18] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_19 br[18] vdd vss bl[18] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_20 br[19] vdd vss bl[19] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_20 br[19] vdd vss bl[19] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_20 br[19] vdd vss bl[19] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_21 br[20] vdd vss bl[20] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_21 br[20] vdd vss bl[20] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_21 br[20] vdd vss bl[20] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_22 br[21] vdd vss bl[21] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_22 br[21] vdd vss bl[21] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_22 br[21] vdd vss bl[21] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_23 br[22] vdd vss bl[22] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_23 br[22] vdd vss bl[22] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_23 br[22] vdd vss bl[22] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_24 br[23] vdd vss bl[23] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_24 br[23] vdd vss bl[23] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_24 br[23] vdd vss bl[23] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_25 br[24] vdd vss bl[24] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_25 br[24] vdd vss bl[24] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_25 br[24] vdd vss bl[24] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_26 br[25] vdd vss bl[25] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_26 br[25] vdd vss bl[25] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_26 br[25] vdd vss bl[25] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_27 br[26] vdd vss bl[26] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_27 br[26] vdd vss bl[26] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_27 br[26] vdd vss bl[26] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_28 br[27] vdd vss bl[27] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_28 br[27] vdd vss bl[27] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_28 br[27] vdd vss bl[27] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_29 br[28] vdd vss bl[28] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_29 br[28] vdd vss bl[28] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_29 br[28] vdd vss bl[28] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_30 br[29] vdd vss bl[29] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_30 br[29] vdd vss bl[29] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_30 br[29] vdd vss bl[29] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_31 br[30] vdd vss bl[30] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_31 br[30] vdd vss bl[30] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_31 br[30] vdd vss bl[30] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_32 br[31] vdd vss bl[31] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_32 br[31] vdd vss bl[31] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_32 br[31] vdd vss bl[31] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_33 br[32] vdd vss bl[32] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_33 br[32] vdd vss bl[32] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_33 br[32] vdd vss bl[32] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_34 br[33] vdd vss bl[33] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_34 br[33] vdd vss bl[33] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_34 br[33] vdd vss bl[33] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_35 br[34] vdd vss bl[34] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_35 br[34] vdd vss bl[34] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_35 br[34] vdd vss bl[34] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_36 br[35] vdd vss bl[35] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_36 br[35] vdd vss bl[35] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_36 br[35] vdd vss bl[35] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_37 br[36] vdd vss bl[36] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_37 br[36] vdd vss bl[36] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_37 br[36] vdd vss bl[36] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_38 br[37] vdd vss bl[37] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_38 br[37] vdd vss bl[37] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_38 br[37] vdd vss bl[37] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_39 br[38] vdd vss bl[38] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_39 br[38] vdd vss bl[38] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_39 br[38] vdd vss bl[38] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_40 br[39] vdd vss bl[39] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_40 br[39] vdd vss bl[39] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_40 br[39] vdd vss bl[39] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_41 br[40] vdd vss bl[40] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_41 br[40] vdd vss bl[40] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_41 br[40] vdd vss bl[40] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_42 br[41] vdd vss bl[41] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_42 br[41] vdd vss bl[41] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_42 br[41] vdd vss bl[41] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_43 br[42] vdd vss bl[42] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_43 br[42] vdd vss bl[42] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_43 br[42] vdd vss bl[42] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_44 br[43] vdd vss bl[43] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_44 br[43] vdd vss bl[43] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_44 br[43] vdd vss bl[43] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_45 br[44] vdd vss bl[44] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_45 br[44] vdd vss bl[44] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_45 br[44] vdd vss bl[44] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_46 br[45] vdd vss bl[45] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_46 br[45] vdd vss bl[45] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_46 br[45] vdd vss bl[45] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_47 br[46] vdd vss bl[46] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_47 br[46] vdd vss bl[46] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_47 br[46] vdd vss bl[46] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_48 br[47] vdd vss bl[47] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_48 br[47] vdd vss bl[47] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_48 br[47] vdd vss bl[47] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_49 br[48] vdd vss bl[48] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_49 br[48] vdd vss bl[48] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_49 br[48] vdd vss bl[48] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_50 br[49] vdd vss bl[49] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_50 br[49] vdd vss bl[49] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_50 br[49] vdd vss bl[49] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_51 br[50] vdd vss bl[50] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_51 br[50] vdd vss bl[50] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_51 br[50] vdd vss bl[50] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_52 br[51] vdd vss bl[51] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_52 br[51] vdd vss bl[51] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_52 br[51] vdd vss bl[51] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_53 br[52] vdd vss bl[52] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_53 br[52] vdd vss bl[52] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_53 br[52] vdd vss bl[52] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_54 br[53] vdd vss bl[53] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_54 br[53] vdd vss bl[53] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_54 br[53] vdd vss bl[53] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_55 br[54] vdd vss bl[54] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_55 br[54] vdd vss bl[54] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_55 br[54] vdd vss bl[54] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_56 br[55] vdd vss bl[55] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_56 br[55] vdd vss bl[55] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_56 br[55] vdd vss bl[55] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_57 br[56] vdd vss bl[56] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_57 br[56] vdd vss bl[56] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_57 br[56] vdd vss bl[56] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_58 br[57] vdd vss bl[57] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_58 br[57] vdd vss bl[57] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_58 br[57] vdd vss bl[57] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_59 br[58] vdd vss bl[58] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_59 br[58] vdd vss bl[58] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_59 br[58] vdd vss bl[58] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_60 br[59] vdd vss bl[59] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_60 br[59] vdd vss bl[59] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_60 br[59] vdd vss bl[59] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_61 br[60] vdd vss bl[60] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_61 br[60] vdd vss bl[60] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_61 br[60] vdd vss bl[60] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_62 br[61] vdd vss bl[61] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_62 br[61] vdd vss bl[61] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_62 br[61] vdd vss bl[61] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_63 br[62] vdd vss bl[62] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_63 br[62] vdd vss bl[62] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_63 br[62] vdd vss bl[62] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_64 br[63] vdd vss bl[63] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_64 br[63] vdd vss bl[63] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_64 br[63] vdd vss bl[63] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_65 br[64] vdd vss bl[64] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_65 br[64] vdd vss bl[64] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_65 br[64] vdd vss bl[64] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_65 br[64] vdd vss bl[64] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_65 br[64] vdd vss bl[64] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_65 br[64] vdd vss bl[64] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_65 br[64] vdd vss bl[64] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_65 br[64] vdd vss bl[64] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_65 br[64] vdd vss bl[64] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_65 br[64] vdd vss bl[64] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_65 br[64] vdd vss bl[64] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_65 br[64] vdd vss bl[64] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_65 br[64] vdd vss bl[64] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_65 br[64] vdd vss bl[64] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_65 br[64] vdd vss bl[64] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_65 br[64] vdd vss bl[64] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_65 br[64] vdd vss bl[64] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_65 br[64] vdd vss bl[64] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_65 br[64] vdd vss bl[64] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_66 br[65] vdd vss bl[65] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_66 br[65] vdd vss bl[65] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_66 br[65] vdd vss bl[65] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_66 br[65] vdd vss bl[65] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_66 br[65] vdd vss bl[65] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_66 br[65] vdd vss bl[65] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_66 br[65] vdd vss bl[65] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_66 br[65] vdd vss bl[65] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_66 br[65] vdd vss bl[65] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_66 br[65] vdd vss bl[65] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_66 br[65] vdd vss bl[65] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_66 br[65] vdd vss bl[65] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_66 br[65] vdd vss bl[65] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_66 br[65] vdd vss bl[65] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_66 br[65] vdd vss bl[65] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_66 br[65] vdd vss bl[65] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_66 br[65] vdd vss bl[65] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_66 br[65] vdd vss bl[65] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_66 br[65] vdd vss bl[65] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_67 br[66] vdd vss bl[66] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_67 br[66] vdd vss bl[66] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_67 br[66] vdd vss bl[66] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_67 br[66] vdd vss bl[66] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_67 br[66] vdd vss bl[66] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_67 br[66] vdd vss bl[66] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_67 br[66] vdd vss bl[66] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_67 br[66] vdd vss bl[66] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_67 br[66] vdd vss bl[66] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_67 br[66] vdd vss bl[66] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_67 br[66] vdd vss bl[66] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_67 br[66] vdd vss bl[66] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_67 br[66] vdd vss bl[66] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_67 br[66] vdd vss bl[66] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_67 br[66] vdd vss bl[66] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_67 br[66] vdd vss bl[66] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_67 br[66] vdd vss bl[66] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_67 br[66] vdd vss bl[66] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_67 br[66] vdd vss bl[66] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_68 br[67] vdd vss bl[67] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_68 br[67] vdd vss bl[67] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_68 br[67] vdd vss bl[67] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_68 br[67] vdd vss bl[67] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_68 br[67] vdd vss bl[67] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_68 br[67] vdd vss bl[67] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_68 br[67] vdd vss bl[67] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_68 br[67] vdd vss bl[67] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_68 br[67] vdd vss bl[67] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_68 br[67] vdd vss bl[67] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_68 br[67] vdd vss bl[67] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_68 br[67] vdd vss bl[67] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_68 br[67] vdd vss bl[67] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_68 br[67] vdd vss bl[67] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_68 br[67] vdd vss bl[67] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_68 br[67] vdd vss bl[67] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_68 br[67] vdd vss bl[67] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_68 br[67] vdd vss bl[67] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_68 br[67] vdd vss bl[67] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_69 br[68] vdd vss bl[68] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_69 br[68] vdd vss bl[68] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_69 br[68] vdd vss bl[68] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_69 br[68] vdd vss bl[68] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_69 br[68] vdd vss bl[68] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_69 br[68] vdd vss bl[68] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_69 br[68] vdd vss bl[68] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_69 br[68] vdd vss bl[68] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_69 br[68] vdd vss bl[68] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_69 br[68] vdd vss bl[68] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_69 br[68] vdd vss bl[68] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_69 br[68] vdd vss bl[68] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_69 br[68] vdd vss bl[68] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_69 br[68] vdd vss bl[68] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_69 br[68] vdd vss bl[68] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_69 br[68] vdd vss bl[68] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_69 br[68] vdd vss bl[68] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_69 br[68] vdd vss bl[68] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_69 br[68] vdd vss bl[68] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_70 br[69] vdd vss bl[69] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_70 br[69] vdd vss bl[69] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_70 br[69] vdd vss bl[69] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_70 br[69] vdd vss bl[69] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_70 br[69] vdd vss bl[69] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_70 br[69] vdd vss bl[69] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_70 br[69] vdd vss bl[69] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_70 br[69] vdd vss bl[69] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_70 br[69] vdd vss bl[69] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_70 br[69] vdd vss bl[69] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_70 br[69] vdd vss bl[69] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_70 br[69] vdd vss bl[69] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_70 br[69] vdd vss bl[69] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_70 br[69] vdd vss bl[69] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_70 br[69] vdd vss bl[69] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_70 br[69] vdd vss bl[69] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_70 br[69] vdd vss bl[69] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_70 br[69] vdd vss bl[69] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_70 br[69] vdd vss bl[69] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_71 br[70] vdd vss bl[70] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_71 br[70] vdd vss bl[70] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_71 br[70] vdd vss bl[70] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_71 br[70] vdd vss bl[70] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_71 br[70] vdd vss bl[70] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_71 br[70] vdd vss bl[70] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_71 br[70] vdd vss bl[70] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_71 br[70] vdd vss bl[70] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_71 br[70] vdd vss bl[70] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_71 br[70] vdd vss bl[70] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_71 br[70] vdd vss bl[70] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_71 br[70] vdd vss bl[70] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_71 br[70] vdd vss bl[70] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_71 br[70] vdd vss bl[70] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_71 br[70] vdd vss bl[70] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_71 br[70] vdd vss bl[70] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_71 br[70] vdd vss bl[70] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_71 br[70] vdd vss bl[70] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_71 br[70] vdd vss bl[70] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_72 br[71] vdd vss bl[71] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_72 br[71] vdd vss bl[71] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_72 br[71] vdd vss bl[71] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_72 br[71] vdd vss bl[71] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_72 br[71] vdd vss bl[71] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_72 br[71] vdd vss bl[71] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_72 br[71] vdd vss bl[71] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_72 br[71] vdd vss bl[71] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_72 br[71] vdd vss bl[71] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_72 br[71] vdd vss bl[71] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_72 br[71] vdd vss bl[71] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_72 br[71] vdd vss bl[71] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_72 br[71] vdd vss bl[71] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_72 br[71] vdd vss bl[71] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_72 br[71] vdd vss bl[71] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_72 br[71] vdd vss bl[71] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_72 br[71] vdd vss bl[71] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_72 br[71] vdd vss bl[71] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_72 br[71] vdd vss bl[71] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_73 br[72] vdd vss bl[72] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_73 br[72] vdd vss bl[72] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_73 br[72] vdd vss bl[72] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_73 br[72] vdd vss bl[72] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_73 br[72] vdd vss bl[72] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_73 br[72] vdd vss bl[72] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_73 br[72] vdd vss bl[72] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_73 br[72] vdd vss bl[72] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_73 br[72] vdd vss bl[72] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_73 br[72] vdd vss bl[72] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_73 br[72] vdd vss bl[72] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_73 br[72] vdd vss bl[72] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_73 br[72] vdd vss bl[72] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_73 br[72] vdd vss bl[72] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_73 br[72] vdd vss bl[72] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_73 br[72] vdd vss bl[72] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_73 br[72] vdd vss bl[72] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_73 br[72] vdd vss bl[72] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_73 br[72] vdd vss bl[72] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_74 br[73] vdd vss bl[73] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_74 br[73] vdd vss bl[73] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_74 br[73] vdd vss bl[73] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_74 br[73] vdd vss bl[73] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_74 br[73] vdd vss bl[73] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_74 br[73] vdd vss bl[73] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_74 br[73] vdd vss bl[73] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_74 br[73] vdd vss bl[73] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_74 br[73] vdd vss bl[73] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_74 br[73] vdd vss bl[73] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_74 br[73] vdd vss bl[73] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_74 br[73] vdd vss bl[73] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_74 br[73] vdd vss bl[73] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_74 br[73] vdd vss bl[73] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_74 br[73] vdd vss bl[73] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_74 br[73] vdd vss bl[73] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_74 br[73] vdd vss bl[73] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_74 br[73] vdd vss bl[73] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_74 br[73] vdd vss bl[73] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_75 br[74] vdd vss bl[74] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_75 br[74] vdd vss bl[74] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_75 br[74] vdd vss bl[74] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_75 br[74] vdd vss bl[74] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_75 br[74] vdd vss bl[74] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_75 br[74] vdd vss bl[74] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_75 br[74] vdd vss bl[74] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_75 br[74] vdd vss bl[74] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_75 br[74] vdd vss bl[74] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_75 br[74] vdd vss bl[74] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_75 br[74] vdd vss bl[74] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_75 br[74] vdd vss bl[74] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_75 br[74] vdd vss bl[74] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_75 br[74] vdd vss bl[74] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_75 br[74] vdd vss bl[74] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_75 br[74] vdd vss bl[74] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_75 br[74] vdd vss bl[74] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_75 br[74] vdd vss bl[74] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_75 br[74] vdd vss bl[74] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_76 br[75] vdd vss bl[75] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_76 br[75] vdd vss bl[75] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_76 br[75] vdd vss bl[75] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_76 br[75] vdd vss bl[75] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_76 br[75] vdd vss bl[75] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_76 br[75] vdd vss bl[75] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_76 br[75] vdd vss bl[75] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_76 br[75] vdd vss bl[75] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_76 br[75] vdd vss bl[75] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_76 br[75] vdd vss bl[75] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_76 br[75] vdd vss bl[75] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_76 br[75] vdd vss bl[75] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_76 br[75] vdd vss bl[75] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_76 br[75] vdd vss bl[75] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_76 br[75] vdd vss bl[75] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_76 br[75] vdd vss bl[75] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_76 br[75] vdd vss bl[75] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_76 br[75] vdd vss bl[75] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_76 br[75] vdd vss bl[75] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_77 br[76] vdd vss bl[76] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_77 br[76] vdd vss bl[76] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_77 br[76] vdd vss bl[76] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_77 br[76] vdd vss bl[76] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_77 br[76] vdd vss bl[76] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_77 br[76] vdd vss bl[76] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_77 br[76] vdd vss bl[76] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_77 br[76] vdd vss bl[76] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_77 br[76] vdd vss bl[76] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_77 br[76] vdd vss bl[76] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_77 br[76] vdd vss bl[76] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_77 br[76] vdd vss bl[76] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_77 br[76] vdd vss bl[76] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_77 br[76] vdd vss bl[76] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_77 br[76] vdd vss bl[76] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_77 br[76] vdd vss bl[76] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_77 br[76] vdd vss bl[76] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_77 br[76] vdd vss bl[76] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_77 br[76] vdd vss bl[76] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_78 br[77] vdd vss bl[77] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_78 br[77] vdd vss bl[77] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_78 br[77] vdd vss bl[77] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_78 br[77] vdd vss bl[77] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_78 br[77] vdd vss bl[77] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_78 br[77] vdd vss bl[77] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_78 br[77] vdd vss bl[77] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_78 br[77] vdd vss bl[77] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_78 br[77] vdd vss bl[77] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_78 br[77] vdd vss bl[77] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_78 br[77] vdd vss bl[77] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_78 br[77] vdd vss bl[77] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_78 br[77] vdd vss bl[77] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_78 br[77] vdd vss bl[77] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_78 br[77] vdd vss bl[77] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_78 br[77] vdd vss bl[77] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_78 br[77] vdd vss bl[77] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_78 br[77] vdd vss bl[77] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_78 br[77] vdd vss bl[77] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_79 br[78] vdd vss bl[78] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_79 br[78] vdd vss bl[78] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_79 br[78] vdd vss bl[78] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_79 br[78] vdd vss bl[78] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_79 br[78] vdd vss bl[78] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_79 br[78] vdd vss bl[78] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_79 br[78] vdd vss bl[78] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_79 br[78] vdd vss bl[78] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_79 br[78] vdd vss bl[78] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_79 br[78] vdd vss bl[78] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_79 br[78] vdd vss bl[78] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_79 br[78] vdd vss bl[78] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_79 br[78] vdd vss bl[78] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_79 br[78] vdd vss bl[78] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_79 br[78] vdd vss bl[78] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_79 br[78] vdd vss bl[78] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_79 br[78] vdd vss bl[78] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_79 br[78] vdd vss bl[78] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_79 br[78] vdd vss bl[78] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_80 br[79] vdd vss bl[79] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_80 br[79] vdd vss bl[79] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_80 br[79] vdd vss bl[79] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_80 br[79] vdd vss bl[79] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_80 br[79] vdd vss bl[79] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_80 br[79] vdd vss bl[79] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_80 br[79] vdd vss bl[79] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_80 br[79] vdd vss bl[79] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_80 br[79] vdd vss bl[79] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_80 br[79] vdd vss bl[79] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_80 br[79] vdd vss bl[79] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_80 br[79] vdd vss bl[79] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_80 br[79] vdd vss bl[79] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_80 br[79] vdd vss bl[79] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_80 br[79] vdd vss bl[79] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_80 br[79] vdd vss bl[79] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_80 br[79] vdd vss bl[79] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_80 br[79] vdd vss bl[79] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_80 br[79] vdd vss bl[79] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_81 br[80] vdd vss bl[80] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_81 br[80] vdd vss bl[80] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_81 br[80] vdd vss bl[80] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_81 br[80] vdd vss bl[80] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_81 br[80] vdd vss bl[80] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_81 br[80] vdd vss bl[80] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_81 br[80] vdd vss bl[80] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_81 br[80] vdd vss bl[80] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_81 br[80] vdd vss bl[80] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_81 br[80] vdd vss bl[80] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_81 br[80] vdd vss bl[80] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_81 br[80] vdd vss bl[80] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_81 br[80] vdd vss bl[80] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_81 br[80] vdd vss bl[80] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_81 br[80] vdd vss bl[80] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_81 br[80] vdd vss bl[80] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_81 br[80] vdd vss bl[80] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_81 br[80] vdd vss bl[80] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_81 br[80] vdd vss bl[80] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_82 br[81] vdd vss bl[81] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_82 br[81] vdd vss bl[81] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_82 br[81] vdd vss bl[81] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_82 br[81] vdd vss bl[81] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_82 br[81] vdd vss bl[81] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_82 br[81] vdd vss bl[81] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_82 br[81] vdd vss bl[81] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_82 br[81] vdd vss bl[81] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_82 br[81] vdd vss bl[81] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_82 br[81] vdd vss bl[81] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_82 br[81] vdd vss bl[81] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_82 br[81] vdd vss bl[81] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_82 br[81] vdd vss bl[81] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_82 br[81] vdd vss bl[81] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_82 br[81] vdd vss bl[81] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_82 br[81] vdd vss bl[81] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_82 br[81] vdd vss bl[81] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_82 br[81] vdd vss bl[81] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_82 br[81] vdd vss bl[81] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_83 br[82] vdd vss bl[82] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_83 br[82] vdd vss bl[82] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_83 br[82] vdd vss bl[82] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_83 br[82] vdd vss bl[82] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_83 br[82] vdd vss bl[82] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_83 br[82] vdd vss bl[82] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_83 br[82] vdd vss bl[82] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_83 br[82] vdd vss bl[82] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_83 br[82] vdd vss bl[82] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_83 br[82] vdd vss bl[82] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_83 br[82] vdd vss bl[82] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_83 br[82] vdd vss bl[82] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_83 br[82] vdd vss bl[82] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_83 br[82] vdd vss bl[82] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_83 br[82] vdd vss bl[82] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_83 br[82] vdd vss bl[82] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_83 br[82] vdd vss bl[82] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_83 br[82] vdd vss bl[82] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_83 br[82] vdd vss bl[82] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_84 br[83] vdd vss bl[83] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_84 br[83] vdd vss bl[83] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_84 br[83] vdd vss bl[83] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_84 br[83] vdd vss bl[83] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_84 br[83] vdd vss bl[83] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_84 br[83] vdd vss bl[83] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_84 br[83] vdd vss bl[83] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_84 br[83] vdd vss bl[83] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_84 br[83] vdd vss bl[83] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_84 br[83] vdd vss bl[83] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_84 br[83] vdd vss bl[83] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_84 br[83] vdd vss bl[83] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_84 br[83] vdd vss bl[83] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_84 br[83] vdd vss bl[83] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_84 br[83] vdd vss bl[83] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_84 br[83] vdd vss bl[83] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_84 br[83] vdd vss bl[83] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_84 br[83] vdd vss bl[83] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_84 br[83] vdd vss bl[83] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_85 br[84] vdd vss bl[84] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_85 br[84] vdd vss bl[84] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_85 br[84] vdd vss bl[84] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_85 br[84] vdd vss bl[84] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_85 br[84] vdd vss bl[84] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_85 br[84] vdd vss bl[84] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_85 br[84] vdd vss bl[84] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_85 br[84] vdd vss bl[84] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_85 br[84] vdd vss bl[84] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_85 br[84] vdd vss bl[84] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_85 br[84] vdd vss bl[84] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_85 br[84] vdd vss bl[84] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_85 br[84] vdd vss bl[84] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_85 br[84] vdd vss bl[84] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_85 br[84] vdd vss bl[84] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_85 br[84] vdd vss bl[84] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_85 br[84] vdd vss bl[84] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_85 br[84] vdd vss bl[84] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_85 br[84] vdd vss bl[84] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_86 br[85] vdd vss bl[85] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_86 br[85] vdd vss bl[85] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_86 br[85] vdd vss bl[85] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_86 br[85] vdd vss bl[85] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_86 br[85] vdd vss bl[85] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_86 br[85] vdd vss bl[85] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_86 br[85] vdd vss bl[85] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_86 br[85] vdd vss bl[85] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_86 br[85] vdd vss bl[85] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_86 br[85] vdd vss bl[85] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_86 br[85] vdd vss bl[85] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_86 br[85] vdd vss bl[85] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_86 br[85] vdd vss bl[85] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_86 br[85] vdd vss bl[85] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_86 br[85] vdd vss bl[85] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_86 br[85] vdd vss bl[85] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_86 br[85] vdd vss bl[85] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_86 br[85] vdd vss bl[85] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_86 br[85] vdd vss bl[85] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_87 br[86] vdd vss bl[86] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_87 br[86] vdd vss bl[86] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_87 br[86] vdd vss bl[86] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_87 br[86] vdd vss bl[86] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_87 br[86] vdd vss bl[86] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_87 br[86] vdd vss bl[86] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_87 br[86] vdd vss bl[86] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_87 br[86] vdd vss bl[86] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_87 br[86] vdd vss bl[86] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_87 br[86] vdd vss bl[86] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_87 br[86] vdd vss bl[86] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_87 br[86] vdd vss bl[86] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_87 br[86] vdd vss bl[86] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_87 br[86] vdd vss bl[86] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_87 br[86] vdd vss bl[86] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_87 br[86] vdd vss bl[86] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_87 br[86] vdd vss bl[86] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_87 br[86] vdd vss bl[86] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_87 br[86] vdd vss bl[86] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_88 br[87] vdd vss bl[87] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_88 br[87] vdd vss bl[87] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_88 br[87] vdd vss bl[87] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_88 br[87] vdd vss bl[87] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_88 br[87] vdd vss bl[87] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_88 br[87] vdd vss bl[87] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_88 br[87] vdd vss bl[87] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_88 br[87] vdd vss bl[87] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_88 br[87] vdd vss bl[87] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_88 br[87] vdd vss bl[87] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_88 br[87] vdd vss bl[87] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_88 br[87] vdd vss bl[87] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_88 br[87] vdd vss bl[87] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_88 br[87] vdd vss bl[87] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_88 br[87] vdd vss bl[87] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_88 br[87] vdd vss bl[87] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_88 br[87] vdd vss bl[87] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_88 br[87] vdd vss bl[87] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_88 br[87] vdd vss bl[87] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_89 br[88] vdd vss bl[88] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_89 br[88] vdd vss bl[88] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_89 br[88] vdd vss bl[88] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_89 br[88] vdd vss bl[88] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_89 br[88] vdd vss bl[88] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_89 br[88] vdd vss bl[88] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_89 br[88] vdd vss bl[88] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_89 br[88] vdd vss bl[88] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_89 br[88] vdd vss bl[88] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_89 br[88] vdd vss bl[88] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_89 br[88] vdd vss bl[88] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_89 br[88] vdd vss bl[88] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_89 br[88] vdd vss bl[88] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_89 br[88] vdd vss bl[88] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_89 br[88] vdd vss bl[88] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_89 br[88] vdd vss bl[88] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_89 br[88] vdd vss bl[88] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_89 br[88] vdd vss bl[88] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_89 br[88] vdd vss bl[88] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_90 br[89] vdd vss bl[89] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_90 br[89] vdd vss bl[89] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_90 br[89] vdd vss bl[89] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_90 br[89] vdd vss bl[89] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_90 br[89] vdd vss bl[89] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_90 br[89] vdd vss bl[89] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_90 br[89] vdd vss bl[89] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_90 br[89] vdd vss bl[89] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_90 br[89] vdd vss bl[89] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_90 br[89] vdd vss bl[89] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_90 br[89] vdd vss bl[89] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_90 br[89] vdd vss bl[89] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_90 br[89] vdd vss bl[89] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_90 br[89] vdd vss bl[89] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_90 br[89] vdd vss bl[89] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_90 br[89] vdd vss bl[89] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_90 br[89] vdd vss bl[89] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_90 br[89] vdd vss bl[89] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_90 br[89] vdd vss bl[89] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_91 br[90] vdd vss bl[90] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_91 br[90] vdd vss bl[90] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_91 br[90] vdd vss bl[90] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_91 br[90] vdd vss bl[90] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_91 br[90] vdd vss bl[90] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_91 br[90] vdd vss bl[90] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_91 br[90] vdd vss bl[90] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_91 br[90] vdd vss bl[90] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_91 br[90] vdd vss bl[90] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_91 br[90] vdd vss bl[90] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_91 br[90] vdd vss bl[90] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_91 br[90] vdd vss bl[90] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_91 br[90] vdd vss bl[90] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_91 br[90] vdd vss bl[90] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_91 br[90] vdd vss bl[90] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_91 br[90] vdd vss bl[90] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_91 br[90] vdd vss bl[90] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_91 br[90] vdd vss bl[90] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_91 br[90] vdd vss bl[90] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_92 br[91] vdd vss bl[91] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_92 br[91] vdd vss bl[91] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_92 br[91] vdd vss bl[91] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_92 br[91] vdd vss bl[91] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_92 br[91] vdd vss bl[91] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_92 br[91] vdd vss bl[91] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_92 br[91] vdd vss bl[91] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_92 br[91] vdd vss bl[91] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_92 br[91] vdd vss bl[91] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_92 br[91] vdd vss bl[91] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_92 br[91] vdd vss bl[91] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_92 br[91] vdd vss bl[91] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_92 br[91] vdd vss bl[91] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_92 br[91] vdd vss bl[91] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_92 br[91] vdd vss bl[91] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_92 br[91] vdd vss bl[91] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_92 br[91] vdd vss bl[91] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_92 br[91] vdd vss bl[91] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_92 br[91] vdd vss bl[91] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_93 br[92] vdd vss bl[92] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_93 br[92] vdd vss bl[92] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_93 br[92] vdd vss bl[92] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_93 br[92] vdd vss bl[92] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_93 br[92] vdd vss bl[92] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_93 br[92] vdd vss bl[92] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_93 br[92] vdd vss bl[92] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_93 br[92] vdd vss bl[92] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_93 br[92] vdd vss bl[92] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_93 br[92] vdd vss bl[92] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_93 br[92] vdd vss bl[92] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_93 br[92] vdd vss bl[92] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_93 br[92] vdd vss bl[92] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_93 br[92] vdd vss bl[92] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_93 br[92] vdd vss bl[92] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_93 br[92] vdd vss bl[92] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_93 br[92] vdd vss bl[92] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_93 br[92] vdd vss bl[92] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_93 br[92] vdd vss bl[92] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_94 br[93] vdd vss bl[93] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_94 br[93] vdd vss bl[93] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_94 br[93] vdd vss bl[93] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_94 br[93] vdd vss bl[93] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_94 br[93] vdd vss bl[93] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_94 br[93] vdd vss bl[93] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_94 br[93] vdd vss bl[93] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_94 br[93] vdd vss bl[93] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_94 br[93] vdd vss bl[93] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_94 br[93] vdd vss bl[93] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_94 br[93] vdd vss bl[93] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_94 br[93] vdd vss bl[93] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_94 br[93] vdd vss bl[93] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_94 br[93] vdd vss bl[93] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_94 br[93] vdd vss bl[93] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_94 br[93] vdd vss bl[93] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_94 br[93] vdd vss bl[93] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_94 br[93] vdd vss bl[93] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_94 br[93] vdd vss bl[93] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_95 br[94] vdd vss bl[94] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_95 br[94] vdd vss bl[94] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_95 br[94] vdd vss bl[94] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_95 br[94] vdd vss bl[94] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_95 br[94] vdd vss bl[94] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_95 br[94] vdd vss bl[94] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_95 br[94] vdd vss bl[94] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_95 br[94] vdd vss bl[94] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_95 br[94] vdd vss bl[94] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_95 br[94] vdd vss bl[94] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_95 br[94] vdd vss bl[94] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_95 br[94] vdd vss bl[94] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_95 br[94] vdd vss bl[94] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_95 br[94] vdd vss bl[94] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_95 br[94] vdd vss bl[94] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_95 br[94] vdd vss bl[94] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_95 br[94] vdd vss bl[94] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_95 br[94] vdd vss bl[94] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_95 br[94] vdd vss bl[94] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_96 br[95] vdd vss bl[95] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_96 br[95] vdd vss bl[95] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_96 br[95] vdd vss bl[95] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_96 br[95] vdd vss bl[95] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_96 br[95] vdd vss bl[95] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_96 br[95] vdd vss bl[95] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_96 br[95] vdd vss bl[95] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_96 br[95] vdd vss bl[95] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_96 br[95] vdd vss bl[95] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_96 br[95] vdd vss bl[95] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_96 br[95] vdd vss bl[95] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_96 br[95] vdd vss bl[95] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_96 br[95] vdd vss bl[95] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_96 br[95] vdd vss bl[95] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_96 br[95] vdd vss bl[95] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_96 br[95] vdd vss bl[95] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_96 br[95] vdd vss bl[95] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_96 br[95] vdd vss bl[95] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_96 br[95] vdd vss bl[95] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_97 br[96] vdd vss bl[96] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_97 br[96] vdd vss bl[96] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_97 br[96] vdd vss bl[96] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_97 br[96] vdd vss bl[96] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_97 br[96] vdd vss bl[96] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_97 br[96] vdd vss bl[96] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_97 br[96] vdd vss bl[96] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_97 br[96] vdd vss bl[96] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_97 br[96] vdd vss bl[96] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_97 br[96] vdd vss bl[96] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_97 br[96] vdd vss bl[96] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_97 br[96] vdd vss bl[96] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_97 br[96] vdd vss bl[96] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_97 br[96] vdd vss bl[96] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_97 br[96] vdd vss bl[96] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_97 br[96] vdd vss bl[96] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_97 br[96] vdd vss bl[96] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_97 br[96] vdd vss bl[96] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_97 br[96] vdd vss bl[96] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_98 br[97] vdd vss bl[97] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_98 br[97] vdd vss bl[97] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_98 br[97] vdd vss bl[97] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_98 br[97] vdd vss bl[97] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_98 br[97] vdd vss bl[97] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_98 br[97] vdd vss bl[97] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_98 br[97] vdd vss bl[97] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_98 br[97] vdd vss bl[97] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_98 br[97] vdd vss bl[97] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_98 br[97] vdd vss bl[97] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_98 br[97] vdd vss bl[97] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_98 br[97] vdd vss bl[97] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_98 br[97] vdd vss bl[97] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_98 br[97] vdd vss bl[97] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_98 br[97] vdd vss bl[97] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_98 br[97] vdd vss bl[97] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_98 br[97] vdd vss bl[97] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_98 br[97] vdd vss bl[97] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_98 br[97] vdd vss bl[97] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_99 br[98] vdd vss bl[98] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_99 br[98] vdd vss bl[98] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_99 br[98] vdd vss bl[98] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_99 br[98] vdd vss bl[98] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_99 br[98] vdd vss bl[98] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_99 br[98] vdd vss bl[98] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_99 br[98] vdd vss bl[98] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_99 br[98] vdd vss bl[98] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_99 br[98] vdd vss bl[98] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_99 br[98] vdd vss bl[98] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_99 br[98] vdd vss bl[98] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_99 br[98] vdd vss bl[98] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_99 br[98] vdd vss bl[98] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_99 br[98] vdd vss bl[98] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_99 br[98] vdd vss bl[98] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_99 br[98] vdd vss bl[98] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_99 br[98] vdd vss bl[98] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_99 br[98] vdd vss bl[98] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_99 br[98] vdd vss bl[98] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_100 br[99] vdd vss bl[99] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_100 br[99] vdd vss bl[99] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_100 br[99] vdd vss bl[99] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_100 br[99] vdd vss bl[99] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_100 br[99] vdd vss bl[99] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_100 br[99] vdd vss bl[99] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_100 br[99] vdd vss bl[99] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_100 br[99] vdd vss bl[99] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_100 br[99] vdd vss bl[99] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_100 br[99] vdd vss bl[99] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_100 br[99] vdd vss bl[99] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_100 br[99] vdd vss bl[99] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_100 br[99] vdd vss bl[99] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_100 br[99] vdd vss bl[99] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_100 br[99] vdd vss bl[99] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_100 br[99] vdd vss bl[99] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_100 br[99] vdd vss bl[99] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_100 br[99] vdd vss bl[99] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_100 br[99] vdd vss bl[99] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_101 br[100] vdd vss bl[100] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_101 br[100] vdd vss bl[100] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_101 br[100] vdd vss bl[100] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_101 br[100] vdd vss bl[100] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_101 br[100] vdd vss bl[100] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_101 br[100] vdd vss bl[100] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_101 br[100] vdd vss bl[100] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_101 br[100] vdd vss bl[100] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_101 br[100] vdd vss bl[100] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_101 br[100] vdd vss bl[100] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_101 br[100] vdd vss bl[100] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_101 br[100] vdd vss bl[100] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_101 br[100] vdd vss bl[100] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_101 br[100] vdd vss bl[100] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_101 br[100] vdd vss bl[100] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_101 br[100] vdd vss bl[100] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_101 br[100] vdd vss bl[100] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_101 br[100] vdd vss bl[100] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_101 br[100] vdd vss bl[100] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_102 br[101] vdd vss bl[101] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_102 br[101] vdd vss bl[101] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_102 br[101] vdd vss bl[101] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_102 br[101] vdd vss bl[101] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_102 br[101] vdd vss bl[101] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_102 br[101] vdd vss bl[101] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_102 br[101] vdd vss bl[101] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_102 br[101] vdd vss bl[101] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_102 br[101] vdd vss bl[101] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_102 br[101] vdd vss bl[101] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_102 br[101] vdd vss bl[101] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_102 br[101] vdd vss bl[101] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_102 br[101] vdd vss bl[101] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_102 br[101] vdd vss bl[101] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_102 br[101] vdd vss bl[101] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_102 br[101] vdd vss bl[101] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_102 br[101] vdd vss bl[101] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_102 br[101] vdd vss bl[101] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_102 br[101] vdd vss bl[101] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_103 br[102] vdd vss bl[102] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_103 br[102] vdd vss bl[102] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_103 br[102] vdd vss bl[102] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_103 br[102] vdd vss bl[102] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_103 br[102] vdd vss bl[102] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_103 br[102] vdd vss bl[102] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_103 br[102] vdd vss bl[102] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_103 br[102] vdd vss bl[102] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_103 br[102] vdd vss bl[102] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_103 br[102] vdd vss bl[102] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_103 br[102] vdd vss bl[102] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_103 br[102] vdd vss bl[102] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_103 br[102] vdd vss bl[102] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_103 br[102] vdd vss bl[102] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_103 br[102] vdd vss bl[102] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_103 br[102] vdd vss bl[102] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_103 br[102] vdd vss bl[102] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_103 br[102] vdd vss bl[102] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_103 br[102] vdd vss bl[102] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_104 br[103] vdd vss bl[103] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_104 br[103] vdd vss bl[103] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_104 br[103] vdd vss bl[103] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_104 br[103] vdd vss bl[103] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_104 br[103] vdd vss bl[103] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_104 br[103] vdd vss bl[103] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_104 br[103] vdd vss bl[103] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_104 br[103] vdd vss bl[103] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_104 br[103] vdd vss bl[103] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_104 br[103] vdd vss bl[103] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_104 br[103] vdd vss bl[103] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_104 br[103] vdd vss bl[103] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_104 br[103] vdd vss bl[103] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_104 br[103] vdd vss bl[103] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_104 br[103] vdd vss bl[103] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_104 br[103] vdd vss bl[103] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_104 br[103] vdd vss bl[103] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_104 br[103] vdd vss bl[103] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_104 br[103] vdd vss bl[103] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_105 br[104] vdd vss bl[104] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_105 br[104] vdd vss bl[104] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_105 br[104] vdd vss bl[104] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_105 br[104] vdd vss bl[104] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_105 br[104] vdd vss bl[104] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_105 br[104] vdd vss bl[104] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_105 br[104] vdd vss bl[104] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_105 br[104] vdd vss bl[104] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_105 br[104] vdd vss bl[104] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_105 br[104] vdd vss bl[104] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_105 br[104] vdd vss bl[104] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_105 br[104] vdd vss bl[104] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_105 br[104] vdd vss bl[104] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_105 br[104] vdd vss bl[104] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_105 br[104] vdd vss bl[104] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_105 br[104] vdd vss bl[104] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_105 br[104] vdd vss bl[104] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_105 br[104] vdd vss bl[104] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_105 br[104] vdd vss bl[104] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_106 br[105] vdd vss bl[105] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_106 br[105] vdd vss bl[105] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_106 br[105] vdd vss bl[105] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_106 br[105] vdd vss bl[105] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_106 br[105] vdd vss bl[105] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_106 br[105] vdd vss bl[105] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_106 br[105] vdd vss bl[105] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_106 br[105] vdd vss bl[105] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_106 br[105] vdd vss bl[105] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_106 br[105] vdd vss bl[105] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_106 br[105] vdd vss bl[105] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_106 br[105] vdd vss bl[105] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_106 br[105] vdd vss bl[105] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_106 br[105] vdd vss bl[105] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_106 br[105] vdd vss bl[105] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_106 br[105] vdd vss bl[105] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_106 br[105] vdd vss bl[105] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_106 br[105] vdd vss bl[105] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_106 br[105] vdd vss bl[105] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_107 br[106] vdd vss bl[106] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_107 br[106] vdd vss bl[106] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_107 br[106] vdd vss bl[106] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_107 br[106] vdd vss bl[106] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_107 br[106] vdd vss bl[106] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_107 br[106] vdd vss bl[106] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_107 br[106] vdd vss bl[106] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_107 br[106] vdd vss bl[106] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_107 br[106] vdd vss bl[106] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_107 br[106] vdd vss bl[106] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_107 br[106] vdd vss bl[106] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_107 br[106] vdd vss bl[106] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_107 br[106] vdd vss bl[106] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_107 br[106] vdd vss bl[106] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_107 br[106] vdd vss bl[106] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_107 br[106] vdd vss bl[106] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_107 br[106] vdd vss bl[106] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_107 br[106] vdd vss bl[106] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_107 br[106] vdd vss bl[106] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_108 br[107] vdd vss bl[107] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_108 br[107] vdd vss bl[107] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_108 br[107] vdd vss bl[107] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_108 br[107] vdd vss bl[107] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_108 br[107] vdd vss bl[107] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_108 br[107] vdd vss bl[107] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_108 br[107] vdd vss bl[107] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_108 br[107] vdd vss bl[107] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_108 br[107] vdd vss bl[107] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_108 br[107] vdd vss bl[107] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_108 br[107] vdd vss bl[107] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_108 br[107] vdd vss bl[107] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_108 br[107] vdd vss bl[107] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_108 br[107] vdd vss bl[107] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_108 br[107] vdd vss bl[107] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_108 br[107] vdd vss bl[107] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_108 br[107] vdd vss bl[107] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_108 br[107] vdd vss bl[107] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_108 br[107] vdd vss bl[107] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_109 br[108] vdd vss bl[108] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_109 br[108] vdd vss bl[108] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_109 br[108] vdd vss bl[108] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_109 br[108] vdd vss bl[108] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_109 br[108] vdd vss bl[108] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_109 br[108] vdd vss bl[108] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_109 br[108] vdd vss bl[108] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_109 br[108] vdd vss bl[108] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_109 br[108] vdd vss bl[108] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_109 br[108] vdd vss bl[108] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_109 br[108] vdd vss bl[108] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_109 br[108] vdd vss bl[108] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_109 br[108] vdd vss bl[108] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_109 br[108] vdd vss bl[108] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_109 br[108] vdd vss bl[108] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_109 br[108] vdd vss bl[108] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_109 br[108] vdd vss bl[108] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_109 br[108] vdd vss bl[108] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_109 br[108] vdd vss bl[108] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_110 br[109] vdd vss bl[109] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_110 br[109] vdd vss bl[109] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_110 br[109] vdd vss bl[109] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_110 br[109] vdd vss bl[109] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_110 br[109] vdd vss bl[109] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_110 br[109] vdd vss bl[109] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_110 br[109] vdd vss bl[109] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_110 br[109] vdd vss bl[109] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_110 br[109] vdd vss bl[109] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_110 br[109] vdd vss bl[109] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_110 br[109] vdd vss bl[109] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_110 br[109] vdd vss bl[109] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_110 br[109] vdd vss bl[109] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_110 br[109] vdd vss bl[109] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_110 br[109] vdd vss bl[109] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_110 br[109] vdd vss bl[109] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_110 br[109] vdd vss bl[109] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_110 br[109] vdd vss bl[109] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_110 br[109] vdd vss bl[109] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_111 br[110] vdd vss bl[110] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_111 br[110] vdd vss bl[110] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_111 br[110] vdd vss bl[110] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_111 br[110] vdd vss bl[110] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_111 br[110] vdd vss bl[110] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_111 br[110] vdd vss bl[110] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_111 br[110] vdd vss bl[110] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_111 br[110] vdd vss bl[110] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_111 br[110] vdd vss bl[110] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_111 br[110] vdd vss bl[110] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_111 br[110] vdd vss bl[110] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_111 br[110] vdd vss bl[110] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_111 br[110] vdd vss bl[110] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_111 br[110] vdd vss bl[110] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_111 br[110] vdd vss bl[110] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_111 br[110] vdd vss bl[110] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_111 br[110] vdd vss bl[110] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_111 br[110] vdd vss bl[110] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_111 br[110] vdd vss bl[110] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_112 br[111] vdd vss bl[111] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_112 br[111] vdd vss bl[111] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_112 br[111] vdd vss bl[111] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_112 br[111] vdd vss bl[111] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_112 br[111] vdd vss bl[111] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_112 br[111] vdd vss bl[111] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_112 br[111] vdd vss bl[111] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_112 br[111] vdd vss bl[111] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_112 br[111] vdd vss bl[111] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_112 br[111] vdd vss bl[111] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_112 br[111] vdd vss bl[111] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_112 br[111] vdd vss bl[111] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_112 br[111] vdd vss bl[111] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_112 br[111] vdd vss bl[111] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_112 br[111] vdd vss bl[111] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_112 br[111] vdd vss bl[111] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_112 br[111] vdd vss bl[111] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_112 br[111] vdd vss bl[111] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_112 br[111] vdd vss bl[111] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_113 br[112] vdd vss bl[112] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_113 br[112] vdd vss bl[112] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_113 br[112] vdd vss bl[112] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_113 br[112] vdd vss bl[112] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_113 br[112] vdd vss bl[112] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_113 br[112] vdd vss bl[112] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_113 br[112] vdd vss bl[112] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_113 br[112] vdd vss bl[112] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_113 br[112] vdd vss bl[112] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_113 br[112] vdd vss bl[112] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_113 br[112] vdd vss bl[112] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_113 br[112] vdd vss bl[112] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_113 br[112] vdd vss bl[112] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_113 br[112] vdd vss bl[112] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_113 br[112] vdd vss bl[112] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_113 br[112] vdd vss bl[112] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_113 br[112] vdd vss bl[112] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_113 br[112] vdd vss bl[112] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_113 br[112] vdd vss bl[112] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_114 br[113] vdd vss bl[113] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_114 br[113] vdd vss bl[113] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_114 br[113] vdd vss bl[113] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_114 br[113] vdd vss bl[113] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_114 br[113] vdd vss bl[113] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_114 br[113] vdd vss bl[113] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_114 br[113] vdd vss bl[113] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_114 br[113] vdd vss bl[113] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_114 br[113] vdd vss bl[113] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_114 br[113] vdd vss bl[113] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_114 br[113] vdd vss bl[113] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_114 br[113] vdd vss bl[113] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_114 br[113] vdd vss bl[113] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_114 br[113] vdd vss bl[113] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_114 br[113] vdd vss bl[113] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_114 br[113] vdd vss bl[113] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_114 br[113] vdd vss bl[113] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_114 br[113] vdd vss bl[113] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_114 br[113] vdd vss bl[113] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_115 br[114] vdd vss bl[114] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_115 br[114] vdd vss bl[114] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_115 br[114] vdd vss bl[114] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_115 br[114] vdd vss bl[114] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_115 br[114] vdd vss bl[114] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_115 br[114] vdd vss bl[114] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_115 br[114] vdd vss bl[114] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_115 br[114] vdd vss bl[114] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_115 br[114] vdd vss bl[114] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_115 br[114] vdd vss bl[114] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_115 br[114] vdd vss bl[114] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_115 br[114] vdd vss bl[114] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_115 br[114] vdd vss bl[114] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_115 br[114] vdd vss bl[114] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_115 br[114] vdd vss bl[114] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_115 br[114] vdd vss bl[114] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_115 br[114] vdd vss bl[114] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_115 br[114] vdd vss bl[114] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_115 br[114] vdd vss bl[114] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_116 br[115] vdd vss bl[115] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_116 br[115] vdd vss bl[115] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_116 br[115] vdd vss bl[115] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_116 br[115] vdd vss bl[115] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_116 br[115] vdd vss bl[115] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_116 br[115] vdd vss bl[115] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_116 br[115] vdd vss bl[115] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_116 br[115] vdd vss bl[115] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_116 br[115] vdd vss bl[115] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_116 br[115] vdd vss bl[115] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_116 br[115] vdd vss bl[115] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_116 br[115] vdd vss bl[115] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_116 br[115] vdd vss bl[115] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_116 br[115] vdd vss bl[115] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_116 br[115] vdd vss bl[115] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_116 br[115] vdd vss bl[115] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_116 br[115] vdd vss bl[115] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_116 br[115] vdd vss bl[115] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_116 br[115] vdd vss bl[115] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_117 br[116] vdd vss bl[116] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_117 br[116] vdd vss bl[116] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_117 br[116] vdd vss bl[116] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_117 br[116] vdd vss bl[116] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_117 br[116] vdd vss bl[116] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_117 br[116] vdd vss bl[116] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_117 br[116] vdd vss bl[116] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_117 br[116] vdd vss bl[116] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_117 br[116] vdd vss bl[116] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_117 br[116] vdd vss bl[116] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_117 br[116] vdd vss bl[116] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_117 br[116] vdd vss bl[116] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_117 br[116] vdd vss bl[116] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_117 br[116] vdd vss bl[116] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_117 br[116] vdd vss bl[116] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_117 br[116] vdd vss bl[116] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_117 br[116] vdd vss bl[116] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_117 br[116] vdd vss bl[116] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_117 br[116] vdd vss bl[116] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_118 br[117] vdd vss bl[117] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_118 br[117] vdd vss bl[117] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_118 br[117] vdd vss bl[117] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_118 br[117] vdd vss bl[117] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_118 br[117] vdd vss bl[117] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_118 br[117] vdd vss bl[117] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_118 br[117] vdd vss bl[117] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_118 br[117] vdd vss bl[117] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_118 br[117] vdd vss bl[117] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_118 br[117] vdd vss bl[117] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_118 br[117] vdd vss bl[117] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_118 br[117] vdd vss bl[117] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_118 br[117] vdd vss bl[117] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_118 br[117] vdd vss bl[117] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_118 br[117] vdd vss bl[117] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_118 br[117] vdd vss bl[117] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_118 br[117] vdd vss bl[117] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_118 br[117] vdd vss bl[117] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_118 br[117] vdd vss bl[117] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_119 br[118] vdd vss bl[118] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_119 br[118] vdd vss bl[118] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_119 br[118] vdd vss bl[118] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_119 br[118] vdd vss bl[118] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_119 br[118] vdd vss bl[118] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_119 br[118] vdd vss bl[118] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_119 br[118] vdd vss bl[118] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_119 br[118] vdd vss bl[118] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_119 br[118] vdd vss bl[118] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_119 br[118] vdd vss bl[118] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_119 br[118] vdd vss bl[118] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_119 br[118] vdd vss bl[118] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_119 br[118] vdd vss bl[118] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_119 br[118] vdd vss bl[118] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_119 br[118] vdd vss bl[118] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_119 br[118] vdd vss bl[118] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_119 br[118] vdd vss bl[118] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_119 br[118] vdd vss bl[118] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_119 br[118] vdd vss bl[118] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_120 br[119] vdd vss bl[119] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_120 br[119] vdd vss bl[119] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_120 br[119] vdd vss bl[119] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_120 br[119] vdd vss bl[119] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_120 br[119] vdd vss bl[119] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_120 br[119] vdd vss bl[119] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_120 br[119] vdd vss bl[119] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_120 br[119] vdd vss bl[119] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_120 br[119] vdd vss bl[119] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_120 br[119] vdd vss bl[119] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_120 br[119] vdd vss bl[119] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_120 br[119] vdd vss bl[119] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_120 br[119] vdd vss bl[119] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_120 br[119] vdd vss bl[119] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_120 br[119] vdd vss bl[119] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_120 br[119] vdd vss bl[119] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_120 br[119] vdd vss bl[119] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_120 br[119] vdd vss bl[119] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_120 br[119] vdd vss bl[119] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_121 br[120] vdd vss bl[120] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_121 br[120] vdd vss bl[120] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_121 br[120] vdd vss bl[120] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_121 br[120] vdd vss bl[120] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_121 br[120] vdd vss bl[120] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_121 br[120] vdd vss bl[120] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_121 br[120] vdd vss bl[120] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_121 br[120] vdd vss bl[120] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_121 br[120] vdd vss bl[120] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_121 br[120] vdd vss bl[120] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_121 br[120] vdd vss bl[120] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_121 br[120] vdd vss bl[120] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_121 br[120] vdd vss bl[120] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_121 br[120] vdd vss bl[120] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_121 br[120] vdd vss bl[120] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_121 br[120] vdd vss bl[120] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_121 br[120] vdd vss bl[120] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_121 br[120] vdd vss bl[120] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_121 br[120] vdd vss bl[120] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_122 br[121] vdd vss bl[121] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_122 br[121] vdd vss bl[121] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_122 br[121] vdd vss bl[121] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_122 br[121] vdd vss bl[121] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_122 br[121] vdd vss bl[121] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_122 br[121] vdd vss bl[121] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_122 br[121] vdd vss bl[121] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_122 br[121] vdd vss bl[121] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_122 br[121] vdd vss bl[121] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_122 br[121] vdd vss bl[121] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_122 br[121] vdd vss bl[121] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_122 br[121] vdd vss bl[121] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_122 br[121] vdd vss bl[121] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_122 br[121] vdd vss bl[121] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_122 br[121] vdd vss bl[121] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_122 br[121] vdd vss bl[121] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_122 br[121] vdd vss bl[121] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_122 br[121] vdd vss bl[121] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_122 br[121] vdd vss bl[121] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_123 br[122] vdd vss bl[122] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_123 br[122] vdd vss bl[122] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_123 br[122] vdd vss bl[122] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_123 br[122] vdd vss bl[122] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_123 br[122] vdd vss bl[122] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_123 br[122] vdd vss bl[122] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_123 br[122] vdd vss bl[122] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_123 br[122] vdd vss bl[122] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_123 br[122] vdd vss bl[122] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_123 br[122] vdd vss bl[122] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_123 br[122] vdd vss bl[122] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_123 br[122] vdd vss bl[122] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_123 br[122] vdd vss bl[122] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_123 br[122] vdd vss bl[122] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_123 br[122] vdd vss bl[122] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_123 br[122] vdd vss bl[122] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_123 br[122] vdd vss bl[122] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_123 br[122] vdd vss bl[122] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_123 br[122] vdd vss bl[122] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_124 br[123] vdd vss bl[123] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_124 br[123] vdd vss bl[123] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_124 br[123] vdd vss bl[123] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_124 br[123] vdd vss bl[123] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_124 br[123] vdd vss bl[123] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_124 br[123] vdd vss bl[123] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_124 br[123] vdd vss bl[123] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_124 br[123] vdd vss bl[123] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_124 br[123] vdd vss bl[123] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_124 br[123] vdd vss bl[123] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_124 br[123] vdd vss bl[123] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_124 br[123] vdd vss bl[123] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_124 br[123] vdd vss bl[123] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_124 br[123] vdd vss bl[123] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_124 br[123] vdd vss bl[123] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_124 br[123] vdd vss bl[123] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_124 br[123] vdd vss bl[123] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_124 br[123] vdd vss bl[123] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_124 br[123] vdd vss bl[123] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_125 br[124] vdd vss bl[124] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_125 br[124] vdd vss bl[124] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_125 br[124] vdd vss bl[124] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_125 br[124] vdd vss bl[124] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_125 br[124] vdd vss bl[124] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_125 br[124] vdd vss bl[124] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_125 br[124] vdd vss bl[124] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_125 br[124] vdd vss bl[124] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_125 br[124] vdd vss bl[124] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_125 br[124] vdd vss bl[124] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_125 br[124] vdd vss bl[124] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_125 br[124] vdd vss bl[124] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_125 br[124] vdd vss bl[124] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_125 br[124] vdd vss bl[124] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_125 br[124] vdd vss bl[124] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_125 br[124] vdd vss bl[124] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_125 br[124] vdd vss bl[124] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_125 br[124] vdd vss bl[124] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_125 br[124] vdd vss bl[124] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_126 br[125] vdd vss bl[125] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_126 br[125] vdd vss bl[125] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_126 br[125] vdd vss bl[125] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_126 br[125] vdd vss bl[125] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_126 br[125] vdd vss bl[125] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_126 br[125] vdd vss bl[125] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_126 br[125] vdd vss bl[125] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_126 br[125] vdd vss bl[125] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_126 br[125] vdd vss bl[125] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_126 br[125] vdd vss bl[125] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_126 br[125] vdd vss bl[125] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_126 br[125] vdd vss bl[125] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_126 br[125] vdd vss bl[125] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_126 br[125] vdd vss bl[125] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_126 br[125] vdd vss bl[125] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_126 br[125] vdd vss bl[125] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_126 br[125] vdd vss bl[125] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_126 br[125] vdd vss bl[125] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_126 br[125] vdd vss bl[125] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_127 br[126] vdd vss bl[126] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_127 br[126] vdd vss bl[126] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_127 br[126] vdd vss bl[126] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_127 br[126] vdd vss bl[126] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_127 br[126] vdd vss bl[126] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_127 br[126] vdd vss bl[126] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_127 br[126] vdd vss bl[126] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_127 br[126] vdd vss bl[126] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_127 br[126] vdd vss bl[126] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_127 br[126] vdd vss bl[126] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_127 br[126] vdd vss bl[126] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_127 br[126] vdd vss bl[126] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_127 br[126] vdd vss bl[126] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_127 br[126] vdd vss bl[126] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_127 br[126] vdd vss bl[126] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_127 br[126] vdd vss bl[126] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_127 br[126] vdd vss bl[126] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_127 br[126] vdd vss bl[126] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_127 br[126] vdd vss bl[126] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_128 br[127] vdd vss bl[127] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_128 br[127] vdd vss bl[127] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_128 br[127] vdd vss bl[127] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_128 br[127] vdd vss bl[127] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_128 br[127] vdd vss bl[127] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_128 br[127] vdd vss bl[127] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_128 br[127] vdd vss bl[127] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_128 br[127] vdd vss bl[127] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_128 br[127] vdd vss bl[127] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_128 br[127] vdd vss bl[127] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_128 br[127] vdd vss bl[127] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_128 br[127] vdd vss bl[127] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_128 br[127] vdd vss bl[127] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_128 br[127] vdd vss bl[127] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_128 br[127] vdd vss bl[127] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_128 br[127] vdd vss bl[127] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_128 br[127] vdd vss bl[127] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_128 br[127] vdd vss bl[127] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_128 br[127] vdd vss bl[127] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_129 br[128] vdd vss bl[128] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_129 br[128] vdd vss bl[128] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_129 br[128] vdd vss bl[128] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_129 br[128] vdd vss bl[128] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_129 br[128] vdd vss bl[128] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_129 br[128] vdd vss bl[128] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_129 br[128] vdd vss bl[128] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_129 br[128] vdd vss bl[128] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_129 br[128] vdd vss bl[128] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_129 br[128] vdd vss bl[128] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_129 br[128] vdd vss bl[128] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_129 br[128] vdd vss bl[128] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_129 br[128] vdd vss bl[128] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_129 br[128] vdd vss bl[128] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_129 br[128] vdd vss bl[128] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_129 br[128] vdd vss bl[128] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_129 br[128] vdd vss bl[128] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_129 br[128] vdd vss bl[128] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_129 br[128] vdd vss bl[128] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_130 br[129] vdd vss bl[129] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_130 br[129] vdd vss bl[129] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_130 br[129] vdd vss bl[129] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_130 br[129] vdd vss bl[129] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_130 br[129] vdd vss bl[129] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_130 br[129] vdd vss bl[129] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_130 br[129] vdd vss bl[129] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_130 br[129] vdd vss bl[129] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_130 br[129] vdd vss bl[129] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_130 br[129] vdd vss bl[129] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_130 br[129] vdd vss bl[129] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_130 br[129] vdd vss bl[129] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_130 br[129] vdd vss bl[129] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_130 br[129] vdd vss bl[129] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_130 br[129] vdd vss bl[129] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_130 br[129] vdd vss bl[129] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_130 br[129] vdd vss bl[129] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_130 br[129] vdd vss bl[129] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_130 br[129] vdd vss bl[129] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_131 br[130] vdd vss bl[130] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_131 br[130] vdd vss bl[130] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_131 br[130] vdd vss bl[130] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_131 br[130] vdd vss bl[130] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_131 br[130] vdd vss bl[130] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_131 br[130] vdd vss bl[130] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_131 br[130] vdd vss bl[130] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_131 br[130] vdd vss bl[130] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_131 br[130] vdd vss bl[130] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_131 br[130] vdd vss bl[130] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_131 br[130] vdd vss bl[130] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_131 br[130] vdd vss bl[130] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_131 br[130] vdd vss bl[130] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_131 br[130] vdd vss bl[130] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_131 br[130] vdd vss bl[130] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_131 br[130] vdd vss bl[130] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_131 br[130] vdd vss bl[130] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_131 br[130] vdd vss bl[130] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_131 br[130] vdd vss bl[130] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_132 br[131] vdd vss bl[131] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_132 br[131] vdd vss bl[131] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_132 br[131] vdd vss bl[131] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_132 br[131] vdd vss bl[131] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_132 br[131] vdd vss bl[131] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_132 br[131] vdd vss bl[131] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_132 br[131] vdd vss bl[131] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_132 br[131] vdd vss bl[131] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_132 br[131] vdd vss bl[131] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_132 br[131] vdd vss bl[131] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_132 br[131] vdd vss bl[131] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_132 br[131] vdd vss bl[131] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_132 br[131] vdd vss bl[131] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_132 br[131] vdd vss bl[131] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_132 br[131] vdd vss bl[131] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_132 br[131] vdd vss bl[131] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_132 br[131] vdd vss bl[131] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_132 br[131] vdd vss bl[131] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_132 br[131] vdd vss bl[131] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_133 br[132] vdd vss bl[132] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_133 br[132] vdd vss bl[132] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_133 br[132] vdd vss bl[132] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_133 br[132] vdd vss bl[132] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_133 br[132] vdd vss bl[132] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_133 br[132] vdd vss bl[132] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_133 br[132] vdd vss bl[132] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_133 br[132] vdd vss bl[132] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_133 br[132] vdd vss bl[132] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_133 br[132] vdd vss bl[132] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_133 br[132] vdd vss bl[132] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_133 br[132] vdd vss bl[132] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_133 br[132] vdd vss bl[132] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_133 br[132] vdd vss bl[132] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_133 br[132] vdd vss bl[132] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_133 br[132] vdd vss bl[132] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_133 br[132] vdd vss bl[132] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_133 br[132] vdd vss bl[132] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_133 br[132] vdd vss bl[132] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_134 br[133] vdd vss bl[133] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_134 br[133] vdd vss bl[133] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_134 br[133] vdd vss bl[133] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_134 br[133] vdd vss bl[133] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_134 br[133] vdd vss bl[133] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_134 br[133] vdd vss bl[133] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_134 br[133] vdd vss bl[133] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_134 br[133] vdd vss bl[133] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_134 br[133] vdd vss bl[133] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_134 br[133] vdd vss bl[133] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_134 br[133] vdd vss bl[133] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_134 br[133] vdd vss bl[133] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_134 br[133] vdd vss bl[133] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_134 br[133] vdd vss bl[133] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_134 br[133] vdd vss bl[133] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_134 br[133] vdd vss bl[133] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_134 br[133] vdd vss bl[133] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_134 br[133] vdd vss bl[133] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_134 br[133] vdd vss bl[133] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_135 br[134] vdd vss bl[134] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_135 br[134] vdd vss bl[134] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_135 br[134] vdd vss bl[134] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_135 br[134] vdd vss bl[134] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_135 br[134] vdd vss bl[134] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_135 br[134] vdd vss bl[134] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_135 br[134] vdd vss bl[134] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_135 br[134] vdd vss bl[134] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_135 br[134] vdd vss bl[134] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_135 br[134] vdd vss bl[134] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_135 br[134] vdd vss bl[134] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_135 br[134] vdd vss bl[134] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_135 br[134] vdd vss bl[134] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_135 br[134] vdd vss bl[134] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_135 br[134] vdd vss bl[134] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_135 br[134] vdd vss bl[134] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_135 br[134] vdd vss bl[134] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_135 br[134] vdd vss bl[134] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_135 br[134] vdd vss bl[134] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_136 br[135] vdd vss bl[135] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_136 br[135] vdd vss bl[135] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_136 br[135] vdd vss bl[135] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_136 br[135] vdd vss bl[135] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_136 br[135] vdd vss bl[135] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_136 br[135] vdd vss bl[135] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_136 br[135] vdd vss bl[135] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_136 br[135] vdd vss bl[135] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_136 br[135] vdd vss bl[135] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_136 br[135] vdd vss bl[135] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_136 br[135] vdd vss bl[135] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_136 br[135] vdd vss bl[135] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_136 br[135] vdd vss bl[135] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_136 br[135] vdd vss bl[135] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_136 br[135] vdd vss bl[135] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_136 br[135] vdd vss bl[135] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_136 br[135] vdd vss bl[135] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_136 br[135] vdd vss bl[135] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_136 br[135] vdd vss bl[135] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_137 br[136] vdd vss bl[136] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_137 br[136] vdd vss bl[136] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_137 br[136] vdd vss bl[136] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_137 br[136] vdd vss bl[136] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_137 br[136] vdd vss bl[136] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_137 br[136] vdd vss bl[136] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_137 br[136] vdd vss bl[136] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_137 br[136] vdd vss bl[136] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_137 br[136] vdd vss bl[136] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_137 br[136] vdd vss bl[136] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_137 br[136] vdd vss bl[136] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_137 br[136] vdd vss bl[136] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_137 br[136] vdd vss bl[136] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_137 br[136] vdd vss bl[136] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_137 br[136] vdd vss bl[136] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_137 br[136] vdd vss bl[136] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_137 br[136] vdd vss bl[136] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_137 br[136] vdd vss bl[136] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_137 br[136] vdd vss bl[136] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_138 br[137] vdd vss bl[137] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_138 br[137] vdd vss bl[137] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_138 br[137] vdd vss bl[137] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_138 br[137] vdd vss bl[137] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_138 br[137] vdd vss bl[137] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_138 br[137] vdd vss bl[137] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_138 br[137] vdd vss bl[137] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_138 br[137] vdd vss bl[137] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_138 br[137] vdd vss bl[137] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_138 br[137] vdd vss bl[137] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_138 br[137] vdd vss bl[137] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_138 br[137] vdd vss bl[137] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_138 br[137] vdd vss bl[137] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_138 br[137] vdd vss bl[137] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_138 br[137] vdd vss bl[137] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_138 br[137] vdd vss bl[137] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_138 br[137] vdd vss bl[137] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_138 br[137] vdd vss bl[137] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_138 br[137] vdd vss bl[137] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_139 br[138] vdd vss bl[138] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_139 br[138] vdd vss bl[138] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_139 br[138] vdd vss bl[138] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_139 br[138] vdd vss bl[138] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_139 br[138] vdd vss bl[138] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_139 br[138] vdd vss bl[138] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_139 br[138] vdd vss bl[138] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_139 br[138] vdd vss bl[138] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_139 br[138] vdd vss bl[138] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_139 br[138] vdd vss bl[138] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_139 br[138] vdd vss bl[138] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_139 br[138] vdd vss bl[138] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_139 br[138] vdd vss bl[138] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_139 br[138] vdd vss bl[138] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_139 br[138] vdd vss bl[138] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_139 br[138] vdd vss bl[138] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_139 br[138] vdd vss bl[138] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_139 br[138] vdd vss bl[138] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_139 br[138] vdd vss bl[138] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_140 br[139] vdd vss bl[139] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_140 br[139] vdd vss bl[139] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_140 br[139] vdd vss bl[139] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_140 br[139] vdd vss bl[139] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_140 br[139] vdd vss bl[139] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_140 br[139] vdd vss bl[139] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_140 br[139] vdd vss bl[139] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_140 br[139] vdd vss bl[139] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_140 br[139] vdd vss bl[139] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_140 br[139] vdd vss bl[139] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_140 br[139] vdd vss bl[139] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_140 br[139] vdd vss bl[139] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_140 br[139] vdd vss bl[139] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_140 br[139] vdd vss bl[139] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_140 br[139] vdd vss bl[139] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_140 br[139] vdd vss bl[139] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_140 br[139] vdd vss bl[139] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_140 br[139] vdd vss bl[139] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_140 br[139] vdd vss bl[139] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_141 br[140] vdd vss bl[140] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_141 br[140] vdd vss bl[140] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_141 br[140] vdd vss bl[140] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_141 br[140] vdd vss bl[140] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_141 br[140] vdd vss bl[140] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_141 br[140] vdd vss bl[140] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_141 br[140] vdd vss bl[140] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_141 br[140] vdd vss bl[140] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_141 br[140] vdd vss bl[140] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_141 br[140] vdd vss bl[140] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_141 br[140] vdd vss bl[140] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_141 br[140] vdd vss bl[140] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_141 br[140] vdd vss bl[140] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_141 br[140] vdd vss bl[140] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_141 br[140] vdd vss bl[140] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_141 br[140] vdd vss bl[140] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_141 br[140] vdd vss bl[140] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_141 br[140] vdd vss bl[140] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_141 br[140] vdd vss bl[140] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_142 br[141] vdd vss bl[141] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_142 br[141] vdd vss bl[141] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_142 br[141] vdd vss bl[141] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_142 br[141] vdd vss bl[141] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_142 br[141] vdd vss bl[141] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_142 br[141] vdd vss bl[141] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_142 br[141] vdd vss bl[141] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_142 br[141] vdd vss bl[141] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_142 br[141] vdd vss bl[141] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_142 br[141] vdd vss bl[141] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_142 br[141] vdd vss bl[141] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_142 br[141] vdd vss bl[141] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_142 br[141] vdd vss bl[141] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_142 br[141] vdd vss bl[141] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_142 br[141] vdd vss bl[141] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_142 br[141] vdd vss bl[141] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_142 br[141] vdd vss bl[141] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_142 br[141] vdd vss bl[141] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_142 br[141] vdd vss bl[141] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_143 br[142] vdd vss bl[142] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_143 br[142] vdd vss bl[142] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_143 br[142] vdd vss bl[142] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_143 br[142] vdd vss bl[142] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_143 br[142] vdd vss bl[142] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_143 br[142] vdd vss bl[142] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_143 br[142] vdd vss bl[142] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_143 br[142] vdd vss bl[142] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_143 br[142] vdd vss bl[142] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_143 br[142] vdd vss bl[142] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_143 br[142] vdd vss bl[142] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_143 br[142] vdd vss bl[142] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_143 br[142] vdd vss bl[142] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_143 br[142] vdd vss bl[142] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_143 br[142] vdd vss bl[142] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_143 br[142] vdd vss bl[142] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_143 br[142] vdd vss bl[142] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_143 br[142] vdd vss bl[142] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_143 br[142] vdd vss bl[142] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_144 br[143] vdd vss bl[143] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_144 br[143] vdd vss bl[143] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_144 br[143] vdd vss bl[143] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_144 br[143] vdd vss bl[143] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_144 br[143] vdd vss bl[143] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_144 br[143] vdd vss bl[143] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_144 br[143] vdd vss bl[143] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_144 br[143] vdd vss bl[143] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_144 br[143] vdd vss bl[143] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_144 br[143] vdd vss bl[143] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_144 br[143] vdd vss bl[143] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_144 br[143] vdd vss bl[143] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_144 br[143] vdd vss bl[143] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_144 br[143] vdd vss bl[143] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_144 br[143] vdd vss bl[143] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_144 br[143] vdd vss bl[143] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_144 br[143] vdd vss bl[143] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_144 br[143] vdd vss bl[143] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_144 br[143] vdd vss bl[143] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_145 br[144] vdd vss bl[144] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_145 br[144] vdd vss bl[144] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_145 br[144] vdd vss bl[144] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_145 br[144] vdd vss bl[144] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_145 br[144] vdd vss bl[144] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_145 br[144] vdd vss bl[144] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_145 br[144] vdd vss bl[144] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_145 br[144] vdd vss bl[144] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_145 br[144] vdd vss bl[144] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_145 br[144] vdd vss bl[144] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_145 br[144] vdd vss bl[144] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_145 br[144] vdd vss bl[144] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_145 br[144] vdd vss bl[144] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_145 br[144] vdd vss bl[144] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_145 br[144] vdd vss bl[144] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_145 br[144] vdd vss bl[144] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_145 br[144] vdd vss bl[144] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_145 br[144] vdd vss bl[144] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_145 br[144] vdd vss bl[144] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_146 br[145] vdd vss bl[145] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_146 br[145] vdd vss bl[145] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_146 br[145] vdd vss bl[145] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_146 br[145] vdd vss bl[145] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_146 br[145] vdd vss bl[145] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_146 br[145] vdd vss bl[145] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_146 br[145] vdd vss bl[145] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_146 br[145] vdd vss bl[145] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_146 br[145] vdd vss bl[145] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_146 br[145] vdd vss bl[145] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_146 br[145] vdd vss bl[145] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_146 br[145] vdd vss bl[145] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_146 br[145] vdd vss bl[145] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_146 br[145] vdd vss bl[145] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_146 br[145] vdd vss bl[145] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_146 br[145] vdd vss bl[145] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_146 br[145] vdd vss bl[145] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_146 br[145] vdd vss bl[145] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_146 br[145] vdd vss bl[145] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_147 br[146] vdd vss bl[146] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_147 br[146] vdd vss bl[146] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_147 br[146] vdd vss bl[146] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_147 br[146] vdd vss bl[146] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_147 br[146] vdd vss bl[146] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_147 br[146] vdd vss bl[146] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_147 br[146] vdd vss bl[146] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_147 br[146] vdd vss bl[146] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_147 br[146] vdd vss bl[146] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_147 br[146] vdd vss bl[146] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_147 br[146] vdd vss bl[146] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_147 br[146] vdd vss bl[146] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_147 br[146] vdd vss bl[146] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_147 br[146] vdd vss bl[146] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_147 br[146] vdd vss bl[146] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_147 br[146] vdd vss bl[146] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_147 br[146] vdd vss bl[146] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_147 br[146] vdd vss bl[146] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_147 br[146] vdd vss bl[146] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_148 br[147] vdd vss bl[147] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_148 br[147] vdd vss bl[147] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_148 br[147] vdd vss bl[147] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_148 br[147] vdd vss bl[147] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_148 br[147] vdd vss bl[147] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_148 br[147] vdd vss bl[147] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_148 br[147] vdd vss bl[147] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_148 br[147] vdd vss bl[147] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_148 br[147] vdd vss bl[147] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_148 br[147] vdd vss bl[147] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_148 br[147] vdd vss bl[147] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_148 br[147] vdd vss bl[147] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_148 br[147] vdd vss bl[147] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_148 br[147] vdd vss bl[147] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_148 br[147] vdd vss bl[147] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_148 br[147] vdd vss bl[147] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_148 br[147] vdd vss bl[147] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_148 br[147] vdd vss bl[147] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_148 br[147] vdd vss bl[147] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_149 br[148] vdd vss bl[148] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_149 br[148] vdd vss bl[148] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_149 br[148] vdd vss bl[148] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_149 br[148] vdd vss bl[148] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_149 br[148] vdd vss bl[148] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_149 br[148] vdd vss bl[148] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_149 br[148] vdd vss bl[148] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_149 br[148] vdd vss bl[148] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_149 br[148] vdd vss bl[148] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_149 br[148] vdd vss bl[148] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_149 br[148] vdd vss bl[148] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_149 br[148] vdd vss bl[148] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_149 br[148] vdd vss bl[148] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_149 br[148] vdd vss bl[148] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_149 br[148] vdd vss bl[148] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_149 br[148] vdd vss bl[148] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_149 br[148] vdd vss bl[148] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_149 br[148] vdd vss bl[148] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_149 br[148] vdd vss bl[148] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_150 br[149] vdd vss bl[149] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_150 br[149] vdd vss bl[149] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_150 br[149] vdd vss bl[149] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_150 br[149] vdd vss bl[149] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_150 br[149] vdd vss bl[149] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_150 br[149] vdd vss bl[149] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_150 br[149] vdd vss bl[149] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_150 br[149] vdd vss bl[149] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_150 br[149] vdd vss bl[149] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_150 br[149] vdd vss bl[149] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_150 br[149] vdd vss bl[149] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_150 br[149] vdd vss bl[149] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_150 br[149] vdd vss bl[149] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_150 br[149] vdd vss bl[149] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_150 br[149] vdd vss bl[149] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_150 br[149] vdd vss bl[149] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_150 br[149] vdd vss bl[149] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_150 br[149] vdd vss bl[149] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_150 br[149] vdd vss bl[149] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_151 br[150] vdd vss bl[150] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_151 br[150] vdd vss bl[150] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_151 br[150] vdd vss bl[150] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_151 br[150] vdd vss bl[150] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_151 br[150] vdd vss bl[150] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_151 br[150] vdd vss bl[150] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_151 br[150] vdd vss bl[150] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_151 br[150] vdd vss bl[150] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_151 br[150] vdd vss bl[150] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_151 br[150] vdd vss bl[150] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_151 br[150] vdd vss bl[150] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_151 br[150] vdd vss bl[150] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_151 br[150] vdd vss bl[150] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_151 br[150] vdd vss bl[150] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_151 br[150] vdd vss bl[150] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_151 br[150] vdd vss bl[150] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_151 br[150] vdd vss bl[150] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_151 br[150] vdd vss bl[150] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_151 br[150] vdd vss bl[150] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_152 br[151] vdd vss bl[151] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_152 br[151] vdd vss bl[151] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_152 br[151] vdd vss bl[151] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_152 br[151] vdd vss bl[151] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_152 br[151] vdd vss bl[151] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_152 br[151] vdd vss bl[151] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_152 br[151] vdd vss bl[151] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_152 br[151] vdd vss bl[151] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_152 br[151] vdd vss bl[151] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_152 br[151] vdd vss bl[151] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_152 br[151] vdd vss bl[151] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_152 br[151] vdd vss bl[151] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_152 br[151] vdd vss bl[151] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_152 br[151] vdd vss bl[151] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_152 br[151] vdd vss bl[151] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_152 br[151] vdd vss bl[151] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_152 br[151] vdd vss bl[151] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_152 br[151] vdd vss bl[151] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_152 br[151] vdd vss bl[151] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_153 br[152] vdd vss bl[152] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_153 br[152] vdd vss bl[152] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_153 br[152] vdd vss bl[152] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_153 br[152] vdd vss bl[152] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_153 br[152] vdd vss bl[152] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_153 br[152] vdd vss bl[152] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_153 br[152] vdd vss bl[152] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_153 br[152] vdd vss bl[152] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_153 br[152] vdd vss bl[152] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_153 br[152] vdd vss bl[152] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_153 br[152] vdd vss bl[152] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_153 br[152] vdd vss bl[152] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_153 br[152] vdd vss bl[152] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_153 br[152] vdd vss bl[152] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_153 br[152] vdd vss bl[152] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_153 br[152] vdd vss bl[152] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_153 br[152] vdd vss bl[152] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_153 br[152] vdd vss bl[152] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_153 br[152] vdd vss bl[152] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_154 br[153] vdd vss bl[153] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_154 br[153] vdd vss bl[153] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_154 br[153] vdd vss bl[153] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_154 br[153] vdd vss bl[153] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_154 br[153] vdd vss bl[153] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_154 br[153] vdd vss bl[153] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_154 br[153] vdd vss bl[153] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_154 br[153] vdd vss bl[153] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_154 br[153] vdd vss bl[153] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_154 br[153] vdd vss bl[153] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_154 br[153] vdd vss bl[153] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_154 br[153] vdd vss bl[153] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_154 br[153] vdd vss bl[153] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_154 br[153] vdd vss bl[153] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_154 br[153] vdd vss bl[153] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_154 br[153] vdd vss bl[153] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_154 br[153] vdd vss bl[153] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_154 br[153] vdd vss bl[153] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_154 br[153] vdd vss bl[153] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_155 br[154] vdd vss bl[154] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_155 br[154] vdd vss bl[154] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_155 br[154] vdd vss bl[154] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_155 br[154] vdd vss bl[154] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_155 br[154] vdd vss bl[154] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_155 br[154] vdd vss bl[154] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_155 br[154] vdd vss bl[154] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_155 br[154] vdd vss bl[154] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_155 br[154] vdd vss bl[154] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_155 br[154] vdd vss bl[154] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_155 br[154] vdd vss bl[154] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_155 br[154] vdd vss bl[154] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_155 br[154] vdd vss bl[154] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_155 br[154] vdd vss bl[154] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_155 br[154] vdd vss bl[154] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_155 br[154] vdd vss bl[154] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_155 br[154] vdd vss bl[154] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_155 br[154] vdd vss bl[154] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_155 br[154] vdd vss bl[154] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_156 br[155] vdd vss bl[155] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_156 br[155] vdd vss bl[155] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_156 br[155] vdd vss bl[155] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_156 br[155] vdd vss bl[155] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_156 br[155] vdd vss bl[155] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_156 br[155] vdd vss bl[155] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_156 br[155] vdd vss bl[155] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_156 br[155] vdd vss bl[155] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_156 br[155] vdd vss bl[155] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_156 br[155] vdd vss bl[155] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_156 br[155] vdd vss bl[155] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_156 br[155] vdd vss bl[155] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_156 br[155] vdd vss bl[155] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_156 br[155] vdd vss bl[155] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_156 br[155] vdd vss bl[155] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_156 br[155] vdd vss bl[155] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_156 br[155] vdd vss bl[155] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_156 br[155] vdd vss bl[155] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_156 br[155] vdd vss bl[155] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_157 br[156] vdd vss bl[156] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_157 br[156] vdd vss bl[156] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_157 br[156] vdd vss bl[156] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_157 br[156] vdd vss bl[156] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_157 br[156] vdd vss bl[156] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_157 br[156] vdd vss bl[156] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_157 br[156] vdd vss bl[156] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_157 br[156] vdd vss bl[156] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_157 br[156] vdd vss bl[156] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_157 br[156] vdd vss bl[156] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_157 br[156] vdd vss bl[156] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_157 br[156] vdd vss bl[156] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_157 br[156] vdd vss bl[156] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_157 br[156] vdd vss bl[156] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_157 br[156] vdd vss bl[156] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_157 br[156] vdd vss bl[156] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_157 br[156] vdd vss bl[156] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_157 br[156] vdd vss bl[156] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_157 br[156] vdd vss bl[156] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_158 br[157] vdd vss bl[157] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_158 br[157] vdd vss bl[157] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_158 br[157] vdd vss bl[157] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_158 br[157] vdd vss bl[157] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_158 br[157] vdd vss bl[157] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_158 br[157] vdd vss bl[157] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_158 br[157] vdd vss bl[157] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_158 br[157] vdd vss bl[157] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_158 br[157] vdd vss bl[157] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_158 br[157] vdd vss bl[157] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_158 br[157] vdd vss bl[157] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_158 br[157] vdd vss bl[157] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_158 br[157] vdd vss bl[157] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_158 br[157] vdd vss bl[157] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_158 br[157] vdd vss bl[157] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_158 br[157] vdd vss bl[157] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_158 br[157] vdd vss bl[157] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_158 br[157] vdd vss bl[157] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_158 br[157] vdd vss bl[157] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_159 br[158] vdd vss bl[158] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_159 br[158] vdd vss bl[158] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_159 br[158] vdd vss bl[158] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_159 br[158] vdd vss bl[158] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_159 br[158] vdd vss bl[158] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_159 br[158] vdd vss bl[158] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_159 br[158] vdd vss bl[158] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_159 br[158] vdd vss bl[158] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_159 br[158] vdd vss bl[158] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_159 br[158] vdd vss bl[158] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_159 br[158] vdd vss bl[158] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_159 br[158] vdd vss bl[158] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_159 br[158] vdd vss bl[158] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_159 br[158] vdd vss bl[158] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_159 br[158] vdd vss bl[158] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_159 br[158] vdd vss bl[158] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_159 br[158] vdd vss bl[158] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_159 br[158] vdd vss bl[158] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_159 br[158] vdd vss bl[158] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_160 br[159] vdd vss bl[159] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_160 br[159] vdd vss bl[159] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_160 br[159] vdd vss bl[159] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_160 br[159] vdd vss bl[159] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_160 br[159] vdd vss bl[159] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_160 br[159] vdd vss bl[159] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_160 br[159] vdd vss bl[159] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_160 br[159] vdd vss bl[159] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_160 br[159] vdd vss bl[159] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_160 br[159] vdd vss bl[159] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_160 br[159] vdd vss bl[159] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_160 br[159] vdd vss bl[159] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_160 br[159] vdd vss bl[159] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_160 br[159] vdd vss bl[159] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_160 br[159] vdd vss bl[159] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_160 br[159] vdd vss bl[159] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_160 br[159] vdd vss bl[159] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_160 br[159] vdd vss bl[159] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_160 br[159] vdd vss bl[159] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_161 br[160] vdd vss bl[160] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_161 br[160] vdd vss bl[160] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_161 br[160] vdd vss bl[160] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_161 br[160] vdd vss bl[160] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_161 br[160] vdd vss bl[160] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_161 br[160] vdd vss bl[160] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_161 br[160] vdd vss bl[160] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_161 br[160] vdd vss bl[160] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_161 br[160] vdd vss bl[160] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_161 br[160] vdd vss bl[160] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_161 br[160] vdd vss bl[160] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_161 br[160] vdd vss bl[160] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_161 br[160] vdd vss bl[160] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_161 br[160] vdd vss bl[160] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_161 br[160] vdd vss bl[160] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_161 br[160] vdd vss bl[160] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_161 br[160] vdd vss bl[160] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_161 br[160] vdd vss bl[160] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_161 br[160] vdd vss bl[160] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_162 br[161] vdd vss bl[161] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_162 br[161] vdd vss bl[161] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_162 br[161] vdd vss bl[161] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_162 br[161] vdd vss bl[161] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_162 br[161] vdd vss bl[161] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_162 br[161] vdd vss bl[161] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_162 br[161] vdd vss bl[161] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_162 br[161] vdd vss bl[161] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_162 br[161] vdd vss bl[161] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_162 br[161] vdd vss bl[161] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_162 br[161] vdd vss bl[161] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_162 br[161] vdd vss bl[161] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_162 br[161] vdd vss bl[161] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_162 br[161] vdd vss bl[161] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_162 br[161] vdd vss bl[161] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_162 br[161] vdd vss bl[161] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_162 br[161] vdd vss bl[161] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_162 br[161] vdd vss bl[161] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_162 br[161] vdd vss bl[161] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_163 br[162] vdd vss bl[162] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_163 br[162] vdd vss bl[162] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_163 br[162] vdd vss bl[162] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_163 br[162] vdd vss bl[162] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_163 br[162] vdd vss bl[162] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_163 br[162] vdd vss bl[162] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_163 br[162] vdd vss bl[162] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_163 br[162] vdd vss bl[162] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_163 br[162] vdd vss bl[162] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_163 br[162] vdd vss bl[162] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_163 br[162] vdd vss bl[162] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_163 br[162] vdd vss bl[162] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_163 br[162] vdd vss bl[162] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_163 br[162] vdd vss bl[162] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_163 br[162] vdd vss bl[162] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_163 br[162] vdd vss bl[162] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_163 br[162] vdd vss bl[162] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_163 br[162] vdd vss bl[162] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_163 br[162] vdd vss bl[162] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_164 br[163] vdd vss bl[163] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_164 br[163] vdd vss bl[163] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_164 br[163] vdd vss bl[163] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_164 br[163] vdd vss bl[163] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_164 br[163] vdd vss bl[163] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_164 br[163] vdd vss bl[163] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_164 br[163] vdd vss bl[163] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_164 br[163] vdd vss bl[163] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_164 br[163] vdd vss bl[163] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_164 br[163] vdd vss bl[163] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_164 br[163] vdd vss bl[163] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_164 br[163] vdd vss bl[163] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_164 br[163] vdd vss bl[163] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_164 br[163] vdd vss bl[163] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_164 br[163] vdd vss bl[163] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_164 br[163] vdd vss bl[163] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_164 br[163] vdd vss bl[163] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_164 br[163] vdd vss bl[163] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_164 br[163] vdd vss bl[163] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_165 br[164] vdd vss bl[164] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_165 br[164] vdd vss bl[164] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_165 br[164] vdd vss bl[164] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_165 br[164] vdd vss bl[164] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_165 br[164] vdd vss bl[164] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_165 br[164] vdd vss bl[164] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_165 br[164] vdd vss bl[164] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_165 br[164] vdd vss bl[164] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_165 br[164] vdd vss bl[164] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_165 br[164] vdd vss bl[164] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_165 br[164] vdd vss bl[164] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_165 br[164] vdd vss bl[164] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_165 br[164] vdd vss bl[164] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_165 br[164] vdd vss bl[164] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_165 br[164] vdd vss bl[164] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_165 br[164] vdd vss bl[164] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_165 br[164] vdd vss bl[164] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_165 br[164] vdd vss bl[164] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_165 br[164] vdd vss bl[164] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_166 br[165] vdd vss bl[165] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_166 br[165] vdd vss bl[165] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_166 br[165] vdd vss bl[165] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_166 br[165] vdd vss bl[165] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_166 br[165] vdd vss bl[165] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_166 br[165] vdd vss bl[165] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_166 br[165] vdd vss bl[165] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_166 br[165] vdd vss bl[165] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_166 br[165] vdd vss bl[165] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_166 br[165] vdd vss bl[165] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_166 br[165] vdd vss bl[165] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_166 br[165] vdd vss bl[165] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_166 br[165] vdd vss bl[165] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_166 br[165] vdd vss bl[165] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_166 br[165] vdd vss bl[165] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_166 br[165] vdd vss bl[165] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_166 br[165] vdd vss bl[165] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_166 br[165] vdd vss bl[165] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_166 br[165] vdd vss bl[165] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_167 br[166] vdd vss bl[166] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_167 br[166] vdd vss bl[166] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_167 br[166] vdd vss bl[166] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_167 br[166] vdd vss bl[166] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_167 br[166] vdd vss bl[166] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_167 br[166] vdd vss bl[166] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_167 br[166] vdd vss bl[166] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_167 br[166] vdd vss bl[166] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_167 br[166] vdd vss bl[166] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_167 br[166] vdd vss bl[166] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_167 br[166] vdd vss bl[166] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_167 br[166] vdd vss bl[166] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_167 br[166] vdd vss bl[166] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_167 br[166] vdd vss bl[166] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_167 br[166] vdd vss bl[166] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_167 br[166] vdd vss bl[166] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_167 br[166] vdd vss bl[166] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_167 br[166] vdd vss bl[166] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_167 br[166] vdd vss bl[166] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_168 br[167] vdd vss bl[167] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_168 br[167] vdd vss bl[167] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_168 br[167] vdd vss bl[167] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_168 br[167] vdd vss bl[167] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_168 br[167] vdd vss bl[167] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_168 br[167] vdd vss bl[167] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_168 br[167] vdd vss bl[167] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_168 br[167] vdd vss bl[167] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_168 br[167] vdd vss bl[167] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_168 br[167] vdd vss bl[167] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_168 br[167] vdd vss bl[167] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_168 br[167] vdd vss bl[167] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_168 br[167] vdd vss bl[167] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_168 br[167] vdd vss bl[167] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_168 br[167] vdd vss bl[167] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_168 br[167] vdd vss bl[167] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_168 br[167] vdd vss bl[167] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_168 br[167] vdd vss bl[167] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_168 br[167] vdd vss bl[167] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_169 br[168] vdd vss bl[168] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_169 br[168] vdd vss bl[168] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_169 br[168] vdd vss bl[168] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_169 br[168] vdd vss bl[168] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_169 br[168] vdd vss bl[168] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_169 br[168] vdd vss bl[168] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_169 br[168] vdd vss bl[168] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_169 br[168] vdd vss bl[168] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_169 br[168] vdd vss bl[168] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_169 br[168] vdd vss bl[168] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_169 br[168] vdd vss bl[168] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_169 br[168] vdd vss bl[168] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_169 br[168] vdd vss bl[168] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_169 br[168] vdd vss bl[168] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_169 br[168] vdd vss bl[168] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_169 br[168] vdd vss bl[168] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_169 br[168] vdd vss bl[168] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_169 br[168] vdd vss bl[168] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_169 br[168] vdd vss bl[168] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_170 br[169] vdd vss bl[169] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_170 br[169] vdd vss bl[169] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_170 br[169] vdd vss bl[169] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_170 br[169] vdd vss bl[169] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_170 br[169] vdd vss bl[169] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_170 br[169] vdd vss bl[169] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_170 br[169] vdd vss bl[169] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_170 br[169] vdd vss bl[169] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_170 br[169] vdd vss bl[169] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_170 br[169] vdd vss bl[169] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_170 br[169] vdd vss bl[169] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_170 br[169] vdd vss bl[169] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_170 br[169] vdd vss bl[169] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_170 br[169] vdd vss bl[169] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_170 br[169] vdd vss bl[169] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_170 br[169] vdd vss bl[169] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_170 br[169] vdd vss bl[169] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_170 br[169] vdd vss bl[169] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_170 br[169] vdd vss bl[169] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_171 br[170] vdd vss bl[170] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_171 br[170] vdd vss bl[170] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_171 br[170] vdd vss bl[170] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_171 br[170] vdd vss bl[170] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_171 br[170] vdd vss bl[170] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_171 br[170] vdd vss bl[170] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_171 br[170] vdd vss bl[170] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_171 br[170] vdd vss bl[170] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_171 br[170] vdd vss bl[170] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_171 br[170] vdd vss bl[170] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_171 br[170] vdd vss bl[170] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_171 br[170] vdd vss bl[170] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_171 br[170] vdd vss bl[170] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_171 br[170] vdd vss bl[170] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_171 br[170] vdd vss bl[170] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_171 br[170] vdd vss bl[170] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_171 br[170] vdd vss bl[170] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_171 br[170] vdd vss bl[170] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_171 br[170] vdd vss bl[170] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_172 br[171] vdd vss bl[171] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_172 br[171] vdd vss bl[171] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_172 br[171] vdd vss bl[171] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_172 br[171] vdd vss bl[171] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_172 br[171] vdd vss bl[171] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_172 br[171] vdd vss bl[171] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_172 br[171] vdd vss bl[171] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_172 br[171] vdd vss bl[171] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_172 br[171] vdd vss bl[171] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_172 br[171] vdd vss bl[171] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_172 br[171] vdd vss bl[171] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_172 br[171] vdd vss bl[171] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_172 br[171] vdd vss bl[171] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_172 br[171] vdd vss bl[171] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_172 br[171] vdd vss bl[171] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_172 br[171] vdd vss bl[171] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_172 br[171] vdd vss bl[171] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_172 br[171] vdd vss bl[171] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_172 br[171] vdd vss bl[171] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_173 br[172] vdd vss bl[172] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_173 br[172] vdd vss bl[172] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_173 br[172] vdd vss bl[172] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_173 br[172] vdd vss bl[172] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_173 br[172] vdd vss bl[172] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_173 br[172] vdd vss bl[172] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_173 br[172] vdd vss bl[172] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_173 br[172] vdd vss bl[172] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_173 br[172] vdd vss bl[172] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_173 br[172] vdd vss bl[172] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_173 br[172] vdd vss bl[172] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_173 br[172] vdd vss bl[172] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_173 br[172] vdd vss bl[172] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_173 br[172] vdd vss bl[172] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_173 br[172] vdd vss bl[172] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_173 br[172] vdd vss bl[172] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_173 br[172] vdd vss bl[172] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_173 br[172] vdd vss bl[172] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_173 br[172] vdd vss bl[172] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_174 br[173] vdd vss bl[173] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_174 br[173] vdd vss bl[173] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_174 br[173] vdd vss bl[173] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_174 br[173] vdd vss bl[173] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_174 br[173] vdd vss bl[173] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_174 br[173] vdd vss bl[173] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_174 br[173] vdd vss bl[173] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_174 br[173] vdd vss bl[173] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_174 br[173] vdd vss bl[173] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_174 br[173] vdd vss bl[173] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_174 br[173] vdd vss bl[173] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_174 br[173] vdd vss bl[173] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_174 br[173] vdd vss bl[173] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_174 br[173] vdd vss bl[173] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_174 br[173] vdd vss bl[173] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_174 br[173] vdd vss bl[173] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_174 br[173] vdd vss bl[173] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_174 br[173] vdd vss bl[173] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_174 br[173] vdd vss bl[173] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_175 br[174] vdd vss bl[174] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_175 br[174] vdd vss bl[174] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_175 br[174] vdd vss bl[174] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_175 br[174] vdd vss bl[174] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_175 br[174] vdd vss bl[174] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_175 br[174] vdd vss bl[174] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_175 br[174] vdd vss bl[174] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_175 br[174] vdd vss bl[174] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_175 br[174] vdd vss bl[174] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_175 br[174] vdd vss bl[174] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_175 br[174] vdd vss bl[174] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_175 br[174] vdd vss bl[174] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_175 br[174] vdd vss bl[174] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_175 br[174] vdd vss bl[174] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_175 br[174] vdd vss bl[174] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_175 br[174] vdd vss bl[174] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_175 br[174] vdd vss bl[174] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_175 br[174] vdd vss bl[174] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_175 br[174] vdd vss bl[174] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_176 br[175] vdd vss bl[175] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_176 br[175] vdd vss bl[175] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_176 br[175] vdd vss bl[175] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_176 br[175] vdd vss bl[175] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_176 br[175] vdd vss bl[175] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_176 br[175] vdd vss bl[175] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_176 br[175] vdd vss bl[175] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_176 br[175] vdd vss bl[175] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_176 br[175] vdd vss bl[175] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_176 br[175] vdd vss bl[175] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_176 br[175] vdd vss bl[175] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_176 br[175] vdd vss bl[175] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_176 br[175] vdd vss bl[175] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_176 br[175] vdd vss bl[175] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_176 br[175] vdd vss bl[175] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_176 br[175] vdd vss bl[175] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_176 br[175] vdd vss bl[175] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_176 br[175] vdd vss bl[175] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_176 br[175] vdd vss bl[175] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_177 br[176] vdd vss bl[176] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_177 br[176] vdd vss bl[176] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_177 br[176] vdd vss bl[176] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_177 br[176] vdd vss bl[176] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_177 br[176] vdd vss bl[176] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_177 br[176] vdd vss bl[176] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_177 br[176] vdd vss bl[176] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_177 br[176] vdd vss bl[176] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_177 br[176] vdd vss bl[176] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_177 br[176] vdd vss bl[176] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_177 br[176] vdd vss bl[176] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_177 br[176] vdd vss bl[176] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_177 br[176] vdd vss bl[176] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_177 br[176] vdd vss bl[176] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_177 br[176] vdd vss bl[176] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_177 br[176] vdd vss bl[176] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_177 br[176] vdd vss bl[176] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_177 br[176] vdd vss bl[176] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_177 br[176] vdd vss bl[176] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_178 br[177] vdd vss bl[177] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_178 br[177] vdd vss bl[177] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_178 br[177] vdd vss bl[177] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_178 br[177] vdd vss bl[177] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_178 br[177] vdd vss bl[177] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_178 br[177] vdd vss bl[177] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_178 br[177] vdd vss bl[177] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_178 br[177] vdd vss bl[177] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_178 br[177] vdd vss bl[177] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_178 br[177] vdd vss bl[177] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_178 br[177] vdd vss bl[177] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_178 br[177] vdd vss bl[177] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_178 br[177] vdd vss bl[177] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_178 br[177] vdd vss bl[177] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_178 br[177] vdd vss bl[177] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_178 br[177] vdd vss bl[177] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_178 br[177] vdd vss bl[177] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_178 br[177] vdd vss bl[177] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_178 br[177] vdd vss bl[177] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_179 br[178] vdd vss bl[178] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_179 br[178] vdd vss bl[178] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_179 br[178] vdd vss bl[178] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_179 br[178] vdd vss bl[178] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_179 br[178] vdd vss bl[178] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_179 br[178] vdd vss bl[178] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_179 br[178] vdd vss bl[178] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_179 br[178] vdd vss bl[178] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_179 br[178] vdd vss bl[178] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_179 br[178] vdd vss bl[178] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_179 br[178] vdd vss bl[178] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_179 br[178] vdd vss bl[178] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_179 br[178] vdd vss bl[178] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_179 br[178] vdd vss bl[178] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_179 br[178] vdd vss bl[178] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_179 br[178] vdd vss bl[178] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_179 br[178] vdd vss bl[178] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_179 br[178] vdd vss bl[178] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_179 br[178] vdd vss bl[178] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_180 br[179] vdd vss bl[179] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_180 br[179] vdd vss bl[179] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_180 br[179] vdd vss bl[179] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_180 br[179] vdd vss bl[179] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_180 br[179] vdd vss bl[179] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_180 br[179] vdd vss bl[179] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_180 br[179] vdd vss bl[179] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_180 br[179] vdd vss bl[179] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_180 br[179] vdd vss bl[179] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_180 br[179] vdd vss bl[179] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_180 br[179] vdd vss bl[179] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_180 br[179] vdd vss bl[179] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_180 br[179] vdd vss bl[179] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_180 br[179] vdd vss bl[179] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_180 br[179] vdd vss bl[179] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_180 br[179] vdd vss bl[179] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_180 br[179] vdd vss bl[179] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_180 br[179] vdd vss bl[179] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_180 br[179] vdd vss bl[179] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_181 br[180] vdd vss bl[180] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_181 br[180] vdd vss bl[180] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_181 br[180] vdd vss bl[180] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_181 br[180] vdd vss bl[180] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_181 br[180] vdd vss bl[180] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_181 br[180] vdd vss bl[180] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_181 br[180] vdd vss bl[180] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_181 br[180] vdd vss bl[180] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_181 br[180] vdd vss bl[180] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_181 br[180] vdd vss bl[180] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_181 br[180] vdd vss bl[180] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_181 br[180] vdd vss bl[180] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_181 br[180] vdd vss bl[180] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_181 br[180] vdd vss bl[180] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_181 br[180] vdd vss bl[180] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_181 br[180] vdd vss bl[180] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_181 br[180] vdd vss bl[180] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_181 br[180] vdd vss bl[180] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_181 br[180] vdd vss bl[180] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_182 br[181] vdd vss bl[181] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_182 br[181] vdd vss bl[181] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_182 br[181] vdd vss bl[181] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_182 br[181] vdd vss bl[181] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_182 br[181] vdd vss bl[181] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_182 br[181] vdd vss bl[181] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_182 br[181] vdd vss bl[181] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_182 br[181] vdd vss bl[181] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_182 br[181] vdd vss bl[181] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_182 br[181] vdd vss bl[181] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_182 br[181] vdd vss bl[181] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_182 br[181] vdd vss bl[181] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_182 br[181] vdd vss bl[181] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_182 br[181] vdd vss bl[181] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_182 br[181] vdd vss bl[181] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_182 br[181] vdd vss bl[181] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_182 br[181] vdd vss bl[181] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_182 br[181] vdd vss bl[181] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_182 br[181] vdd vss bl[181] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_183 br[182] vdd vss bl[182] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_183 br[182] vdd vss bl[182] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_183 br[182] vdd vss bl[182] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_183 br[182] vdd vss bl[182] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_183 br[182] vdd vss bl[182] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_183 br[182] vdd vss bl[182] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_183 br[182] vdd vss bl[182] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_183 br[182] vdd vss bl[182] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_183 br[182] vdd vss bl[182] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_183 br[182] vdd vss bl[182] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_183 br[182] vdd vss bl[182] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_183 br[182] vdd vss bl[182] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_183 br[182] vdd vss bl[182] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_183 br[182] vdd vss bl[182] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_183 br[182] vdd vss bl[182] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_183 br[182] vdd vss bl[182] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_183 br[182] vdd vss bl[182] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_183 br[182] vdd vss bl[182] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_183 br[182] vdd vss bl[182] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_184 br[183] vdd vss bl[183] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_184 br[183] vdd vss bl[183] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_184 br[183] vdd vss bl[183] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_184 br[183] vdd vss bl[183] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_184 br[183] vdd vss bl[183] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_184 br[183] vdd vss bl[183] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_184 br[183] vdd vss bl[183] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_184 br[183] vdd vss bl[183] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_184 br[183] vdd vss bl[183] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_184 br[183] vdd vss bl[183] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_184 br[183] vdd vss bl[183] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_184 br[183] vdd vss bl[183] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_184 br[183] vdd vss bl[183] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_184 br[183] vdd vss bl[183] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_184 br[183] vdd vss bl[183] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_184 br[183] vdd vss bl[183] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_184 br[183] vdd vss bl[183] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_184 br[183] vdd vss bl[183] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_184 br[183] vdd vss bl[183] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_185 br[184] vdd vss bl[184] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_185 br[184] vdd vss bl[184] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_185 br[184] vdd vss bl[184] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_185 br[184] vdd vss bl[184] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_185 br[184] vdd vss bl[184] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_185 br[184] vdd vss bl[184] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_185 br[184] vdd vss bl[184] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_185 br[184] vdd vss bl[184] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_185 br[184] vdd vss bl[184] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_185 br[184] vdd vss bl[184] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_185 br[184] vdd vss bl[184] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_185 br[184] vdd vss bl[184] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_185 br[184] vdd vss bl[184] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_185 br[184] vdd vss bl[184] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_185 br[184] vdd vss bl[184] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_185 br[184] vdd vss bl[184] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_185 br[184] vdd vss bl[184] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_185 br[184] vdd vss bl[184] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_185 br[184] vdd vss bl[184] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_186 br[185] vdd vss bl[185] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_186 br[185] vdd vss bl[185] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_186 br[185] vdd vss bl[185] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_186 br[185] vdd vss bl[185] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_186 br[185] vdd vss bl[185] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_186 br[185] vdd vss bl[185] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_186 br[185] vdd vss bl[185] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_186 br[185] vdd vss bl[185] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_186 br[185] vdd vss bl[185] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_186 br[185] vdd vss bl[185] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_186 br[185] vdd vss bl[185] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_186 br[185] vdd vss bl[185] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_186 br[185] vdd vss bl[185] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_186 br[185] vdd vss bl[185] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_186 br[185] vdd vss bl[185] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_186 br[185] vdd vss bl[185] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_186 br[185] vdd vss bl[185] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_186 br[185] vdd vss bl[185] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_186 br[185] vdd vss bl[185] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_187 br[186] vdd vss bl[186] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_187 br[186] vdd vss bl[186] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_187 br[186] vdd vss bl[186] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_187 br[186] vdd vss bl[186] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_187 br[186] vdd vss bl[186] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_187 br[186] vdd vss bl[186] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_187 br[186] vdd vss bl[186] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_187 br[186] vdd vss bl[186] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_187 br[186] vdd vss bl[186] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_187 br[186] vdd vss bl[186] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_187 br[186] vdd vss bl[186] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_187 br[186] vdd vss bl[186] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_187 br[186] vdd vss bl[186] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_187 br[186] vdd vss bl[186] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_187 br[186] vdd vss bl[186] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_187 br[186] vdd vss bl[186] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_187 br[186] vdd vss bl[186] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_187 br[186] vdd vss bl[186] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_187 br[186] vdd vss bl[186] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_188 br[187] vdd vss bl[187] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_188 br[187] vdd vss bl[187] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_188 br[187] vdd vss bl[187] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_188 br[187] vdd vss bl[187] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_188 br[187] vdd vss bl[187] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_188 br[187] vdd vss bl[187] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_188 br[187] vdd vss bl[187] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_188 br[187] vdd vss bl[187] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_188 br[187] vdd vss bl[187] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_188 br[187] vdd vss bl[187] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_188 br[187] vdd vss bl[187] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_188 br[187] vdd vss bl[187] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_188 br[187] vdd vss bl[187] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_188 br[187] vdd vss bl[187] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_188 br[187] vdd vss bl[187] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_188 br[187] vdd vss bl[187] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_188 br[187] vdd vss bl[187] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_188 br[187] vdd vss bl[187] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_188 br[187] vdd vss bl[187] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_189 br[188] vdd vss bl[188] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_189 br[188] vdd vss bl[188] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_189 br[188] vdd vss bl[188] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_189 br[188] vdd vss bl[188] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_189 br[188] vdd vss bl[188] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_189 br[188] vdd vss bl[188] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_189 br[188] vdd vss bl[188] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_189 br[188] vdd vss bl[188] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_189 br[188] vdd vss bl[188] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_189 br[188] vdd vss bl[188] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_189 br[188] vdd vss bl[188] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_189 br[188] vdd vss bl[188] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_189 br[188] vdd vss bl[188] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_189 br[188] vdd vss bl[188] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_189 br[188] vdd vss bl[188] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_189 br[188] vdd vss bl[188] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_189 br[188] vdd vss bl[188] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_189 br[188] vdd vss bl[188] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_189 br[188] vdd vss bl[188] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_190 br[189] vdd vss bl[189] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_190 br[189] vdd vss bl[189] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_190 br[189] vdd vss bl[189] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_190 br[189] vdd vss bl[189] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_190 br[189] vdd vss bl[189] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_190 br[189] vdd vss bl[189] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_190 br[189] vdd vss bl[189] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_190 br[189] vdd vss bl[189] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_190 br[189] vdd vss bl[189] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_190 br[189] vdd vss bl[189] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_190 br[189] vdd vss bl[189] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_190 br[189] vdd vss bl[189] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_190 br[189] vdd vss bl[189] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_190 br[189] vdd vss bl[189] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_190 br[189] vdd vss bl[189] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_190 br[189] vdd vss bl[189] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_190 br[189] vdd vss bl[189] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_190 br[189] vdd vss bl[189] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_190 br[189] vdd vss bl[189] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_191 br[190] vdd vss bl[190] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_191 br[190] vdd vss bl[190] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_191 br[190] vdd vss bl[190] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_191 br[190] vdd vss bl[190] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_191 br[190] vdd vss bl[190] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_191 br[190] vdd vss bl[190] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_191 br[190] vdd vss bl[190] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_191 br[190] vdd vss bl[190] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_191 br[190] vdd vss bl[190] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_191 br[190] vdd vss bl[190] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_191 br[190] vdd vss bl[190] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_191 br[190] vdd vss bl[190] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_191 br[190] vdd vss bl[190] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_191 br[190] vdd vss bl[190] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_191 br[190] vdd vss bl[190] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_191 br[190] vdd vss bl[190] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_191 br[190] vdd vss bl[190] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_191 br[190] vdd vss bl[190] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_191 br[190] vdd vss bl[190] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_192 br[191] vdd vss bl[191] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_192 br[191] vdd vss bl[191] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_192 br[191] vdd vss bl[191] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_192 br[191] vdd vss bl[191] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_192 br[191] vdd vss bl[191] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_192 br[191] vdd vss bl[191] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_192 br[191] vdd vss bl[191] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_192 br[191] vdd vss bl[191] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_192 br[191] vdd vss bl[191] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_192 br[191] vdd vss bl[191] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_192 br[191] vdd vss bl[191] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_192 br[191] vdd vss bl[191] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_192 br[191] vdd vss bl[191] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_192 br[191] vdd vss bl[191] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_192 br[191] vdd vss bl[191] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_192 br[191] vdd vss bl[191] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_192 br[191] vdd vss bl[191] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_192 br[191] vdd vss bl[191] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_192 br[191] vdd vss bl[191] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_193 br[192] vdd vss bl[192] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_193 br[192] vdd vss bl[192] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_193 br[192] vdd vss bl[192] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_193 br[192] vdd vss bl[192] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_193 br[192] vdd vss bl[192] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_193 br[192] vdd vss bl[192] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_193 br[192] vdd vss bl[192] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_193 br[192] vdd vss bl[192] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_193 br[192] vdd vss bl[192] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_193 br[192] vdd vss bl[192] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_193 br[192] vdd vss bl[192] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_193 br[192] vdd vss bl[192] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_193 br[192] vdd vss bl[192] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_193 br[192] vdd vss bl[192] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_193 br[192] vdd vss bl[192] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_193 br[192] vdd vss bl[192] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_193 br[192] vdd vss bl[192] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_193 br[192] vdd vss bl[192] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_193 br[192] vdd vss bl[192] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_194 br[193] vdd vss bl[193] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_194 br[193] vdd vss bl[193] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_194 br[193] vdd vss bl[193] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_194 br[193] vdd vss bl[193] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_194 br[193] vdd vss bl[193] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_194 br[193] vdd vss bl[193] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_194 br[193] vdd vss bl[193] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_194 br[193] vdd vss bl[193] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_194 br[193] vdd vss bl[193] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_194 br[193] vdd vss bl[193] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_194 br[193] vdd vss bl[193] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_194 br[193] vdd vss bl[193] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_194 br[193] vdd vss bl[193] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_194 br[193] vdd vss bl[193] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_194 br[193] vdd vss bl[193] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_194 br[193] vdd vss bl[193] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_194 br[193] vdd vss bl[193] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_194 br[193] vdd vss bl[193] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_194 br[193] vdd vss bl[193] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_195 br[194] vdd vss bl[194] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_195 br[194] vdd vss bl[194] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_195 br[194] vdd vss bl[194] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_195 br[194] vdd vss bl[194] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_195 br[194] vdd vss bl[194] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_195 br[194] vdd vss bl[194] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_195 br[194] vdd vss bl[194] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_195 br[194] vdd vss bl[194] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_195 br[194] vdd vss bl[194] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_195 br[194] vdd vss bl[194] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_195 br[194] vdd vss bl[194] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_195 br[194] vdd vss bl[194] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_195 br[194] vdd vss bl[194] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_195 br[194] vdd vss bl[194] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_195 br[194] vdd vss bl[194] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_195 br[194] vdd vss bl[194] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_195 br[194] vdd vss bl[194] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_195 br[194] vdd vss bl[194] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_195 br[194] vdd vss bl[194] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_196 br[195] vdd vss bl[195] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_196 br[195] vdd vss bl[195] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_196 br[195] vdd vss bl[195] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_196 br[195] vdd vss bl[195] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_196 br[195] vdd vss bl[195] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_196 br[195] vdd vss bl[195] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_196 br[195] vdd vss bl[195] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_196 br[195] vdd vss bl[195] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_196 br[195] vdd vss bl[195] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_196 br[195] vdd vss bl[195] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_196 br[195] vdd vss bl[195] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_196 br[195] vdd vss bl[195] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_196 br[195] vdd vss bl[195] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_196 br[195] vdd vss bl[195] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_196 br[195] vdd vss bl[195] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_196 br[195] vdd vss bl[195] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_196 br[195] vdd vss bl[195] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_196 br[195] vdd vss bl[195] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_196 br[195] vdd vss bl[195] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_197 br[196] vdd vss bl[196] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_197 br[196] vdd vss bl[196] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_197 br[196] vdd vss bl[196] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_197 br[196] vdd vss bl[196] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_197 br[196] vdd vss bl[196] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_197 br[196] vdd vss bl[196] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_197 br[196] vdd vss bl[196] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_197 br[196] vdd vss bl[196] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_197 br[196] vdd vss bl[196] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_197 br[196] vdd vss bl[196] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_197 br[196] vdd vss bl[196] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_197 br[196] vdd vss bl[196] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_197 br[196] vdd vss bl[196] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_197 br[196] vdd vss bl[196] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_197 br[196] vdd vss bl[196] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_197 br[196] vdd vss bl[196] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_197 br[196] vdd vss bl[196] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_197 br[196] vdd vss bl[196] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_197 br[196] vdd vss bl[196] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_198 br[197] vdd vss bl[197] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_198 br[197] vdd vss bl[197] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_198 br[197] vdd vss bl[197] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_198 br[197] vdd vss bl[197] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_198 br[197] vdd vss bl[197] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_198 br[197] vdd vss bl[197] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_198 br[197] vdd vss bl[197] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_198 br[197] vdd vss bl[197] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_198 br[197] vdd vss bl[197] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_198 br[197] vdd vss bl[197] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_198 br[197] vdd vss bl[197] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_198 br[197] vdd vss bl[197] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_198 br[197] vdd vss bl[197] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_198 br[197] vdd vss bl[197] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_198 br[197] vdd vss bl[197] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_198 br[197] vdd vss bl[197] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_198 br[197] vdd vss bl[197] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_198 br[197] vdd vss bl[197] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_198 br[197] vdd vss bl[197] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_199 br[198] vdd vss bl[198] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_199 br[198] vdd vss bl[198] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_199 br[198] vdd vss bl[198] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_199 br[198] vdd vss bl[198] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_199 br[198] vdd vss bl[198] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_199 br[198] vdd vss bl[198] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_199 br[198] vdd vss bl[198] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_199 br[198] vdd vss bl[198] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_199 br[198] vdd vss bl[198] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_199 br[198] vdd vss bl[198] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_199 br[198] vdd vss bl[198] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_199 br[198] vdd vss bl[198] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_199 br[198] vdd vss bl[198] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_199 br[198] vdd vss bl[198] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_199 br[198] vdd vss bl[198] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_199 br[198] vdd vss bl[198] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_199 br[198] vdd vss bl[198] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_199 br[198] vdd vss bl[198] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_199 br[198] vdd vss bl[198] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_200 br[199] vdd vss bl[199] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_200 br[199] vdd vss bl[199] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_200 br[199] vdd vss bl[199] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_200 br[199] vdd vss bl[199] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_200 br[199] vdd vss bl[199] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_200 br[199] vdd vss bl[199] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_200 br[199] vdd vss bl[199] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_200 br[199] vdd vss bl[199] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_200 br[199] vdd vss bl[199] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_200 br[199] vdd vss bl[199] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_200 br[199] vdd vss bl[199] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_200 br[199] vdd vss bl[199] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_200 br[199] vdd vss bl[199] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_200 br[199] vdd vss bl[199] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_200 br[199] vdd vss bl[199] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_200 br[199] vdd vss bl[199] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_200 br[199] vdd vss bl[199] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_200 br[199] vdd vss bl[199] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_200 br[199] vdd vss bl[199] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_201 br[200] vdd vss bl[200] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_201 br[200] vdd vss bl[200] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_201 br[200] vdd vss bl[200] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_201 br[200] vdd vss bl[200] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_201 br[200] vdd vss bl[200] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_201 br[200] vdd vss bl[200] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_201 br[200] vdd vss bl[200] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_201 br[200] vdd vss bl[200] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_201 br[200] vdd vss bl[200] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_201 br[200] vdd vss bl[200] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_201 br[200] vdd vss bl[200] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_201 br[200] vdd vss bl[200] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_201 br[200] vdd vss bl[200] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_201 br[200] vdd vss bl[200] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_201 br[200] vdd vss bl[200] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_201 br[200] vdd vss bl[200] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_201 br[200] vdd vss bl[200] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_201 br[200] vdd vss bl[200] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_201 br[200] vdd vss bl[200] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_202 br[201] vdd vss bl[201] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_202 br[201] vdd vss bl[201] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_202 br[201] vdd vss bl[201] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_202 br[201] vdd vss bl[201] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_202 br[201] vdd vss bl[201] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_202 br[201] vdd vss bl[201] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_202 br[201] vdd vss bl[201] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_202 br[201] vdd vss bl[201] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_202 br[201] vdd vss bl[201] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_202 br[201] vdd vss bl[201] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_202 br[201] vdd vss bl[201] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_202 br[201] vdd vss bl[201] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_202 br[201] vdd vss bl[201] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_202 br[201] vdd vss bl[201] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_202 br[201] vdd vss bl[201] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_202 br[201] vdd vss bl[201] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_202 br[201] vdd vss bl[201] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_202 br[201] vdd vss bl[201] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_202 br[201] vdd vss bl[201] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_203 br[202] vdd vss bl[202] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_203 br[202] vdd vss bl[202] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_203 br[202] vdd vss bl[202] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_203 br[202] vdd vss bl[202] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_203 br[202] vdd vss bl[202] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_203 br[202] vdd vss bl[202] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_203 br[202] vdd vss bl[202] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_203 br[202] vdd vss bl[202] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_203 br[202] vdd vss bl[202] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_203 br[202] vdd vss bl[202] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_203 br[202] vdd vss bl[202] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_203 br[202] vdd vss bl[202] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_203 br[202] vdd vss bl[202] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_203 br[202] vdd vss bl[202] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_203 br[202] vdd vss bl[202] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_203 br[202] vdd vss bl[202] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_203 br[202] vdd vss bl[202] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_203 br[202] vdd vss bl[202] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_203 br[202] vdd vss bl[202] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_204 br[203] vdd vss bl[203] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_204 br[203] vdd vss bl[203] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_204 br[203] vdd vss bl[203] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_204 br[203] vdd vss bl[203] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_204 br[203] vdd vss bl[203] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_204 br[203] vdd vss bl[203] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_204 br[203] vdd vss bl[203] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_204 br[203] vdd vss bl[203] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_204 br[203] vdd vss bl[203] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_204 br[203] vdd vss bl[203] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_204 br[203] vdd vss bl[203] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_204 br[203] vdd vss bl[203] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_204 br[203] vdd vss bl[203] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_204 br[203] vdd vss bl[203] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_204 br[203] vdd vss bl[203] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_204 br[203] vdd vss bl[203] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_204 br[203] vdd vss bl[203] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_204 br[203] vdd vss bl[203] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_204 br[203] vdd vss bl[203] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_205 br[204] vdd vss bl[204] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_205 br[204] vdd vss bl[204] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_205 br[204] vdd vss bl[204] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_205 br[204] vdd vss bl[204] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_205 br[204] vdd vss bl[204] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_205 br[204] vdd vss bl[204] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_205 br[204] vdd vss bl[204] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_205 br[204] vdd vss bl[204] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_205 br[204] vdd vss bl[204] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_205 br[204] vdd vss bl[204] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_205 br[204] vdd vss bl[204] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_205 br[204] vdd vss bl[204] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_205 br[204] vdd vss bl[204] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_205 br[204] vdd vss bl[204] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_205 br[204] vdd vss bl[204] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_205 br[204] vdd vss bl[204] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_205 br[204] vdd vss bl[204] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_205 br[204] vdd vss bl[204] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_205 br[204] vdd vss bl[204] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_206 br[205] vdd vss bl[205] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_206 br[205] vdd vss bl[205] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_206 br[205] vdd vss bl[205] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_206 br[205] vdd vss bl[205] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_206 br[205] vdd vss bl[205] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_206 br[205] vdd vss bl[205] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_206 br[205] vdd vss bl[205] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_206 br[205] vdd vss bl[205] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_206 br[205] vdd vss bl[205] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_206 br[205] vdd vss bl[205] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_206 br[205] vdd vss bl[205] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_206 br[205] vdd vss bl[205] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_206 br[205] vdd vss bl[205] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_206 br[205] vdd vss bl[205] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_206 br[205] vdd vss bl[205] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_206 br[205] vdd vss bl[205] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_206 br[205] vdd vss bl[205] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_206 br[205] vdd vss bl[205] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_206 br[205] vdd vss bl[205] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_207 br[206] vdd vss bl[206] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_207 br[206] vdd vss bl[206] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_207 br[206] vdd vss bl[206] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_207 br[206] vdd vss bl[206] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_207 br[206] vdd vss bl[206] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_207 br[206] vdd vss bl[206] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_207 br[206] vdd vss bl[206] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_207 br[206] vdd vss bl[206] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_207 br[206] vdd vss bl[206] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_207 br[206] vdd vss bl[206] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_207 br[206] vdd vss bl[206] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_207 br[206] vdd vss bl[206] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_207 br[206] vdd vss bl[206] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_207 br[206] vdd vss bl[206] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_207 br[206] vdd vss bl[206] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_207 br[206] vdd vss bl[206] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_207 br[206] vdd vss bl[206] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_207 br[206] vdd vss bl[206] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_207 br[206] vdd vss bl[206] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_208 br[207] vdd vss bl[207] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_208 br[207] vdd vss bl[207] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_208 br[207] vdd vss bl[207] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_208 br[207] vdd vss bl[207] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_208 br[207] vdd vss bl[207] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_208 br[207] vdd vss bl[207] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_208 br[207] vdd vss bl[207] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_208 br[207] vdd vss bl[207] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_208 br[207] vdd vss bl[207] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_208 br[207] vdd vss bl[207] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_208 br[207] vdd vss bl[207] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_208 br[207] vdd vss bl[207] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_208 br[207] vdd vss bl[207] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_208 br[207] vdd vss bl[207] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_208 br[207] vdd vss bl[207] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_208 br[207] vdd vss bl[207] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_208 br[207] vdd vss bl[207] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_208 br[207] vdd vss bl[207] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_208 br[207] vdd vss bl[207] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_209 br[208] vdd vss bl[208] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_209 br[208] vdd vss bl[208] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_209 br[208] vdd vss bl[208] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_209 br[208] vdd vss bl[208] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_209 br[208] vdd vss bl[208] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_209 br[208] vdd vss bl[208] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_209 br[208] vdd vss bl[208] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_209 br[208] vdd vss bl[208] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_209 br[208] vdd vss bl[208] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_209 br[208] vdd vss bl[208] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_209 br[208] vdd vss bl[208] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_209 br[208] vdd vss bl[208] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_209 br[208] vdd vss bl[208] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_209 br[208] vdd vss bl[208] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_209 br[208] vdd vss bl[208] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_209 br[208] vdd vss bl[208] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_209 br[208] vdd vss bl[208] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_209 br[208] vdd vss bl[208] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_209 br[208] vdd vss bl[208] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_210 br[209] vdd vss bl[209] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_210 br[209] vdd vss bl[209] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_210 br[209] vdd vss bl[209] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_210 br[209] vdd vss bl[209] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_210 br[209] vdd vss bl[209] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_210 br[209] vdd vss bl[209] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_210 br[209] vdd vss bl[209] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_210 br[209] vdd vss bl[209] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_210 br[209] vdd vss bl[209] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_210 br[209] vdd vss bl[209] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_210 br[209] vdd vss bl[209] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_210 br[209] vdd vss bl[209] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_210 br[209] vdd vss bl[209] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_210 br[209] vdd vss bl[209] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_210 br[209] vdd vss bl[209] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_210 br[209] vdd vss bl[209] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_210 br[209] vdd vss bl[209] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_210 br[209] vdd vss bl[209] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_210 br[209] vdd vss bl[209] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_211 br[210] vdd vss bl[210] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_211 br[210] vdd vss bl[210] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_211 br[210] vdd vss bl[210] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_211 br[210] vdd vss bl[210] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_211 br[210] vdd vss bl[210] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_211 br[210] vdd vss bl[210] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_211 br[210] vdd vss bl[210] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_211 br[210] vdd vss bl[210] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_211 br[210] vdd vss bl[210] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_211 br[210] vdd vss bl[210] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_211 br[210] vdd vss bl[210] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_211 br[210] vdd vss bl[210] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_211 br[210] vdd vss bl[210] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_211 br[210] vdd vss bl[210] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_211 br[210] vdd vss bl[210] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_211 br[210] vdd vss bl[210] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_211 br[210] vdd vss bl[210] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_211 br[210] vdd vss bl[210] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_211 br[210] vdd vss bl[210] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_212 br[211] vdd vss bl[211] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_212 br[211] vdd vss bl[211] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_212 br[211] vdd vss bl[211] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_212 br[211] vdd vss bl[211] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_212 br[211] vdd vss bl[211] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_212 br[211] vdd vss bl[211] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_212 br[211] vdd vss bl[211] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_212 br[211] vdd vss bl[211] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_212 br[211] vdd vss bl[211] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_212 br[211] vdd vss bl[211] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_212 br[211] vdd vss bl[211] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_212 br[211] vdd vss bl[211] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_212 br[211] vdd vss bl[211] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_212 br[211] vdd vss bl[211] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_212 br[211] vdd vss bl[211] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_212 br[211] vdd vss bl[211] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_212 br[211] vdd vss bl[211] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_212 br[211] vdd vss bl[211] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_212 br[211] vdd vss bl[211] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_213 br[212] vdd vss bl[212] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_213 br[212] vdd vss bl[212] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_213 br[212] vdd vss bl[212] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_213 br[212] vdd vss bl[212] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_213 br[212] vdd vss bl[212] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_213 br[212] vdd vss bl[212] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_213 br[212] vdd vss bl[212] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_213 br[212] vdd vss bl[212] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_213 br[212] vdd vss bl[212] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_213 br[212] vdd vss bl[212] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_213 br[212] vdd vss bl[212] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_213 br[212] vdd vss bl[212] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_213 br[212] vdd vss bl[212] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_213 br[212] vdd vss bl[212] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_213 br[212] vdd vss bl[212] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_213 br[212] vdd vss bl[212] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_213 br[212] vdd vss bl[212] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_213 br[212] vdd vss bl[212] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_213 br[212] vdd vss bl[212] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_214 br[213] vdd vss bl[213] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_214 br[213] vdd vss bl[213] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_214 br[213] vdd vss bl[213] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_214 br[213] vdd vss bl[213] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_214 br[213] vdd vss bl[213] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_214 br[213] vdd vss bl[213] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_214 br[213] vdd vss bl[213] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_214 br[213] vdd vss bl[213] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_214 br[213] vdd vss bl[213] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_214 br[213] vdd vss bl[213] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_214 br[213] vdd vss bl[213] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_214 br[213] vdd vss bl[213] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_214 br[213] vdd vss bl[213] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_214 br[213] vdd vss bl[213] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_214 br[213] vdd vss bl[213] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_214 br[213] vdd vss bl[213] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_214 br[213] vdd vss bl[213] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_214 br[213] vdd vss bl[213] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_214 br[213] vdd vss bl[213] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_215 br[214] vdd vss bl[214] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_215 br[214] vdd vss bl[214] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_215 br[214] vdd vss bl[214] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_215 br[214] vdd vss bl[214] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_215 br[214] vdd vss bl[214] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_215 br[214] vdd vss bl[214] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_215 br[214] vdd vss bl[214] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_215 br[214] vdd vss bl[214] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_215 br[214] vdd vss bl[214] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_215 br[214] vdd vss bl[214] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_215 br[214] vdd vss bl[214] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_215 br[214] vdd vss bl[214] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_215 br[214] vdd vss bl[214] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_215 br[214] vdd vss bl[214] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_215 br[214] vdd vss bl[214] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_215 br[214] vdd vss bl[214] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_215 br[214] vdd vss bl[214] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_215 br[214] vdd vss bl[214] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_215 br[214] vdd vss bl[214] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_216 br[215] vdd vss bl[215] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_216 br[215] vdd vss bl[215] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_216 br[215] vdd vss bl[215] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_216 br[215] vdd vss bl[215] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_216 br[215] vdd vss bl[215] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_216 br[215] vdd vss bl[215] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_216 br[215] vdd vss bl[215] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_216 br[215] vdd vss bl[215] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_216 br[215] vdd vss bl[215] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_216 br[215] vdd vss bl[215] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_216 br[215] vdd vss bl[215] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_216 br[215] vdd vss bl[215] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_216 br[215] vdd vss bl[215] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_216 br[215] vdd vss bl[215] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_216 br[215] vdd vss bl[215] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_216 br[215] vdd vss bl[215] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_216 br[215] vdd vss bl[215] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_216 br[215] vdd vss bl[215] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_216 br[215] vdd vss bl[215] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_217 br[216] vdd vss bl[216] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_217 br[216] vdd vss bl[216] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_217 br[216] vdd vss bl[216] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_217 br[216] vdd vss bl[216] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_217 br[216] vdd vss bl[216] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_217 br[216] vdd vss bl[216] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_217 br[216] vdd vss bl[216] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_217 br[216] vdd vss bl[216] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_217 br[216] vdd vss bl[216] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_217 br[216] vdd vss bl[216] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_217 br[216] vdd vss bl[216] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_217 br[216] vdd vss bl[216] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_217 br[216] vdd vss bl[216] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_217 br[216] vdd vss bl[216] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_217 br[216] vdd vss bl[216] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_217 br[216] vdd vss bl[216] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_217 br[216] vdd vss bl[216] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_217 br[216] vdd vss bl[216] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_217 br[216] vdd vss bl[216] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_218 br[217] vdd vss bl[217] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_218 br[217] vdd vss bl[217] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_218 br[217] vdd vss bl[217] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_218 br[217] vdd vss bl[217] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_218 br[217] vdd vss bl[217] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_218 br[217] vdd vss bl[217] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_218 br[217] vdd vss bl[217] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_218 br[217] vdd vss bl[217] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_218 br[217] vdd vss bl[217] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_218 br[217] vdd vss bl[217] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_218 br[217] vdd vss bl[217] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_218 br[217] vdd vss bl[217] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_218 br[217] vdd vss bl[217] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_218 br[217] vdd vss bl[217] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_218 br[217] vdd vss bl[217] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_218 br[217] vdd vss bl[217] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_218 br[217] vdd vss bl[217] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_218 br[217] vdd vss bl[217] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_218 br[217] vdd vss bl[217] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_219 br[218] vdd vss bl[218] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_219 br[218] vdd vss bl[218] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_219 br[218] vdd vss bl[218] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_219 br[218] vdd vss bl[218] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_219 br[218] vdd vss bl[218] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_219 br[218] vdd vss bl[218] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_219 br[218] vdd vss bl[218] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_219 br[218] vdd vss bl[218] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_219 br[218] vdd vss bl[218] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_219 br[218] vdd vss bl[218] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_219 br[218] vdd vss bl[218] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_219 br[218] vdd vss bl[218] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_219 br[218] vdd vss bl[218] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_219 br[218] vdd vss bl[218] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_219 br[218] vdd vss bl[218] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_219 br[218] vdd vss bl[218] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_219 br[218] vdd vss bl[218] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_219 br[218] vdd vss bl[218] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_219 br[218] vdd vss bl[218] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_220 br[219] vdd vss bl[219] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_220 br[219] vdd vss bl[219] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_220 br[219] vdd vss bl[219] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_220 br[219] vdd vss bl[219] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_220 br[219] vdd vss bl[219] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_220 br[219] vdd vss bl[219] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_220 br[219] vdd vss bl[219] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_220 br[219] vdd vss bl[219] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_220 br[219] vdd vss bl[219] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_220 br[219] vdd vss bl[219] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_220 br[219] vdd vss bl[219] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_220 br[219] vdd vss bl[219] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_220 br[219] vdd vss bl[219] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_220 br[219] vdd vss bl[219] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_220 br[219] vdd vss bl[219] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_220 br[219] vdd vss bl[219] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_220 br[219] vdd vss bl[219] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_220 br[219] vdd vss bl[219] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_220 br[219] vdd vss bl[219] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_221 br[220] vdd vss bl[220] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_221 br[220] vdd vss bl[220] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_221 br[220] vdd vss bl[220] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_221 br[220] vdd vss bl[220] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_221 br[220] vdd vss bl[220] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_221 br[220] vdd vss bl[220] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_221 br[220] vdd vss bl[220] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_221 br[220] vdd vss bl[220] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_221 br[220] vdd vss bl[220] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_221 br[220] vdd vss bl[220] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_221 br[220] vdd vss bl[220] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_221 br[220] vdd vss bl[220] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_221 br[220] vdd vss bl[220] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_221 br[220] vdd vss bl[220] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_221 br[220] vdd vss bl[220] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_221 br[220] vdd vss bl[220] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_221 br[220] vdd vss bl[220] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_221 br[220] vdd vss bl[220] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_221 br[220] vdd vss bl[220] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_222 br[221] vdd vss bl[221] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_222 br[221] vdd vss bl[221] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_222 br[221] vdd vss bl[221] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_222 br[221] vdd vss bl[221] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_222 br[221] vdd vss bl[221] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_222 br[221] vdd vss bl[221] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_222 br[221] vdd vss bl[221] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_222 br[221] vdd vss bl[221] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_222 br[221] vdd vss bl[221] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_222 br[221] vdd vss bl[221] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_222 br[221] vdd vss bl[221] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_222 br[221] vdd vss bl[221] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_222 br[221] vdd vss bl[221] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_222 br[221] vdd vss bl[221] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_222 br[221] vdd vss bl[221] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_222 br[221] vdd vss bl[221] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_222 br[221] vdd vss bl[221] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_222 br[221] vdd vss bl[221] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_222 br[221] vdd vss bl[221] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_223 br[222] vdd vss bl[222] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_223 br[222] vdd vss bl[222] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_223 br[222] vdd vss bl[222] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_223 br[222] vdd vss bl[222] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_223 br[222] vdd vss bl[222] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_223 br[222] vdd vss bl[222] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_223 br[222] vdd vss bl[222] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_223 br[222] vdd vss bl[222] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_223 br[222] vdd vss bl[222] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_223 br[222] vdd vss bl[222] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_223 br[222] vdd vss bl[222] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_223 br[222] vdd vss bl[222] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_223 br[222] vdd vss bl[222] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_223 br[222] vdd vss bl[222] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_223 br[222] vdd vss bl[222] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_223 br[222] vdd vss bl[222] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_223 br[222] vdd vss bl[222] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_223 br[222] vdd vss bl[222] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_223 br[222] vdd vss bl[222] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_224 br[223] vdd vss bl[223] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_224 br[223] vdd vss bl[223] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_224 br[223] vdd vss bl[223] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_224 br[223] vdd vss bl[223] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_224 br[223] vdd vss bl[223] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_224 br[223] vdd vss bl[223] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_224 br[223] vdd vss bl[223] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_224 br[223] vdd vss bl[223] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_224 br[223] vdd vss bl[223] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_224 br[223] vdd vss bl[223] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_224 br[223] vdd vss bl[223] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_224 br[223] vdd vss bl[223] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_224 br[223] vdd vss bl[223] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_224 br[223] vdd vss bl[223] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_224 br[223] vdd vss bl[223] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_224 br[223] vdd vss bl[223] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_224 br[223] vdd vss bl[223] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_224 br[223] vdd vss bl[223] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_224 br[223] vdd vss bl[223] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_225 br[224] vdd vss bl[224] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_225 br[224] vdd vss bl[224] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_225 br[224] vdd vss bl[224] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_225 br[224] vdd vss bl[224] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_225 br[224] vdd vss bl[224] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_225 br[224] vdd vss bl[224] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_225 br[224] vdd vss bl[224] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_225 br[224] vdd vss bl[224] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_225 br[224] vdd vss bl[224] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_225 br[224] vdd vss bl[224] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_225 br[224] vdd vss bl[224] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_225 br[224] vdd vss bl[224] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_225 br[224] vdd vss bl[224] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_225 br[224] vdd vss bl[224] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_225 br[224] vdd vss bl[224] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_225 br[224] vdd vss bl[224] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_225 br[224] vdd vss bl[224] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_225 br[224] vdd vss bl[224] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_225 br[224] vdd vss bl[224] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_226 br[225] vdd vss bl[225] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_226 br[225] vdd vss bl[225] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_226 br[225] vdd vss bl[225] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_226 br[225] vdd vss bl[225] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_226 br[225] vdd vss bl[225] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_226 br[225] vdd vss bl[225] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_226 br[225] vdd vss bl[225] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_226 br[225] vdd vss bl[225] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_226 br[225] vdd vss bl[225] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_226 br[225] vdd vss bl[225] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_226 br[225] vdd vss bl[225] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_226 br[225] vdd vss bl[225] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_226 br[225] vdd vss bl[225] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_226 br[225] vdd vss bl[225] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_226 br[225] vdd vss bl[225] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_226 br[225] vdd vss bl[225] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_226 br[225] vdd vss bl[225] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_226 br[225] vdd vss bl[225] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_226 br[225] vdd vss bl[225] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_227 br[226] vdd vss bl[226] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_227 br[226] vdd vss bl[226] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_227 br[226] vdd vss bl[226] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_227 br[226] vdd vss bl[226] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_227 br[226] vdd vss bl[226] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_227 br[226] vdd vss bl[226] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_227 br[226] vdd vss bl[226] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_227 br[226] vdd vss bl[226] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_227 br[226] vdd vss bl[226] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_227 br[226] vdd vss bl[226] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_227 br[226] vdd vss bl[226] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_227 br[226] vdd vss bl[226] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_227 br[226] vdd vss bl[226] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_227 br[226] vdd vss bl[226] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_227 br[226] vdd vss bl[226] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_227 br[226] vdd vss bl[226] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_227 br[226] vdd vss bl[226] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_227 br[226] vdd vss bl[226] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_227 br[226] vdd vss bl[226] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_228 br[227] vdd vss bl[227] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_228 br[227] vdd vss bl[227] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_228 br[227] vdd vss bl[227] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_228 br[227] vdd vss bl[227] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_228 br[227] vdd vss bl[227] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_228 br[227] vdd vss bl[227] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_228 br[227] vdd vss bl[227] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_228 br[227] vdd vss bl[227] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_228 br[227] vdd vss bl[227] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_228 br[227] vdd vss bl[227] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_228 br[227] vdd vss bl[227] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_228 br[227] vdd vss bl[227] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_228 br[227] vdd vss bl[227] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_228 br[227] vdd vss bl[227] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_228 br[227] vdd vss bl[227] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_228 br[227] vdd vss bl[227] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_228 br[227] vdd vss bl[227] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_228 br[227] vdd vss bl[227] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_228 br[227] vdd vss bl[227] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_229 br[228] vdd vss bl[228] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_229 br[228] vdd vss bl[228] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_229 br[228] vdd vss bl[228] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_229 br[228] vdd vss bl[228] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_229 br[228] vdd vss bl[228] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_229 br[228] vdd vss bl[228] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_229 br[228] vdd vss bl[228] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_229 br[228] vdd vss bl[228] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_229 br[228] vdd vss bl[228] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_229 br[228] vdd vss bl[228] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_229 br[228] vdd vss bl[228] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_229 br[228] vdd vss bl[228] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_229 br[228] vdd vss bl[228] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_229 br[228] vdd vss bl[228] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_229 br[228] vdd vss bl[228] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_229 br[228] vdd vss bl[228] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_229 br[228] vdd vss bl[228] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_229 br[228] vdd vss bl[228] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_229 br[228] vdd vss bl[228] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_230 br[229] vdd vss bl[229] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_230 br[229] vdd vss bl[229] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_230 br[229] vdd vss bl[229] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_230 br[229] vdd vss bl[229] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_230 br[229] vdd vss bl[229] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_230 br[229] vdd vss bl[229] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_230 br[229] vdd vss bl[229] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_230 br[229] vdd vss bl[229] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_230 br[229] vdd vss bl[229] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_230 br[229] vdd vss bl[229] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_230 br[229] vdd vss bl[229] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_230 br[229] vdd vss bl[229] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_230 br[229] vdd vss bl[229] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_230 br[229] vdd vss bl[229] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_230 br[229] vdd vss bl[229] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_230 br[229] vdd vss bl[229] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_230 br[229] vdd vss bl[229] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_230 br[229] vdd vss bl[229] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_230 br[229] vdd vss bl[229] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_231 br[230] vdd vss bl[230] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_231 br[230] vdd vss bl[230] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_231 br[230] vdd vss bl[230] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_231 br[230] vdd vss bl[230] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_231 br[230] vdd vss bl[230] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_231 br[230] vdd vss bl[230] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_231 br[230] vdd vss bl[230] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_231 br[230] vdd vss bl[230] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_231 br[230] vdd vss bl[230] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_231 br[230] vdd vss bl[230] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_231 br[230] vdd vss bl[230] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_231 br[230] vdd vss bl[230] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_231 br[230] vdd vss bl[230] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_231 br[230] vdd vss bl[230] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_231 br[230] vdd vss bl[230] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_231 br[230] vdd vss bl[230] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_231 br[230] vdd vss bl[230] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_231 br[230] vdd vss bl[230] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_231 br[230] vdd vss bl[230] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_232 br[231] vdd vss bl[231] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_232 br[231] vdd vss bl[231] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_232 br[231] vdd vss bl[231] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_232 br[231] vdd vss bl[231] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_232 br[231] vdd vss bl[231] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_232 br[231] vdd vss bl[231] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_232 br[231] vdd vss bl[231] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_232 br[231] vdd vss bl[231] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_232 br[231] vdd vss bl[231] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_232 br[231] vdd vss bl[231] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_232 br[231] vdd vss bl[231] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_232 br[231] vdd vss bl[231] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_232 br[231] vdd vss bl[231] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_232 br[231] vdd vss bl[231] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_232 br[231] vdd vss bl[231] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_232 br[231] vdd vss bl[231] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_232 br[231] vdd vss bl[231] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_232 br[231] vdd vss bl[231] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_232 br[231] vdd vss bl[231] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_233 br[232] vdd vss bl[232] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_233 br[232] vdd vss bl[232] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_233 br[232] vdd vss bl[232] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_233 br[232] vdd vss bl[232] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_233 br[232] vdd vss bl[232] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_233 br[232] vdd vss bl[232] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_233 br[232] vdd vss bl[232] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_233 br[232] vdd vss bl[232] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_233 br[232] vdd vss bl[232] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_233 br[232] vdd vss bl[232] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_233 br[232] vdd vss bl[232] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_233 br[232] vdd vss bl[232] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_233 br[232] vdd vss bl[232] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_233 br[232] vdd vss bl[232] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_233 br[232] vdd vss bl[232] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_233 br[232] vdd vss bl[232] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_233 br[232] vdd vss bl[232] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_233 br[232] vdd vss bl[232] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_233 br[232] vdd vss bl[232] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_234 br[233] vdd vss bl[233] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_234 br[233] vdd vss bl[233] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_234 br[233] vdd vss bl[233] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_234 br[233] vdd vss bl[233] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_234 br[233] vdd vss bl[233] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_234 br[233] vdd vss bl[233] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_234 br[233] vdd vss bl[233] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_234 br[233] vdd vss bl[233] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_234 br[233] vdd vss bl[233] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_234 br[233] vdd vss bl[233] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_234 br[233] vdd vss bl[233] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_234 br[233] vdd vss bl[233] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_234 br[233] vdd vss bl[233] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_234 br[233] vdd vss bl[233] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_234 br[233] vdd vss bl[233] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_234 br[233] vdd vss bl[233] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_234 br[233] vdd vss bl[233] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_234 br[233] vdd vss bl[233] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_234 br[233] vdd vss bl[233] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_235 br[234] vdd vss bl[234] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_235 br[234] vdd vss bl[234] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_235 br[234] vdd vss bl[234] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_235 br[234] vdd vss bl[234] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_235 br[234] vdd vss bl[234] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_235 br[234] vdd vss bl[234] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_235 br[234] vdd vss bl[234] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_235 br[234] vdd vss bl[234] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_235 br[234] vdd vss bl[234] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_235 br[234] vdd vss bl[234] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_235 br[234] vdd vss bl[234] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_235 br[234] vdd vss bl[234] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_235 br[234] vdd vss bl[234] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_235 br[234] vdd vss bl[234] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_235 br[234] vdd vss bl[234] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_235 br[234] vdd vss bl[234] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_235 br[234] vdd vss bl[234] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_235 br[234] vdd vss bl[234] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_235 br[234] vdd vss bl[234] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_236 br[235] vdd vss bl[235] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_236 br[235] vdd vss bl[235] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_236 br[235] vdd vss bl[235] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_236 br[235] vdd vss bl[235] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_236 br[235] vdd vss bl[235] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_236 br[235] vdd vss bl[235] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_236 br[235] vdd vss bl[235] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_236 br[235] vdd vss bl[235] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_236 br[235] vdd vss bl[235] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_236 br[235] vdd vss bl[235] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_236 br[235] vdd vss bl[235] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_236 br[235] vdd vss bl[235] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_236 br[235] vdd vss bl[235] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_236 br[235] vdd vss bl[235] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_236 br[235] vdd vss bl[235] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_236 br[235] vdd vss bl[235] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_236 br[235] vdd vss bl[235] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_236 br[235] vdd vss bl[235] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_236 br[235] vdd vss bl[235] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_237 br[236] vdd vss bl[236] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_237 br[236] vdd vss bl[236] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_237 br[236] vdd vss bl[236] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_237 br[236] vdd vss bl[236] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_237 br[236] vdd vss bl[236] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_237 br[236] vdd vss bl[236] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_237 br[236] vdd vss bl[236] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_237 br[236] vdd vss bl[236] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_237 br[236] vdd vss bl[236] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_237 br[236] vdd vss bl[236] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_237 br[236] vdd vss bl[236] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_237 br[236] vdd vss bl[236] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_237 br[236] vdd vss bl[236] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_237 br[236] vdd vss bl[236] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_237 br[236] vdd vss bl[236] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_237 br[236] vdd vss bl[236] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_237 br[236] vdd vss bl[236] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_237 br[236] vdd vss bl[236] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_237 br[236] vdd vss bl[236] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_238 br[237] vdd vss bl[237] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_238 br[237] vdd vss bl[237] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_238 br[237] vdd vss bl[237] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_238 br[237] vdd vss bl[237] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_238 br[237] vdd vss bl[237] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_238 br[237] vdd vss bl[237] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_238 br[237] vdd vss bl[237] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_238 br[237] vdd vss bl[237] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_238 br[237] vdd vss bl[237] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_238 br[237] vdd vss bl[237] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_238 br[237] vdd vss bl[237] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_238 br[237] vdd vss bl[237] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_238 br[237] vdd vss bl[237] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_238 br[237] vdd vss bl[237] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_238 br[237] vdd vss bl[237] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_238 br[237] vdd vss bl[237] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_238 br[237] vdd vss bl[237] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_238 br[237] vdd vss bl[237] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_238 br[237] vdd vss bl[237] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_239 br[238] vdd vss bl[238] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_239 br[238] vdd vss bl[238] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_239 br[238] vdd vss bl[238] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_239 br[238] vdd vss bl[238] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_239 br[238] vdd vss bl[238] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_239 br[238] vdd vss bl[238] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_239 br[238] vdd vss bl[238] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_239 br[238] vdd vss bl[238] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_239 br[238] vdd vss bl[238] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_239 br[238] vdd vss bl[238] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_239 br[238] vdd vss bl[238] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_239 br[238] vdd vss bl[238] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_239 br[238] vdd vss bl[238] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_239 br[238] vdd vss bl[238] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_239 br[238] vdd vss bl[238] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_239 br[238] vdd vss bl[238] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_239 br[238] vdd vss bl[238] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_239 br[238] vdd vss bl[238] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_239 br[238] vdd vss bl[238] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_240 br[239] vdd vss bl[239] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_240 br[239] vdd vss bl[239] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_240 br[239] vdd vss bl[239] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_240 br[239] vdd vss bl[239] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_240 br[239] vdd vss bl[239] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_240 br[239] vdd vss bl[239] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_240 br[239] vdd vss bl[239] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_240 br[239] vdd vss bl[239] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_240 br[239] vdd vss bl[239] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_240 br[239] vdd vss bl[239] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_240 br[239] vdd vss bl[239] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_240 br[239] vdd vss bl[239] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_240 br[239] vdd vss bl[239] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_240 br[239] vdd vss bl[239] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_240 br[239] vdd vss bl[239] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_240 br[239] vdd vss bl[239] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_240 br[239] vdd vss bl[239] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_240 br[239] vdd vss bl[239] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_240 br[239] vdd vss bl[239] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_241 br[240] vdd vss bl[240] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_241 br[240] vdd vss bl[240] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_241 br[240] vdd vss bl[240] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_241 br[240] vdd vss bl[240] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_241 br[240] vdd vss bl[240] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_241 br[240] vdd vss bl[240] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_241 br[240] vdd vss bl[240] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_241 br[240] vdd vss bl[240] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_241 br[240] vdd vss bl[240] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_241 br[240] vdd vss bl[240] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_241 br[240] vdd vss bl[240] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_241 br[240] vdd vss bl[240] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_241 br[240] vdd vss bl[240] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_241 br[240] vdd vss bl[240] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_241 br[240] vdd vss bl[240] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_241 br[240] vdd vss bl[240] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_241 br[240] vdd vss bl[240] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_241 br[240] vdd vss bl[240] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_241 br[240] vdd vss bl[240] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_242 br[241] vdd vss bl[241] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_242 br[241] vdd vss bl[241] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_242 br[241] vdd vss bl[241] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_242 br[241] vdd vss bl[241] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_242 br[241] vdd vss bl[241] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_242 br[241] vdd vss bl[241] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_242 br[241] vdd vss bl[241] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_242 br[241] vdd vss bl[241] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_242 br[241] vdd vss bl[241] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_242 br[241] vdd vss bl[241] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_242 br[241] vdd vss bl[241] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_242 br[241] vdd vss bl[241] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_242 br[241] vdd vss bl[241] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_242 br[241] vdd vss bl[241] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_242 br[241] vdd vss bl[241] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_242 br[241] vdd vss bl[241] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_242 br[241] vdd vss bl[241] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_242 br[241] vdd vss bl[241] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_242 br[241] vdd vss bl[241] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_243 br[242] vdd vss bl[242] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_243 br[242] vdd vss bl[242] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_243 br[242] vdd vss bl[242] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_243 br[242] vdd vss bl[242] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_243 br[242] vdd vss bl[242] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_243 br[242] vdd vss bl[242] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_243 br[242] vdd vss bl[242] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_243 br[242] vdd vss bl[242] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_243 br[242] vdd vss bl[242] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_243 br[242] vdd vss bl[242] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_243 br[242] vdd vss bl[242] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_243 br[242] vdd vss bl[242] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_243 br[242] vdd vss bl[242] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_243 br[242] vdd vss bl[242] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_243 br[242] vdd vss bl[242] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_243 br[242] vdd vss bl[242] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_243 br[242] vdd vss bl[242] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_243 br[242] vdd vss bl[242] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_243 br[242] vdd vss bl[242] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_244 br[243] vdd vss bl[243] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_244 br[243] vdd vss bl[243] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_244 br[243] vdd vss bl[243] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_244 br[243] vdd vss bl[243] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_244 br[243] vdd vss bl[243] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_244 br[243] vdd vss bl[243] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_244 br[243] vdd vss bl[243] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_244 br[243] vdd vss bl[243] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_244 br[243] vdd vss bl[243] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_244 br[243] vdd vss bl[243] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_244 br[243] vdd vss bl[243] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_244 br[243] vdd vss bl[243] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_244 br[243] vdd vss bl[243] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_244 br[243] vdd vss bl[243] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_244 br[243] vdd vss bl[243] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_244 br[243] vdd vss bl[243] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_244 br[243] vdd vss bl[243] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_244 br[243] vdd vss bl[243] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_244 br[243] vdd vss bl[243] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_245 br[244] vdd vss bl[244] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_245 br[244] vdd vss bl[244] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_245 br[244] vdd vss bl[244] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_245 br[244] vdd vss bl[244] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_245 br[244] vdd vss bl[244] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_245 br[244] vdd vss bl[244] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_245 br[244] vdd vss bl[244] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_245 br[244] vdd vss bl[244] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_245 br[244] vdd vss bl[244] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_245 br[244] vdd vss bl[244] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_245 br[244] vdd vss bl[244] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_245 br[244] vdd vss bl[244] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_245 br[244] vdd vss bl[244] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_245 br[244] vdd vss bl[244] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_245 br[244] vdd vss bl[244] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_245 br[244] vdd vss bl[244] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_245 br[244] vdd vss bl[244] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_245 br[244] vdd vss bl[244] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_245 br[244] vdd vss bl[244] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_246 br[245] vdd vss bl[245] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_246 br[245] vdd vss bl[245] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_246 br[245] vdd vss bl[245] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_246 br[245] vdd vss bl[245] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_246 br[245] vdd vss bl[245] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_246 br[245] vdd vss bl[245] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_246 br[245] vdd vss bl[245] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_246 br[245] vdd vss bl[245] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_246 br[245] vdd vss bl[245] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_246 br[245] vdd vss bl[245] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_246 br[245] vdd vss bl[245] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_246 br[245] vdd vss bl[245] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_246 br[245] vdd vss bl[245] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_246 br[245] vdd vss bl[245] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_246 br[245] vdd vss bl[245] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_246 br[245] vdd vss bl[245] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_246 br[245] vdd vss bl[245] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_246 br[245] vdd vss bl[245] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_246 br[245] vdd vss bl[245] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_247 br[246] vdd vss bl[246] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_247 br[246] vdd vss bl[246] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_247 br[246] vdd vss bl[246] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_247 br[246] vdd vss bl[246] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_247 br[246] vdd vss bl[246] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_247 br[246] vdd vss bl[246] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_247 br[246] vdd vss bl[246] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_247 br[246] vdd vss bl[246] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_247 br[246] vdd vss bl[246] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_247 br[246] vdd vss bl[246] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_247 br[246] vdd vss bl[246] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_247 br[246] vdd vss bl[246] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_247 br[246] vdd vss bl[246] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_247 br[246] vdd vss bl[246] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_247 br[246] vdd vss bl[246] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_247 br[246] vdd vss bl[246] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_247 br[246] vdd vss bl[246] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_247 br[246] vdd vss bl[246] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_247 br[246] vdd vss bl[246] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_248 br[247] vdd vss bl[247] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_248 br[247] vdd vss bl[247] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_248 br[247] vdd vss bl[247] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_248 br[247] vdd vss bl[247] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_248 br[247] vdd vss bl[247] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_248 br[247] vdd vss bl[247] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_248 br[247] vdd vss bl[247] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_248 br[247] vdd vss bl[247] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_248 br[247] vdd vss bl[247] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_248 br[247] vdd vss bl[247] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_248 br[247] vdd vss bl[247] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_248 br[247] vdd vss bl[247] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_248 br[247] vdd vss bl[247] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_248 br[247] vdd vss bl[247] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_248 br[247] vdd vss bl[247] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_248 br[247] vdd vss bl[247] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_248 br[247] vdd vss bl[247] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_248 br[247] vdd vss bl[247] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_248 br[247] vdd vss bl[247] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_249 br[248] vdd vss bl[248] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_249 br[248] vdd vss bl[248] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_249 br[248] vdd vss bl[248] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_249 br[248] vdd vss bl[248] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_249 br[248] vdd vss bl[248] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_249 br[248] vdd vss bl[248] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_249 br[248] vdd vss bl[248] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_249 br[248] vdd vss bl[248] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_249 br[248] vdd vss bl[248] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_249 br[248] vdd vss bl[248] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_249 br[248] vdd vss bl[248] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_249 br[248] vdd vss bl[248] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_249 br[248] vdd vss bl[248] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_249 br[248] vdd vss bl[248] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_249 br[248] vdd vss bl[248] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_249 br[248] vdd vss bl[248] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_249 br[248] vdd vss bl[248] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_249 br[248] vdd vss bl[248] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_249 br[248] vdd vss bl[248] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_250 br[249] vdd vss bl[249] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_250 br[249] vdd vss bl[249] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_250 br[249] vdd vss bl[249] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_250 br[249] vdd vss bl[249] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_250 br[249] vdd vss bl[249] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_250 br[249] vdd vss bl[249] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_250 br[249] vdd vss bl[249] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_250 br[249] vdd vss bl[249] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_250 br[249] vdd vss bl[249] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_250 br[249] vdd vss bl[249] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_250 br[249] vdd vss bl[249] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_250 br[249] vdd vss bl[249] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_250 br[249] vdd vss bl[249] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_250 br[249] vdd vss bl[249] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_250 br[249] vdd vss bl[249] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_250 br[249] vdd vss bl[249] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_250 br[249] vdd vss bl[249] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_250 br[249] vdd vss bl[249] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_250 br[249] vdd vss bl[249] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_251 br[250] vdd vss bl[250] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_251 br[250] vdd vss bl[250] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_251 br[250] vdd vss bl[250] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_251 br[250] vdd vss bl[250] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_251 br[250] vdd vss bl[250] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_251 br[250] vdd vss bl[250] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_251 br[250] vdd vss bl[250] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_251 br[250] vdd vss bl[250] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_251 br[250] vdd vss bl[250] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_251 br[250] vdd vss bl[250] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_251 br[250] vdd vss bl[250] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_251 br[250] vdd vss bl[250] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_251 br[250] vdd vss bl[250] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_251 br[250] vdd vss bl[250] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_251 br[250] vdd vss bl[250] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_251 br[250] vdd vss bl[250] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_251 br[250] vdd vss bl[250] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_251 br[250] vdd vss bl[250] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_251 br[250] vdd vss bl[250] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_252 br[251] vdd vss bl[251] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_252 br[251] vdd vss bl[251] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_252 br[251] vdd vss bl[251] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_252 br[251] vdd vss bl[251] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_252 br[251] vdd vss bl[251] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_252 br[251] vdd vss bl[251] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_252 br[251] vdd vss bl[251] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_252 br[251] vdd vss bl[251] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_252 br[251] vdd vss bl[251] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_252 br[251] vdd vss bl[251] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_252 br[251] vdd vss bl[251] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_252 br[251] vdd vss bl[251] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_252 br[251] vdd vss bl[251] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_252 br[251] vdd vss bl[251] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_252 br[251] vdd vss bl[251] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_252 br[251] vdd vss bl[251] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_252 br[251] vdd vss bl[251] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_252 br[251] vdd vss bl[251] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_252 br[251] vdd vss bl[251] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_253 br[252] vdd vss bl[252] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_253 br[252] vdd vss bl[252] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_253 br[252] vdd vss bl[252] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_253 br[252] vdd vss bl[252] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_253 br[252] vdd vss bl[252] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_253 br[252] vdd vss bl[252] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_253 br[252] vdd vss bl[252] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_253 br[252] vdd vss bl[252] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_253 br[252] vdd vss bl[252] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_253 br[252] vdd vss bl[252] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_253 br[252] vdd vss bl[252] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_253 br[252] vdd vss bl[252] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_253 br[252] vdd vss bl[252] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_253 br[252] vdd vss bl[252] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_253 br[252] vdd vss bl[252] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_253 br[252] vdd vss bl[252] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_253 br[252] vdd vss bl[252] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_253 br[252] vdd vss bl[252] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_253 br[252] vdd vss bl[252] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_254 br[253] vdd vss bl[253] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_254 br[253] vdd vss bl[253] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_254 br[253] vdd vss bl[253] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_254 br[253] vdd vss bl[253] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_254 br[253] vdd vss bl[253] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_254 br[253] vdd vss bl[253] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_254 br[253] vdd vss bl[253] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_254 br[253] vdd vss bl[253] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_254 br[253] vdd vss bl[253] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_254 br[253] vdd vss bl[253] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_254 br[253] vdd vss bl[253] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_254 br[253] vdd vss bl[253] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_254 br[253] vdd vss bl[253] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_254 br[253] vdd vss bl[253] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_254 br[253] vdd vss bl[253] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_254 br[253] vdd vss bl[253] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_254 br[253] vdd vss bl[253] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_254 br[253] vdd vss bl[253] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_254 br[253] vdd vss bl[253] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_255 br[254] vdd vss bl[254] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_255 br[254] vdd vss bl[254] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_255 br[254] vdd vss bl[254] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_255 br[254] vdd vss bl[254] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_255 br[254] vdd vss bl[254] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_255 br[254] vdd vss bl[254] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_255 br[254] vdd vss bl[254] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_255 br[254] vdd vss bl[254] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_255 br[254] vdd vss bl[254] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_255 br[254] vdd vss bl[254] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_255 br[254] vdd vss bl[254] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_255 br[254] vdd vss bl[254] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_255 br[254] vdd vss bl[254] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_255 br[254] vdd vss bl[254] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_255 br[254] vdd vss bl[254] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_255 br[254] vdd vss bl[254] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_255 br[254] vdd vss bl[254] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_255 br[254] vdd vss bl[254] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_255 br[254] vdd vss bl[254] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_256 br[255] vdd vss bl[255] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_256 br[255] vdd vss bl[255] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_256 br[255] vdd vss bl[255] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_256 br[255] vdd vss bl[255] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_256 br[255] vdd vss bl[255] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_256 br[255] vdd vss bl[255] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_256 br[255] vdd vss bl[255] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_256 br[255] vdd vss bl[255] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_256 br[255] vdd vss bl[255] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_256 br[255] vdd vss bl[255] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_256 br[255] vdd vss bl[255] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_256 br[255] vdd vss bl[255] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_256 br[255] vdd vss bl[255] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_256 br[255] vdd vss bl[255] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_256 br[255] vdd vss bl[255] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_256 br[255] vdd vss bl[255] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_256 br[255] vdd vss bl[255] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_256 br[255] vdd vss bl[255] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_256 br[255] vdd vss bl[255] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_257 br[256] vdd vss bl[256] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_257 br[256] vdd vss bl[256] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_257 br[256] vdd vss bl[256] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_257 br[256] vdd vss bl[256] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_257 br[256] vdd vss bl[256] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_257 br[256] vdd vss bl[256] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_257 br[256] vdd vss bl[256] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_257 br[256] vdd vss bl[256] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_257 br[256] vdd vss bl[256] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_257 br[256] vdd vss bl[256] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_257 br[256] vdd vss bl[256] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_257 br[256] vdd vss bl[256] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_257 br[256] vdd vss bl[256] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_257 br[256] vdd vss bl[256] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_257 br[256] vdd vss bl[256] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_257 br[256] vdd vss bl[256] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_257 br[256] vdd vss bl[256] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_257 br[256] vdd vss bl[256] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_257 br[256] vdd vss bl[256] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_258 br[257] vdd vss bl[257] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_258 br[257] vdd vss bl[257] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_258 br[257] vdd vss bl[257] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_258 br[257] vdd vss bl[257] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_258 br[257] vdd vss bl[257] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_258 br[257] vdd vss bl[257] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_258 br[257] vdd vss bl[257] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_258 br[257] vdd vss bl[257] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_258 br[257] vdd vss bl[257] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_258 br[257] vdd vss bl[257] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_258 br[257] vdd vss bl[257] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_258 br[257] vdd vss bl[257] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_258 br[257] vdd vss bl[257] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_258 br[257] vdd vss bl[257] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_258 br[257] vdd vss bl[257] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_258 br[257] vdd vss bl[257] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_258 br[257] vdd vss bl[257] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_258 br[257] vdd vss bl[257] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_258 br[257] vdd vss bl[257] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_259 br[258] vdd vss bl[258] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_259 br[258] vdd vss bl[258] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_259 br[258] vdd vss bl[258] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_259 br[258] vdd vss bl[258] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_259 br[258] vdd vss bl[258] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_259 br[258] vdd vss bl[258] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_259 br[258] vdd vss bl[258] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_259 br[258] vdd vss bl[258] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_259 br[258] vdd vss bl[258] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_259 br[258] vdd vss bl[258] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_259 br[258] vdd vss bl[258] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_259 br[258] vdd vss bl[258] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_259 br[258] vdd vss bl[258] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_259 br[258] vdd vss bl[258] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_259 br[258] vdd vss bl[258] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_259 br[258] vdd vss bl[258] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_259 br[258] vdd vss bl[258] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_259 br[258] vdd vss bl[258] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_259 br[258] vdd vss bl[258] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_260 br[259] vdd vss bl[259] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_260 br[259] vdd vss bl[259] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_260 br[259] vdd vss bl[259] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_260 br[259] vdd vss bl[259] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_260 br[259] vdd vss bl[259] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_260 br[259] vdd vss bl[259] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_260 br[259] vdd vss bl[259] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_260 br[259] vdd vss bl[259] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_260 br[259] vdd vss bl[259] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_260 br[259] vdd vss bl[259] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_260 br[259] vdd vss bl[259] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_260 br[259] vdd vss bl[259] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_260 br[259] vdd vss bl[259] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_260 br[259] vdd vss bl[259] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_260 br[259] vdd vss bl[259] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_260 br[259] vdd vss bl[259] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_260 br[259] vdd vss bl[259] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_260 br[259] vdd vss bl[259] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_260 br[259] vdd vss bl[259] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_261 br[260] vdd vss bl[260] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_261 br[260] vdd vss bl[260] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_261 br[260] vdd vss bl[260] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_261 br[260] vdd vss bl[260] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_261 br[260] vdd vss bl[260] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_261 br[260] vdd vss bl[260] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_261 br[260] vdd vss bl[260] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_261 br[260] vdd vss bl[260] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_261 br[260] vdd vss bl[260] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_261 br[260] vdd vss bl[260] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_261 br[260] vdd vss bl[260] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_261 br[260] vdd vss bl[260] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_261 br[260] vdd vss bl[260] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_261 br[260] vdd vss bl[260] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_261 br[260] vdd vss bl[260] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_261 br[260] vdd vss bl[260] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_261 br[260] vdd vss bl[260] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_261 br[260] vdd vss bl[260] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_261 br[260] vdd vss bl[260] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_262 br[261] vdd vss bl[261] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_262 br[261] vdd vss bl[261] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_262 br[261] vdd vss bl[261] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_262 br[261] vdd vss bl[261] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_262 br[261] vdd vss bl[261] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_262 br[261] vdd vss bl[261] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_262 br[261] vdd vss bl[261] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_262 br[261] vdd vss bl[261] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_262 br[261] vdd vss bl[261] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_262 br[261] vdd vss bl[261] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_262 br[261] vdd vss bl[261] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_262 br[261] vdd vss bl[261] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_262 br[261] vdd vss bl[261] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_262 br[261] vdd vss bl[261] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_262 br[261] vdd vss bl[261] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_262 br[261] vdd vss bl[261] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_262 br[261] vdd vss bl[261] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_262 br[261] vdd vss bl[261] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_262 br[261] vdd vss bl[261] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_263 br[262] vdd vss bl[262] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_263 br[262] vdd vss bl[262] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_263 br[262] vdd vss bl[262] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_263 br[262] vdd vss bl[262] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_263 br[262] vdd vss bl[262] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_263 br[262] vdd vss bl[262] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_263 br[262] vdd vss bl[262] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_263 br[262] vdd vss bl[262] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_263 br[262] vdd vss bl[262] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_263 br[262] vdd vss bl[262] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_263 br[262] vdd vss bl[262] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_263 br[262] vdd vss bl[262] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_263 br[262] vdd vss bl[262] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_263 br[262] vdd vss bl[262] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_263 br[262] vdd vss bl[262] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_263 br[262] vdd vss bl[262] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_263 br[262] vdd vss bl[262] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_263 br[262] vdd vss bl[262] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_263 br[262] vdd vss bl[262] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_264 br[263] vdd vss bl[263] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_264 br[263] vdd vss bl[263] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_264 br[263] vdd vss bl[263] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_264 br[263] vdd vss bl[263] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_264 br[263] vdd vss bl[263] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_264 br[263] vdd vss bl[263] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_264 br[263] vdd vss bl[263] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_264 br[263] vdd vss bl[263] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_264 br[263] vdd vss bl[263] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_264 br[263] vdd vss bl[263] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_264 br[263] vdd vss bl[263] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_264 br[263] vdd vss bl[263] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_264 br[263] vdd vss bl[263] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_264 br[263] vdd vss bl[263] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_264 br[263] vdd vss bl[263] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_264 br[263] vdd vss bl[263] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_264 br[263] vdd vss bl[263] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_264 br[263] vdd vss bl[263] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_264 br[263] vdd vss bl[263] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_265 br[264] vdd vss bl[264] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_265 br[264] vdd vss bl[264] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_265 br[264] vdd vss bl[264] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_265 br[264] vdd vss bl[264] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_265 br[264] vdd vss bl[264] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_265 br[264] vdd vss bl[264] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_265 br[264] vdd vss bl[264] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_265 br[264] vdd vss bl[264] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_265 br[264] vdd vss bl[264] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_265 br[264] vdd vss bl[264] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_265 br[264] vdd vss bl[264] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_265 br[264] vdd vss bl[264] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_265 br[264] vdd vss bl[264] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_265 br[264] vdd vss bl[264] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_265 br[264] vdd vss bl[264] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_265 br[264] vdd vss bl[264] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_265 br[264] vdd vss bl[264] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_265 br[264] vdd vss bl[264] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_265 br[264] vdd vss bl[264] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_266 br[265] vdd vss bl[265] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_266 br[265] vdd vss bl[265] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_266 br[265] vdd vss bl[265] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_266 br[265] vdd vss bl[265] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_266 br[265] vdd vss bl[265] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_266 br[265] vdd vss bl[265] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_266 br[265] vdd vss bl[265] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_266 br[265] vdd vss bl[265] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_266 br[265] vdd vss bl[265] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_266 br[265] vdd vss bl[265] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_266 br[265] vdd vss bl[265] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_266 br[265] vdd vss bl[265] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_266 br[265] vdd vss bl[265] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_266 br[265] vdd vss bl[265] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_266 br[265] vdd vss bl[265] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_266 br[265] vdd vss bl[265] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_266 br[265] vdd vss bl[265] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_266 br[265] vdd vss bl[265] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_266 br[265] vdd vss bl[265] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_267 br[266] vdd vss bl[266] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_267 br[266] vdd vss bl[266] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_267 br[266] vdd vss bl[266] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_267 br[266] vdd vss bl[266] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_267 br[266] vdd vss bl[266] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_267 br[266] vdd vss bl[266] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_267 br[266] vdd vss bl[266] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_267 br[266] vdd vss bl[266] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_267 br[266] vdd vss bl[266] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_267 br[266] vdd vss bl[266] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_267 br[266] vdd vss bl[266] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_267 br[266] vdd vss bl[266] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_267 br[266] vdd vss bl[266] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_267 br[266] vdd vss bl[266] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_267 br[266] vdd vss bl[266] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_267 br[266] vdd vss bl[266] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_267 br[266] vdd vss bl[266] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_267 br[266] vdd vss bl[266] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_267 br[266] vdd vss bl[266] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_268 br[267] vdd vss bl[267] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_268 br[267] vdd vss bl[267] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_268 br[267] vdd vss bl[267] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_268 br[267] vdd vss bl[267] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_268 br[267] vdd vss bl[267] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_268 br[267] vdd vss bl[267] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_268 br[267] vdd vss bl[267] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_268 br[267] vdd vss bl[267] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_268 br[267] vdd vss bl[267] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_268 br[267] vdd vss bl[267] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_268 br[267] vdd vss bl[267] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_268 br[267] vdd vss bl[267] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_268 br[267] vdd vss bl[267] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_268 br[267] vdd vss bl[267] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_268 br[267] vdd vss bl[267] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_268 br[267] vdd vss bl[267] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_268 br[267] vdd vss bl[267] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_268 br[267] vdd vss bl[267] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_268 br[267] vdd vss bl[267] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_269 br[268] vdd vss bl[268] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_269 br[268] vdd vss bl[268] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_269 br[268] vdd vss bl[268] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_269 br[268] vdd vss bl[268] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_269 br[268] vdd vss bl[268] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_269 br[268] vdd vss bl[268] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_269 br[268] vdd vss bl[268] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_269 br[268] vdd vss bl[268] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_269 br[268] vdd vss bl[268] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_269 br[268] vdd vss bl[268] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_269 br[268] vdd vss bl[268] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_269 br[268] vdd vss bl[268] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_269 br[268] vdd vss bl[268] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_269 br[268] vdd vss bl[268] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_269 br[268] vdd vss bl[268] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_269 br[268] vdd vss bl[268] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_269 br[268] vdd vss bl[268] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_269 br[268] vdd vss bl[268] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_269 br[268] vdd vss bl[268] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_270 br[269] vdd vss bl[269] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_270 br[269] vdd vss bl[269] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_270 br[269] vdd vss bl[269] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_270 br[269] vdd vss bl[269] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_270 br[269] vdd vss bl[269] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_270 br[269] vdd vss bl[269] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_270 br[269] vdd vss bl[269] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_270 br[269] vdd vss bl[269] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_270 br[269] vdd vss bl[269] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_270 br[269] vdd vss bl[269] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_270 br[269] vdd vss bl[269] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_270 br[269] vdd vss bl[269] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_270 br[269] vdd vss bl[269] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_270 br[269] vdd vss bl[269] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_270 br[269] vdd vss bl[269] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_270 br[269] vdd vss bl[269] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_270 br[269] vdd vss bl[269] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_270 br[269] vdd vss bl[269] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_270 br[269] vdd vss bl[269] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_271 br[270] vdd vss bl[270] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_271 br[270] vdd vss bl[270] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_271 br[270] vdd vss bl[270] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_271 br[270] vdd vss bl[270] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_271 br[270] vdd vss bl[270] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_271 br[270] vdd vss bl[270] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_271 br[270] vdd vss bl[270] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_271 br[270] vdd vss bl[270] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_271 br[270] vdd vss bl[270] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_271 br[270] vdd vss bl[270] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_271 br[270] vdd vss bl[270] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_271 br[270] vdd vss bl[270] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_271 br[270] vdd vss bl[270] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_271 br[270] vdd vss bl[270] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_271 br[270] vdd vss bl[270] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_271 br[270] vdd vss bl[270] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_271 br[270] vdd vss bl[270] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_271 br[270] vdd vss bl[270] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_271 br[270] vdd vss bl[270] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_272 br[271] vdd vss bl[271] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_272 br[271] vdd vss bl[271] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_272 br[271] vdd vss bl[271] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_272 br[271] vdd vss bl[271] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_272 br[271] vdd vss bl[271] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_272 br[271] vdd vss bl[271] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_272 br[271] vdd vss bl[271] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_272 br[271] vdd vss bl[271] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_272 br[271] vdd vss bl[271] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_272 br[271] vdd vss bl[271] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_272 br[271] vdd vss bl[271] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_272 br[271] vdd vss bl[271] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_272 br[271] vdd vss bl[271] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_272 br[271] vdd vss bl[271] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_272 br[271] vdd vss bl[271] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_272 br[271] vdd vss bl[271] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_272 br[271] vdd vss bl[271] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_272 br[271] vdd vss bl[271] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_272 br[271] vdd vss bl[271] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_273 br[272] vdd vss bl[272] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_273 br[272] vdd vss bl[272] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_273 br[272] vdd vss bl[272] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_273 br[272] vdd vss bl[272] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_273 br[272] vdd vss bl[272] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_273 br[272] vdd vss bl[272] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_273 br[272] vdd vss bl[272] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_273 br[272] vdd vss bl[272] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_273 br[272] vdd vss bl[272] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_273 br[272] vdd vss bl[272] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_273 br[272] vdd vss bl[272] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_273 br[272] vdd vss bl[272] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_273 br[272] vdd vss bl[272] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_273 br[272] vdd vss bl[272] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_273 br[272] vdd vss bl[272] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_273 br[272] vdd vss bl[272] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_273 br[272] vdd vss bl[272] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_273 br[272] vdd vss bl[272] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_273 br[272] vdd vss bl[272] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_274 br[273] vdd vss bl[273] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_274 br[273] vdd vss bl[273] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_274 br[273] vdd vss bl[273] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_274 br[273] vdd vss bl[273] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_274 br[273] vdd vss bl[273] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_274 br[273] vdd vss bl[273] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_274 br[273] vdd vss bl[273] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_274 br[273] vdd vss bl[273] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_274 br[273] vdd vss bl[273] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_274 br[273] vdd vss bl[273] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_274 br[273] vdd vss bl[273] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_274 br[273] vdd vss bl[273] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_274 br[273] vdd vss bl[273] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_274 br[273] vdd vss bl[273] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_274 br[273] vdd vss bl[273] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_274 br[273] vdd vss bl[273] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_274 br[273] vdd vss bl[273] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_274 br[273] vdd vss bl[273] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_274 br[273] vdd vss bl[273] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_275 br[274] vdd vss bl[274] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_275 br[274] vdd vss bl[274] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_275 br[274] vdd vss bl[274] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_275 br[274] vdd vss bl[274] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_275 br[274] vdd vss bl[274] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_275 br[274] vdd vss bl[274] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_275 br[274] vdd vss bl[274] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_275 br[274] vdd vss bl[274] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_275 br[274] vdd vss bl[274] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_275 br[274] vdd vss bl[274] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_275 br[274] vdd vss bl[274] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_275 br[274] vdd vss bl[274] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_275 br[274] vdd vss bl[274] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_275 br[274] vdd vss bl[274] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_275 br[274] vdd vss bl[274] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_275 br[274] vdd vss bl[274] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_275 br[274] vdd vss bl[274] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_275 br[274] vdd vss bl[274] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_275 br[274] vdd vss bl[274] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_276 br[275] vdd vss bl[275] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_276 br[275] vdd vss bl[275] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_276 br[275] vdd vss bl[275] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_276 br[275] vdd vss bl[275] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_276 br[275] vdd vss bl[275] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_276 br[275] vdd vss bl[275] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_276 br[275] vdd vss bl[275] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_276 br[275] vdd vss bl[275] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_276 br[275] vdd vss bl[275] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_276 br[275] vdd vss bl[275] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_276 br[275] vdd vss bl[275] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_276 br[275] vdd vss bl[275] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_276 br[275] vdd vss bl[275] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_276 br[275] vdd vss bl[275] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_276 br[275] vdd vss bl[275] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_276 br[275] vdd vss bl[275] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_276 br[275] vdd vss bl[275] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_276 br[275] vdd vss bl[275] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_276 br[275] vdd vss bl[275] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_277 br[276] vdd vss bl[276] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_277 br[276] vdd vss bl[276] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_277 br[276] vdd vss bl[276] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_277 br[276] vdd vss bl[276] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_277 br[276] vdd vss bl[276] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_277 br[276] vdd vss bl[276] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_277 br[276] vdd vss bl[276] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_277 br[276] vdd vss bl[276] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_277 br[276] vdd vss bl[276] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_277 br[276] vdd vss bl[276] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_277 br[276] vdd vss bl[276] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_277 br[276] vdd vss bl[276] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_277 br[276] vdd vss bl[276] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_277 br[276] vdd vss bl[276] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_277 br[276] vdd vss bl[276] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_277 br[276] vdd vss bl[276] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_277 br[276] vdd vss bl[276] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_277 br[276] vdd vss bl[276] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_277 br[276] vdd vss bl[276] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_278 br[277] vdd vss bl[277] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_278 br[277] vdd vss bl[277] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_278 br[277] vdd vss bl[277] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_278 br[277] vdd vss bl[277] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_278 br[277] vdd vss bl[277] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_278 br[277] vdd vss bl[277] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_278 br[277] vdd vss bl[277] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_278 br[277] vdd vss bl[277] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_278 br[277] vdd vss bl[277] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_278 br[277] vdd vss bl[277] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_278 br[277] vdd vss bl[277] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_278 br[277] vdd vss bl[277] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_278 br[277] vdd vss bl[277] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_278 br[277] vdd vss bl[277] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_278 br[277] vdd vss bl[277] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_278 br[277] vdd vss bl[277] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_278 br[277] vdd vss bl[277] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_278 br[277] vdd vss bl[277] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_278 br[277] vdd vss bl[277] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_279 br[278] vdd vss bl[278] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_279 br[278] vdd vss bl[278] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_279 br[278] vdd vss bl[278] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_279 br[278] vdd vss bl[278] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_279 br[278] vdd vss bl[278] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_279 br[278] vdd vss bl[278] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_279 br[278] vdd vss bl[278] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_279 br[278] vdd vss bl[278] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_279 br[278] vdd vss bl[278] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_279 br[278] vdd vss bl[278] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_279 br[278] vdd vss bl[278] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_279 br[278] vdd vss bl[278] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_279 br[278] vdd vss bl[278] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_279 br[278] vdd vss bl[278] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_279 br[278] vdd vss bl[278] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_279 br[278] vdd vss bl[278] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_279 br[278] vdd vss bl[278] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_279 br[278] vdd vss bl[278] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_279 br[278] vdd vss bl[278] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_280 br[279] vdd vss bl[279] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_280 br[279] vdd vss bl[279] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_280 br[279] vdd vss bl[279] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_280 br[279] vdd vss bl[279] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_280 br[279] vdd vss bl[279] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_280 br[279] vdd vss bl[279] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_280 br[279] vdd vss bl[279] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_280 br[279] vdd vss bl[279] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_280 br[279] vdd vss bl[279] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_280 br[279] vdd vss bl[279] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_280 br[279] vdd vss bl[279] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_280 br[279] vdd vss bl[279] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_280 br[279] vdd vss bl[279] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_280 br[279] vdd vss bl[279] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_280 br[279] vdd vss bl[279] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_280 br[279] vdd vss bl[279] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_280 br[279] vdd vss bl[279] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_280 br[279] vdd vss bl[279] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_280 br[279] vdd vss bl[279] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_281 br[280] vdd vss bl[280] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_281 br[280] vdd vss bl[280] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_281 br[280] vdd vss bl[280] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_281 br[280] vdd vss bl[280] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_281 br[280] vdd vss bl[280] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_281 br[280] vdd vss bl[280] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_281 br[280] vdd vss bl[280] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_281 br[280] vdd vss bl[280] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_281 br[280] vdd vss bl[280] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_281 br[280] vdd vss bl[280] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_281 br[280] vdd vss bl[280] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_281 br[280] vdd vss bl[280] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_281 br[280] vdd vss bl[280] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_281 br[280] vdd vss bl[280] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_281 br[280] vdd vss bl[280] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_281 br[280] vdd vss bl[280] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_281 br[280] vdd vss bl[280] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_281 br[280] vdd vss bl[280] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_281 br[280] vdd vss bl[280] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_282 br[281] vdd vss bl[281] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_282 br[281] vdd vss bl[281] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_282 br[281] vdd vss bl[281] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_282 br[281] vdd vss bl[281] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_282 br[281] vdd vss bl[281] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_282 br[281] vdd vss bl[281] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_282 br[281] vdd vss bl[281] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_282 br[281] vdd vss bl[281] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_282 br[281] vdd vss bl[281] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_282 br[281] vdd vss bl[281] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_282 br[281] vdd vss bl[281] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_282 br[281] vdd vss bl[281] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_282 br[281] vdd vss bl[281] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_282 br[281] vdd vss bl[281] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_282 br[281] vdd vss bl[281] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_282 br[281] vdd vss bl[281] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_282 br[281] vdd vss bl[281] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_282 br[281] vdd vss bl[281] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_282 br[281] vdd vss bl[281] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_283 br[282] vdd vss bl[282] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_283 br[282] vdd vss bl[282] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_283 br[282] vdd vss bl[282] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_283 br[282] vdd vss bl[282] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_283 br[282] vdd vss bl[282] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_283 br[282] vdd vss bl[282] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_283 br[282] vdd vss bl[282] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_283 br[282] vdd vss bl[282] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_283 br[282] vdd vss bl[282] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_283 br[282] vdd vss bl[282] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_283 br[282] vdd vss bl[282] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_283 br[282] vdd vss bl[282] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_283 br[282] vdd vss bl[282] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_283 br[282] vdd vss bl[282] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_283 br[282] vdd vss bl[282] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_283 br[282] vdd vss bl[282] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_283 br[282] vdd vss bl[282] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_283 br[282] vdd vss bl[282] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_283 br[282] vdd vss bl[282] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_284 br[283] vdd vss bl[283] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_284 br[283] vdd vss bl[283] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_284 br[283] vdd vss bl[283] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_284 br[283] vdd vss bl[283] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_284 br[283] vdd vss bl[283] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_284 br[283] vdd vss bl[283] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_284 br[283] vdd vss bl[283] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_284 br[283] vdd vss bl[283] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_284 br[283] vdd vss bl[283] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_284 br[283] vdd vss bl[283] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_284 br[283] vdd vss bl[283] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_284 br[283] vdd vss bl[283] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_284 br[283] vdd vss bl[283] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_284 br[283] vdd vss bl[283] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_284 br[283] vdd vss bl[283] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_284 br[283] vdd vss bl[283] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_284 br[283] vdd vss bl[283] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_284 br[283] vdd vss bl[283] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_284 br[283] vdd vss bl[283] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_285 br[284] vdd vss bl[284] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_285 br[284] vdd vss bl[284] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_285 br[284] vdd vss bl[284] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_285 br[284] vdd vss bl[284] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_285 br[284] vdd vss bl[284] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_285 br[284] vdd vss bl[284] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_285 br[284] vdd vss bl[284] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_285 br[284] vdd vss bl[284] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_285 br[284] vdd vss bl[284] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_285 br[284] vdd vss bl[284] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_285 br[284] vdd vss bl[284] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_285 br[284] vdd vss bl[284] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_285 br[284] vdd vss bl[284] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_285 br[284] vdd vss bl[284] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_285 br[284] vdd vss bl[284] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_285 br[284] vdd vss bl[284] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_285 br[284] vdd vss bl[284] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_285 br[284] vdd vss bl[284] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_285 br[284] vdd vss bl[284] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_286 br[285] vdd vss bl[285] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_286 br[285] vdd vss bl[285] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_286 br[285] vdd vss bl[285] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_286 br[285] vdd vss bl[285] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_286 br[285] vdd vss bl[285] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_286 br[285] vdd vss bl[285] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_286 br[285] vdd vss bl[285] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_286 br[285] vdd vss bl[285] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_286 br[285] vdd vss bl[285] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_286 br[285] vdd vss bl[285] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_286 br[285] vdd vss bl[285] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_286 br[285] vdd vss bl[285] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_286 br[285] vdd vss bl[285] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_286 br[285] vdd vss bl[285] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_286 br[285] vdd vss bl[285] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_286 br[285] vdd vss bl[285] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_286 br[285] vdd vss bl[285] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_286 br[285] vdd vss bl[285] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_286 br[285] vdd vss bl[285] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_287 br[286] vdd vss bl[286] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_287 br[286] vdd vss bl[286] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_287 br[286] vdd vss bl[286] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_287 br[286] vdd vss bl[286] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_287 br[286] vdd vss bl[286] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_287 br[286] vdd vss bl[286] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_287 br[286] vdd vss bl[286] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_287 br[286] vdd vss bl[286] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_287 br[286] vdd vss bl[286] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_287 br[286] vdd vss bl[286] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_287 br[286] vdd vss bl[286] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_287 br[286] vdd vss bl[286] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_287 br[286] vdd vss bl[286] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_287 br[286] vdd vss bl[286] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_287 br[286] vdd vss bl[286] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_287 br[286] vdd vss bl[286] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_287 br[286] vdd vss bl[286] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_287 br[286] vdd vss bl[286] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_287 br[286] vdd vss bl[286] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_288 br[287] vdd vss bl[287] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_288 br[287] vdd vss bl[287] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_288 br[287] vdd vss bl[287] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_288 br[287] vdd vss bl[287] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_288 br[287] vdd vss bl[287] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_288 br[287] vdd vss bl[287] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_288 br[287] vdd vss bl[287] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_288 br[287] vdd vss bl[287] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_288 br[287] vdd vss bl[287] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_288 br[287] vdd vss bl[287] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_288 br[287] vdd vss bl[287] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_288 br[287] vdd vss bl[287] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_288 br[287] vdd vss bl[287] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_288 br[287] vdd vss bl[287] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_288 br[287] vdd vss bl[287] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_288 br[287] vdd vss bl[287] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_288 br[287] vdd vss bl[287] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_288 br[287] vdd vss bl[287] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_288 br[287] vdd vss bl[287] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_289 br[288] vdd vss bl[288] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_289 br[288] vdd vss bl[288] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_289 br[288] vdd vss bl[288] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_289 br[288] vdd vss bl[288] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_289 br[288] vdd vss bl[288] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_289 br[288] vdd vss bl[288] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_289 br[288] vdd vss bl[288] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_289 br[288] vdd vss bl[288] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_289 br[288] vdd vss bl[288] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_289 br[288] vdd vss bl[288] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_289 br[288] vdd vss bl[288] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_289 br[288] vdd vss bl[288] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_289 br[288] vdd vss bl[288] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_289 br[288] vdd vss bl[288] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_289 br[288] vdd vss bl[288] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_289 br[288] vdd vss bl[288] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_289 br[288] vdd vss bl[288] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_289 br[288] vdd vss bl[288] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_289 br[288] vdd vss bl[288] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_290 br[289] vdd vss bl[289] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_290 br[289] vdd vss bl[289] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_290 br[289] vdd vss bl[289] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_290 br[289] vdd vss bl[289] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_290 br[289] vdd vss bl[289] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_290 br[289] vdd vss bl[289] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_290 br[289] vdd vss bl[289] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_290 br[289] vdd vss bl[289] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_290 br[289] vdd vss bl[289] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_290 br[289] vdd vss bl[289] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_290 br[289] vdd vss bl[289] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_290 br[289] vdd vss bl[289] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_290 br[289] vdd vss bl[289] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_290 br[289] vdd vss bl[289] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_290 br[289] vdd vss bl[289] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_290 br[289] vdd vss bl[289] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_290 br[289] vdd vss bl[289] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_290 br[289] vdd vss bl[289] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_290 br[289] vdd vss bl[289] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_291 br[290] vdd vss bl[290] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_291 br[290] vdd vss bl[290] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_291 br[290] vdd vss bl[290] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_291 br[290] vdd vss bl[290] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_291 br[290] vdd vss bl[290] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_291 br[290] vdd vss bl[290] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_291 br[290] vdd vss bl[290] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_291 br[290] vdd vss bl[290] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_291 br[290] vdd vss bl[290] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_291 br[290] vdd vss bl[290] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_291 br[290] vdd vss bl[290] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_291 br[290] vdd vss bl[290] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_291 br[290] vdd vss bl[290] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_291 br[290] vdd vss bl[290] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_291 br[290] vdd vss bl[290] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_291 br[290] vdd vss bl[290] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_291 br[290] vdd vss bl[290] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_291 br[290] vdd vss bl[290] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_291 br[290] vdd vss bl[290] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_292 br[291] vdd vss bl[291] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_292 br[291] vdd vss bl[291] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_292 br[291] vdd vss bl[291] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_292 br[291] vdd vss bl[291] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_292 br[291] vdd vss bl[291] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_292 br[291] vdd vss bl[291] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_292 br[291] vdd vss bl[291] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_292 br[291] vdd vss bl[291] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_292 br[291] vdd vss bl[291] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_292 br[291] vdd vss bl[291] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_292 br[291] vdd vss bl[291] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_292 br[291] vdd vss bl[291] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_292 br[291] vdd vss bl[291] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_292 br[291] vdd vss bl[291] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_292 br[291] vdd vss bl[291] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_292 br[291] vdd vss bl[291] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_292 br[291] vdd vss bl[291] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_292 br[291] vdd vss bl[291] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_292 br[291] vdd vss bl[291] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_293 br[292] vdd vss bl[292] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_293 br[292] vdd vss bl[292] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_293 br[292] vdd vss bl[292] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_293 br[292] vdd vss bl[292] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_293 br[292] vdd vss bl[292] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_293 br[292] vdd vss bl[292] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_293 br[292] vdd vss bl[292] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_293 br[292] vdd vss bl[292] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_293 br[292] vdd vss bl[292] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_293 br[292] vdd vss bl[292] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_293 br[292] vdd vss bl[292] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_293 br[292] vdd vss bl[292] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_293 br[292] vdd vss bl[292] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_293 br[292] vdd vss bl[292] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_293 br[292] vdd vss bl[292] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_293 br[292] vdd vss bl[292] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_293 br[292] vdd vss bl[292] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_293 br[292] vdd vss bl[292] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_293 br[292] vdd vss bl[292] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_294 br[293] vdd vss bl[293] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_294 br[293] vdd vss bl[293] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_294 br[293] vdd vss bl[293] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_294 br[293] vdd vss bl[293] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_294 br[293] vdd vss bl[293] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_294 br[293] vdd vss bl[293] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_294 br[293] vdd vss bl[293] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_294 br[293] vdd vss bl[293] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_294 br[293] vdd vss bl[293] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_294 br[293] vdd vss bl[293] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_294 br[293] vdd vss bl[293] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_294 br[293] vdd vss bl[293] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_294 br[293] vdd vss bl[293] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_294 br[293] vdd vss bl[293] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_294 br[293] vdd vss bl[293] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_294 br[293] vdd vss bl[293] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_294 br[293] vdd vss bl[293] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_294 br[293] vdd vss bl[293] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_294 br[293] vdd vss bl[293] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_295 br[294] vdd vss bl[294] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_295 br[294] vdd vss bl[294] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_295 br[294] vdd vss bl[294] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_295 br[294] vdd vss bl[294] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_295 br[294] vdd vss bl[294] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_295 br[294] vdd vss bl[294] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_295 br[294] vdd vss bl[294] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_295 br[294] vdd vss bl[294] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_295 br[294] vdd vss bl[294] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_295 br[294] vdd vss bl[294] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_295 br[294] vdd vss bl[294] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_295 br[294] vdd vss bl[294] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_295 br[294] vdd vss bl[294] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_295 br[294] vdd vss bl[294] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_295 br[294] vdd vss bl[294] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_295 br[294] vdd vss bl[294] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_295 br[294] vdd vss bl[294] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_295 br[294] vdd vss bl[294] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_295 br[294] vdd vss bl[294] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_296 br[295] vdd vss bl[295] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_296 br[295] vdd vss bl[295] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_296 br[295] vdd vss bl[295] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_296 br[295] vdd vss bl[295] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_296 br[295] vdd vss bl[295] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_296 br[295] vdd vss bl[295] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_296 br[295] vdd vss bl[295] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_296 br[295] vdd vss bl[295] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_296 br[295] vdd vss bl[295] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_296 br[295] vdd vss bl[295] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_296 br[295] vdd vss bl[295] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_296 br[295] vdd vss bl[295] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_296 br[295] vdd vss bl[295] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_296 br[295] vdd vss bl[295] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_296 br[295] vdd vss bl[295] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_296 br[295] vdd vss bl[295] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_296 br[295] vdd vss bl[295] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_296 br[295] vdd vss bl[295] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_296 br[295] vdd vss bl[295] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_297 br[296] vdd vss bl[296] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_297 br[296] vdd vss bl[296] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_297 br[296] vdd vss bl[296] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_297 br[296] vdd vss bl[296] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_297 br[296] vdd vss bl[296] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_297 br[296] vdd vss bl[296] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_297 br[296] vdd vss bl[296] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_297 br[296] vdd vss bl[296] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_297 br[296] vdd vss bl[296] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_297 br[296] vdd vss bl[296] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_297 br[296] vdd vss bl[296] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_297 br[296] vdd vss bl[296] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_297 br[296] vdd vss bl[296] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_297 br[296] vdd vss bl[296] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_297 br[296] vdd vss bl[296] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_297 br[296] vdd vss bl[296] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_297 br[296] vdd vss bl[296] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_297 br[296] vdd vss bl[296] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_297 br[296] vdd vss bl[296] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_298 br[297] vdd vss bl[297] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_298 br[297] vdd vss bl[297] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_298 br[297] vdd vss bl[297] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_298 br[297] vdd vss bl[297] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_298 br[297] vdd vss bl[297] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_298 br[297] vdd vss bl[297] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_298 br[297] vdd vss bl[297] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_298 br[297] vdd vss bl[297] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_298 br[297] vdd vss bl[297] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_298 br[297] vdd vss bl[297] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_298 br[297] vdd vss bl[297] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_298 br[297] vdd vss bl[297] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_298 br[297] vdd vss bl[297] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_298 br[297] vdd vss bl[297] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_298 br[297] vdd vss bl[297] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_298 br[297] vdd vss bl[297] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_298 br[297] vdd vss bl[297] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_298 br[297] vdd vss bl[297] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_298 br[297] vdd vss bl[297] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_299 br[298] vdd vss bl[298] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_299 br[298] vdd vss bl[298] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_299 br[298] vdd vss bl[298] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_299 br[298] vdd vss bl[298] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_299 br[298] vdd vss bl[298] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_299 br[298] vdd vss bl[298] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_299 br[298] vdd vss bl[298] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_299 br[298] vdd vss bl[298] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_299 br[298] vdd vss bl[298] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_299 br[298] vdd vss bl[298] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_299 br[298] vdd vss bl[298] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_299 br[298] vdd vss bl[298] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_299 br[298] vdd vss bl[298] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_299 br[298] vdd vss bl[298] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_299 br[298] vdd vss bl[298] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_299 br[298] vdd vss bl[298] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_299 br[298] vdd vss bl[298] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_299 br[298] vdd vss bl[298] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_299 br[298] vdd vss bl[298] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_300 br[299] vdd vss bl[299] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_300 br[299] vdd vss bl[299] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_300 br[299] vdd vss bl[299] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_300 br[299] vdd vss bl[299] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_300 br[299] vdd vss bl[299] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_300 br[299] vdd vss bl[299] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_300 br[299] vdd vss bl[299] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_300 br[299] vdd vss bl[299] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_300 br[299] vdd vss bl[299] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_300 br[299] vdd vss bl[299] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_300 br[299] vdd vss bl[299] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_300 br[299] vdd vss bl[299] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_300 br[299] vdd vss bl[299] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_300 br[299] vdd vss bl[299] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_300 br[299] vdd vss bl[299] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_300 br[299] vdd vss bl[299] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_300 br[299] vdd vss bl[299] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_300 br[299] vdd vss bl[299] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_300 br[299] vdd vss bl[299] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_301 br[300] vdd vss bl[300] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_301 br[300] vdd vss bl[300] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_301 br[300] vdd vss bl[300] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_301 br[300] vdd vss bl[300] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_301 br[300] vdd vss bl[300] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_301 br[300] vdd vss bl[300] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_301 br[300] vdd vss bl[300] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_301 br[300] vdd vss bl[300] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_301 br[300] vdd vss bl[300] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_301 br[300] vdd vss bl[300] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_301 br[300] vdd vss bl[300] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_301 br[300] vdd vss bl[300] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_301 br[300] vdd vss bl[300] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_301 br[300] vdd vss bl[300] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_301 br[300] vdd vss bl[300] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_301 br[300] vdd vss bl[300] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_301 br[300] vdd vss bl[300] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_301 br[300] vdd vss bl[300] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_301 br[300] vdd vss bl[300] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_302 br[301] vdd vss bl[301] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_302 br[301] vdd vss bl[301] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_302 br[301] vdd vss bl[301] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_302 br[301] vdd vss bl[301] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_302 br[301] vdd vss bl[301] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_302 br[301] vdd vss bl[301] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_302 br[301] vdd vss bl[301] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_302 br[301] vdd vss bl[301] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_302 br[301] vdd vss bl[301] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_302 br[301] vdd vss bl[301] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_302 br[301] vdd vss bl[301] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_302 br[301] vdd vss bl[301] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_302 br[301] vdd vss bl[301] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_302 br[301] vdd vss bl[301] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_302 br[301] vdd vss bl[301] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_302 br[301] vdd vss bl[301] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_302 br[301] vdd vss bl[301] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_302 br[301] vdd vss bl[301] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_302 br[301] vdd vss bl[301] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_303 br[302] vdd vss bl[302] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_303 br[302] vdd vss bl[302] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_303 br[302] vdd vss bl[302] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_303 br[302] vdd vss bl[302] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_303 br[302] vdd vss bl[302] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_303 br[302] vdd vss bl[302] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_303 br[302] vdd vss bl[302] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_303 br[302] vdd vss bl[302] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_303 br[302] vdd vss bl[302] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_303 br[302] vdd vss bl[302] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_303 br[302] vdd vss bl[302] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_303 br[302] vdd vss bl[302] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_303 br[302] vdd vss bl[302] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_303 br[302] vdd vss bl[302] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_303 br[302] vdd vss bl[302] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_303 br[302] vdd vss bl[302] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_303 br[302] vdd vss bl[302] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_303 br[302] vdd vss bl[302] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_303 br[302] vdd vss bl[302] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_304 br[303] vdd vss bl[303] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_304 br[303] vdd vss bl[303] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_304 br[303] vdd vss bl[303] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_304 br[303] vdd vss bl[303] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_304 br[303] vdd vss bl[303] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_304 br[303] vdd vss bl[303] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_304 br[303] vdd vss bl[303] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_304 br[303] vdd vss bl[303] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_304 br[303] vdd vss bl[303] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_304 br[303] vdd vss bl[303] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_304 br[303] vdd vss bl[303] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_304 br[303] vdd vss bl[303] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_304 br[303] vdd vss bl[303] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_304 br[303] vdd vss bl[303] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_304 br[303] vdd vss bl[303] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_304 br[303] vdd vss bl[303] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_304 br[303] vdd vss bl[303] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_304 br[303] vdd vss bl[303] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_304 br[303] vdd vss bl[303] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_305 br[304] vdd vss bl[304] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_305 br[304] vdd vss bl[304] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_305 br[304] vdd vss bl[304] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_305 br[304] vdd vss bl[304] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_305 br[304] vdd vss bl[304] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_305 br[304] vdd vss bl[304] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_305 br[304] vdd vss bl[304] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_305 br[304] vdd vss bl[304] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_305 br[304] vdd vss bl[304] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_305 br[304] vdd vss bl[304] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_305 br[304] vdd vss bl[304] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_305 br[304] vdd vss bl[304] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_305 br[304] vdd vss bl[304] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_305 br[304] vdd vss bl[304] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_305 br[304] vdd vss bl[304] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_305 br[304] vdd vss bl[304] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_305 br[304] vdd vss bl[304] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_305 br[304] vdd vss bl[304] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_305 br[304] vdd vss bl[304] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_306 br[305] vdd vss bl[305] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_306 br[305] vdd vss bl[305] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_306 br[305] vdd vss bl[305] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_306 br[305] vdd vss bl[305] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_306 br[305] vdd vss bl[305] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_306 br[305] vdd vss bl[305] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_306 br[305] vdd vss bl[305] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_306 br[305] vdd vss bl[305] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_306 br[305] vdd vss bl[305] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_306 br[305] vdd vss bl[305] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_306 br[305] vdd vss bl[305] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_306 br[305] vdd vss bl[305] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_306 br[305] vdd vss bl[305] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_306 br[305] vdd vss bl[305] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_306 br[305] vdd vss bl[305] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_306 br[305] vdd vss bl[305] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_306 br[305] vdd vss bl[305] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_306 br[305] vdd vss bl[305] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_306 br[305] vdd vss bl[305] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_307 br[306] vdd vss bl[306] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_307 br[306] vdd vss bl[306] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_307 br[306] vdd vss bl[306] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_307 br[306] vdd vss bl[306] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_307 br[306] vdd vss bl[306] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_307 br[306] vdd vss bl[306] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_307 br[306] vdd vss bl[306] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_307 br[306] vdd vss bl[306] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_307 br[306] vdd vss bl[306] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_307 br[306] vdd vss bl[306] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_307 br[306] vdd vss bl[306] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_307 br[306] vdd vss bl[306] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_307 br[306] vdd vss bl[306] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_307 br[306] vdd vss bl[306] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_307 br[306] vdd vss bl[306] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_307 br[306] vdd vss bl[306] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_307 br[306] vdd vss bl[306] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_307 br[306] vdd vss bl[306] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_307 br[306] vdd vss bl[306] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_308 br[307] vdd vss bl[307] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_308 br[307] vdd vss bl[307] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_308 br[307] vdd vss bl[307] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_308 br[307] vdd vss bl[307] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_308 br[307] vdd vss bl[307] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_308 br[307] vdd vss bl[307] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_308 br[307] vdd vss bl[307] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_308 br[307] vdd vss bl[307] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_308 br[307] vdd vss bl[307] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_308 br[307] vdd vss bl[307] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_308 br[307] vdd vss bl[307] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_308 br[307] vdd vss bl[307] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_308 br[307] vdd vss bl[307] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_308 br[307] vdd vss bl[307] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_308 br[307] vdd vss bl[307] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_308 br[307] vdd vss bl[307] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_308 br[307] vdd vss bl[307] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_308 br[307] vdd vss bl[307] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_308 br[307] vdd vss bl[307] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_309 br[308] vdd vss bl[308] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_309 br[308] vdd vss bl[308] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_309 br[308] vdd vss bl[308] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_309 br[308] vdd vss bl[308] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_309 br[308] vdd vss bl[308] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_309 br[308] vdd vss bl[308] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_309 br[308] vdd vss bl[308] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_309 br[308] vdd vss bl[308] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_309 br[308] vdd vss bl[308] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_309 br[308] vdd vss bl[308] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_309 br[308] vdd vss bl[308] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_309 br[308] vdd vss bl[308] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_309 br[308] vdd vss bl[308] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_309 br[308] vdd vss bl[308] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_309 br[308] vdd vss bl[308] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_309 br[308] vdd vss bl[308] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_309 br[308] vdd vss bl[308] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_309 br[308] vdd vss bl[308] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_309 br[308] vdd vss bl[308] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_310 br[309] vdd vss bl[309] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_310 br[309] vdd vss bl[309] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_310 br[309] vdd vss bl[309] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_310 br[309] vdd vss bl[309] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_310 br[309] vdd vss bl[309] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_310 br[309] vdd vss bl[309] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_310 br[309] vdd vss bl[309] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_310 br[309] vdd vss bl[309] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_310 br[309] vdd vss bl[309] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_310 br[309] vdd vss bl[309] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_310 br[309] vdd vss bl[309] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_310 br[309] vdd vss bl[309] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_310 br[309] vdd vss bl[309] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_310 br[309] vdd vss bl[309] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_310 br[309] vdd vss bl[309] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_310 br[309] vdd vss bl[309] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_310 br[309] vdd vss bl[309] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_310 br[309] vdd vss bl[309] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_310 br[309] vdd vss bl[309] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_311 br[310] vdd vss bl[310] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_311 br[310] vdd vss bl[310] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_311 br[310] vdd vss bl[310] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_311 br[310] vdd vss bl[310] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_311 br[310] vdd vss bl[310] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_311 br[310] vdd vss bl[310] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_311 br[310] vdd vss bl[310] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_311 br[310] vdd vss bl[310] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_311 br[310] vdd vss bl[310] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_311 br[310] vdd vss bl[310] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_311 br[310] vdd vss bl[310] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_311 br[310] vdd vss bl[310] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_311 br[310] vdd vss bl[310] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_311 br[310] vdd vss bl[310] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_311 br[310] vdd vss bl[310] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_311 br[310] vdd vss bl[310] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_311 br[310] vdd vss bl[310] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_311 br[310] vdd vss bl[310] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_311 br[310] vdd vss bl[310] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_312 br[311] vdd vss bl[311] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_312 br[311] vdd vss bl[311] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_312 br[311] vdd vss bl[311] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_312 br[311] vdd vss bl[311] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_312 br[311] vdd vss bl[311] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_312 br[311] vdd vss bl[311] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_312 br[311] vdd vss bl[311] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_312 br[311] vdd vss bl[311] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_312 br[311] vdd vss bl[311] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_312 br[311] vdd vss bl[311] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_312 br[311] vdd vss bl[311] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_312 br[311] vdd vss bl[311] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_312 br[311] vdd vss bl[311] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_312 br[311] vdd vss bl[311] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_312 br[311] vdd vss bl[311] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_312 br[311] vdd vss bl[311] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_312 br[311] vdd vss bl[311] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_312 br[311] vdd vss bl[311] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_312 br[311] vdd vss bl[311] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_313 br[312] vdd vss bl[312] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_313 br[312] vdd vss bl[312] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_313 br[312] vdd vss bl[312] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_313 br[312] vdd vss bl[312] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_313 br[312] vdd vss bl[312] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_313 br[312] vdd vss bl[312] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_313 br[312] vdd vss bl[312] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_313 br[312] vdd vss bl[312] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_313 br[312] vdd vss bl[312] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_313 br[312] vdd vss bl[312] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_313 br[312] vdd vss bl[312] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_313 br[312] vdd vss bl[312] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_313 br[312] vdd vss bl[312] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_313 br[312] vdd vss bl[312] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_313 br[312] vdd vss bl[312] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_313 br[312] vdd vss bl[312] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_313 br[312] vdd vss bl[312] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_313 br[312] vdd vss bl[312] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_313 br[312] vdd vss bl[312] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_314 br[313] vdd vss bl[313] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_314 br[313] vdd vss bl[313] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_314 br[313] vdd vss bl[313] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_314 br[313] vdd vss bl[313] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_314 br[313] vdd vss bl[313] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_314 br[313] vdd vss bl[313] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_314 br[313] vdd vss bl[313] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_314 br[313] vdd vss bl[313] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_314 br[313] vdd vss bl[313] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_314 br[313] vdd vss bl[313] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_314 br[313] vdd vss bl[313] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_314 br[313] vdd vss bl[313] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_314 br[313] vdd vss bl[313] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_314 br[313] vdd vss bl[313] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_314 br[313] vdd vss bl[313] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_314 br[313] vdd vss bl[313] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_314 br[313] vdd vss bl[313] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_314 br[313] vdd vss bl[313] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_314 br[313] vdd vss bl[313] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_315 br[314] vdd vss bl[314] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_315 br[314] vdd vss bl[314] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_315 br[314] vdd vss bl[314] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_315 br[314] vdd vss bl[314] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_315 br[314] vdd vss bl[314] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_315 br[314] vdd vss bl[314] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_315 br[314] vdd vss bl[314] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_315 br[314] vdd vss bl[314] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_315 br[314] vdd vss bl[314] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_315 br[314] vdd vss bl[314] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_315 br[314] vdd vss bl[314] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_315 br[314] vdd vss bl[314] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_315 br[314] vdd vss bl[314] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_315 br[314] vdd vss bl[314] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_315 br[314] vdd vss bl[314] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_315 br[314] vdd vss bl[314] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_315 br[314] vdd vss bl[314] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_315 br[314] vdd vss bl[314] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_315 br[314] vdd vss bl[314] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_316 br[315] vdd vss bl[315] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_316 br[315] vdd vss bl[315] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_316 br[315] vdd vss bl[315] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_316 br[315] vdd vss bl[315] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_316 br[315] vdd vss bl[315] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_316 br[315] vdd vss bl[315] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_316 br[315] vdd vss bl[315] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_316 br[315] vdd vss bl[315] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_316 br[315] vdd vss bl[315] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_316 br[315] vdd vss bl[315] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_316 br[315] vdd vss bl[315] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_316 br[315] vdd vss bl[315] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_316 br[315] vdd vss bl[315] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_316 br[315] vdd vss bl[315] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_316 br[315] vdd vss bl[315] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_316 br[315] vdd vss bl[315] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_316 br[315] vdd vss bl[315] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_316 br[315] vdd vss bl[315] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_316 br[315] vdd vss bl[315] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_317 br[316] vdd vss bl[316] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_317 br[316] vdd vss bl[316] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_317 br[316] vdd vss bl[316] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_317 br[316] vdd vss bl[316] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_317 br[316] vdd vss bl[316] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_317 br[316] vdd vss bl[316] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_317 br[316] vdd vss bl[316] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_317 br[316] vdd vss bl[316] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_317 br[316] vdd vss bl[316] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_317 br[316] vdd vss bl[316] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_317 br[316] vdd vss bl[316] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_317 br[316] vdd vss bl[316] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_317 br[316] vdd vss bl[316] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_317 br[316] vdd vss bl[316] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_317 br[316] vdd vss bl[316] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_317 br[316] vdd vss bl[316] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_317 br[316] vdd vss bl[316] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_317 br[316] vdd vss bl[316] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_317 br[316] vdd vss bl[316] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_318 br[317] vdd vss bl[317] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_318 br[317] vdd vss bl[317] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_318 br[317] vdd vss bl[317] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_318 br[317] vdd vss bl[317] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_318 br[317] vdd vss bl[317] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_318 br[317] vdd vss bl[317] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_318 br[317] vdd vss bl[317] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_318 br[317] vdd vss bl[317] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_318 br[317] vdd vss bl[317] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_318 br[317] vdd vss bl[317] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_318 br[317] vdd vss bl[317] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_318 br[317] vdd vss bl[317] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_318 br[317] vdd vss bl[317] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_318 br[317] vdd vss bl[317] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_318 br[317] vdd vss bl[317] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_318 br[317] vdd vss bl[317] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_318 br[317] vdd vss bl[317] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_318 br[317] vdd vss bl[317] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_318 br[317] vdd vss bl[317] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_319 br[318] vdd vss bl[318] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_319 br[318] vdd vss bl[318] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_319 br[318] vdd vss bl[318] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_319 br[318] vdd vss bl[318] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_319 br[318] vdd vss bl[318] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_319 br[318] vdd vss bl[318] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_319 br[318] vdd vss bl[318] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_319 br[318] vdd vss bl[318] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_319 br[318] vdd vss bl[318] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_319 br[318] vdd vss bl[318] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_319 br[318] vdd vss bl[318] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_319 br[318] vdd vss bl[318] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_319 br[318] vdd vss bl[318] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_319 br[318] vdd vss bl[318] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_319 br[318] vdd vss bl[318] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_319 br[318] vdd vss bl[318] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_319 br[318] vdd vss bl[318] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_319 br[318] vdd vss bl[318] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_319 br[318] vdd vss bl[318] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_320 br[319] vdd vss bl[319] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_320 br[319] vdd vss bl[319] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_320 br[319] vdd vss bl[319] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_320 br[319] vdd vss bl[319] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_320 br[319] vdd vss bl[319] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_320 br[319] vdd vss bl[319] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_320 br[319] vdd vss bl[319] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_320 br[319] vdd vss bl[319] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_320 br[319] vdd vss bl[319] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_320 br[319] vdd vss bl[319] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_320 br[319] vdd vss bl[319] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_320 br[319] vdd vss bl[319] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_320 br[319] vdd vss bl[319] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_320 br[319] vdd vss bl[319] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_320 br[319] vdd vss bl[319] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_320 br[319] vdd vss bl[319] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_320 br[319] vdd vss bl[319] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_320 br[319] vdd vss bl[319] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_320 br[319] vdd vss bl[319] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_321 br[320] vdd vss bl[320] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_321 br[320] vdd vss bl[320] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_321 br[320] vdd vss bl[320] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_321 br[320] vdd vss bl[320] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_321 br[320] vdd vss bl[320] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_321 br[320] vdd vss bl[320] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_321 br[320] vdd vss bl[320] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_321 br[320] vdd vss bl[320] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_321 br[320] vdd vss bl[320] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_321 br[320] vdd vss bl[320] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_321 br[320] vdd vss bl[320] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_321 br[320] vdd vss bl[320] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_321 br[320] vdd vss bl[320] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_321 br[320] vdd vss bl[320] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_321 br[320] vdd vss bl[320] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_321 br[320] vdd vss bl[320] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_321 br[320] vdd vss bl[320] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_321 br[320] vdd vss bl[320] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_321 br[320] vdd vss bl[320] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_322 br[321] vdd vss bl[321] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_322 br[321] vdd vss bl[321] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_322 br[321] vdd vss bl[321] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_322 br[321] vdd vss bl[321] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_322 br[321] vdd vss bl[321] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_322 br[321] vdd vss bl[321] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_322 br[321] vdd vss bl[321] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_322 br[321] vdd vss bl[321] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_322 br[321] vdd vss bl[321] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_322 br[321] vdd vss bl[321] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_322 br[321] vdd vss bl[321] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_322 br[321] vdd vss bl[321] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_322 br[321] vdd vss bl[321] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_322 br[321] vdd vss bl[321] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_322 br[321] vdd vss bl[321] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_322 br[321] vdd vss bl[321] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_322 br[321] vdd vss bl[321] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_322 br[321] vdd vss bl[321] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_322 br[321] vdd vss bl[321] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_323 br[322] vdd vss bl[322] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_323 br[322] vdd vss bl[322] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_323 br[322] vdd vss bl[322] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_323 br[322] vdd vss bl[322] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_323 br[322] vdd vss bl[322] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_323 br[322] vdd vss bl[322] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_323 br[322] vdd vss bl[322] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_323 br[322] vdd vss bl[322] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_323 br[322] vdd vss bl[322] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_323 br[322] vdd vss bl[322] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_323 br[322] vdd vss bl[322] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_323 br[322] vdd vss bl[322] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_323 br[322] vdd vss bl[322] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_323 br[322] vdd vss bl[322] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_323 br[322] vdd vss bl[322] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_323 br[322] vdd vss bl[322] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_323 br[322] vdd vss bl[322] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_323 br[322] vdd vss bl[322] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_323 br[322] vdd vss bl[322] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_324 br[323] vdd vss bl[323] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_324 br[323] vdd vss bl[323] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_324 br[323] vdd vss bl[323] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_324 br[323] vdd vss bl[323] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_324 br[323] vdd vss bl[323] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_324 br[323] vdd vss bl[323] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_324 br[323] vdd vss bl[323] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_324 br[323] vdd vss bl[323] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_324 br[323] vdd vss bl[323] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_324 br[323] vdd vss bl[323] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_324 br[323] vdd vss bl[323] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_324 br[323] vdd vss bl[323] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_324 br[323] vdd vss bl[323] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_324 br[323] vdd vss bl[323] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_324 br[323] vdd vss bl[323] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_324 br[323] vdd vss bl[323] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_324 br[323] vdd vss bl[323] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_324 br[323] vdd vss bl[323] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_324 br[323] vdd vss bl[323] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_325 br[324] vdd vss bl[324] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_325 br[324] vdd vss bl[324] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_325 br[324] vdd vss bl[324] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_325 br[324] vdd vss bl[324] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_325 br[324] vdd vss bl[324] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_325 br[324] vdd vss bl[324] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_325 br[324] vdd vss bl[324] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_325 br[324] vdd vss bl[324] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_325 br[324] vdd vss bl[324] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_325 br[324] vdd vss bl[324] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_325 br[324] vdd vss bl[324] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_325 br[324] vdd vss bl[324] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_325 br[324] vdd vss bl[324] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_325 br[324] vdd vss bl[324] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_325 br[324] vdd vss bl[324] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_325 br[324] vdd vss bl[324] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_325 br[324] vdd vss bl[324] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_325 br[324] vdd vss bl[324] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_325 br[324] vdd vss bl[324] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_326 br[325] vdd vss bl[325] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_326 br[325] vdd vss bl[325] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_326 br[325] vdd vss bl[325] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_326 br[325] vdd vss bl[325] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_326 br[325] vdd vss bl[325] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_326 br[325] vdd vss bl[325] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_326 br[325] vdd vss bl[325] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_326 br[325] vdd vss bl[325] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_326 br[325] vdd vss bl[325] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_326 br[325] vdd vss bl[325] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_326 br[325] vdd vss bl[325] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_326 br[325] vdd vss bl[325] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_326 br[325] vdd vss bl[325] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_326 br[325] vdd vss bl[325] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_326 br[325] vdd vss bl[325] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_326 br[325] vdd vss bl[325] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_326 br[325] vdd vss bl[325] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_326 br[325] vdd vss bl[325] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_326 br[325] vdd vss bl[325] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_327 br[326] vdd vss bl[326] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_327 br[326] vdd vss bl[326] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_327 br[326] vdd vss bl[326] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_327 br[326] vdd vss bl[326] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_327 br[326] vdd vss bl[326] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_327 br[326] vdd vss bl[326] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_327 br[326] vdd vss bl[326] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_327 br[326] vdd vss bl[326] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_327 br[326] vdd vss bl[326] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_327 br[326] vdd vss bl[326] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_327 br[326] vdd vss bl[326] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_327 br[326] vdd vss bl[326] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_327 br[326] vdd vss bl[326] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_327 br[326] vdd vss bl[326] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_327 br[326] vdd vss bl[326] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_327 br[326] vdd vss bl[326] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_327 br[326] vdd vss bl[326] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_327 br[326] vdd vss bl[326] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_327 br[326] vdd vss bl[326] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_328 br[327] vdd vss bl[327] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_328 br[327] vdd vss bl[327] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_328 br[327] vdd vss bl[327] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_328 br[327] vdd vss bl[327] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_328 br[327] vdd vss bl[327] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_328 br[327] vdd vss bl[327] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_328 br[327] vdd vss bl[327] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_328 br[327] vdd vss bl[327] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_328 br[327] vdd vss bl[327] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_328 br[327] vdd vss bl[327] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_328 br[327] vdd vss bl[327] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_328 br[327] vdd vss bl[327] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_328 br[327] vdd vss bl[327] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_328 br[327] vdd vss bl[327] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_328 br[327] vdd vss bl[327] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_328 br[327] vdd vss bl[327] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_328 br[327] vdd vss bl[327] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_328 br[327] vdd vss bl[327] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_328 br[327] vdd vss bl[327] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_329 br[328] vdd vss bl[328] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_329 br[328] vdd vss bl[328] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_329 br[328] vdd vss bl[328] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_329 br[328] vdd vss bl[328] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_329 br[328] vdd vss bl[328] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_329 br[328] vdd vss bl[328] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_329 br[328] vdd vss bl[328] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_329 br[328] vdd vss bl[328] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_329 br[328] vdd vss bl[328] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_329 br[328] vdd vss bl[328] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_329 br[328] vdd vss bl[328] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_329 br[328] vdd vss bl[328] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_329 br[328] vdd vss bl[328] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_329 br[328] vdd vss bl[328] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_329 br[328] vdd vss bl[328] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_329 br[328] vdd vss bl[328] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_329 br[328] vdd vss bl[328] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_329 br[328] vdd vss bl[328] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_329 br[328] vdd vss bl[328] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_330 br[329] vdd vss bl[329] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_330 br[329] vdd vss bl[329] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_330 br[329] vdd vss bl[329] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_330 br[329] vdd vss bl[329] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_330 br[329] vdd vss bl[329] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_330 br[329] vdd vss bl[329] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_330 br[329] vdd vss bl[329] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_330 br[329] vdd vss bl[329] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_330 br[329] vdd vss bl[329] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_330 br[329] vdd vss bl[329] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_330 br[329] vdd vss bl[329] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_330 br[329] vdd vss bl[329] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_330 br[329] vdd vss bl[329] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_330 br[329] vdd vss bl[329] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_330 br[329] vdd vss bl[329] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_330 br[329] vdd vss bl[329] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_330 br[329] vdd vss bl[329] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_330 br[329] vdd vss bl[329] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_330 br[329] vdd vss bl[329] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_331 br[330] vdd vss bl[330] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_331 br[330] vdd vss bl[330] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_331 br[330] vdd vss bl[330] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_331 br[330] vdd vss bl[330] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_331 br[330] vdd vss bl[330] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_331 br[330] vdd vss bl[330] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_331 br[330] vdd vss bl[330] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_331 br[330] vdd vss bl[330] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_331 br[330] vdd vss bl[330] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_331 br[330] vdd vss bl[330] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_331 br[330] vdd vss bl[330] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_331 br[330] vdd vss bl[330] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_331 br[330] vdd vss bl[330] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_331 br[330] vdd vss bl[330] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_331 br[330] vdd vss bl[330] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_331 br[330] vdd vss bl[330] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_331 br[330] vdd vss bl[330] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_331 br[330] vdd vss bl[330] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_331 br[330] vdd vss bl[330] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_332 br[331] vdd vss bl[331] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_332 br[331] vdd vss bl[331] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_332 br[331] vdd vss bl[331] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_332 br[331] vdd vss bl[331] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_332 br[331] vdd vss bl[331] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_332 br[331] vdd vss bl[331] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_332 br[331] vdd vss bl[331] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_332 br[331] vdd vss bl[331] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_332 br[331] vdd vss bl[331] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_332 br[331] vdd vss bl[331] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_332 br[331] vdd vss bl[331] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_332 br[331] vdd vss bl[331] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_332 br[331] vdd vss bl[331] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_332 br[331] vdd vss bl[331] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_332 br[331] vdd vss bl[331] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_332 br[331] vdd vss bl[331] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_332 br[331] vdd vss bl[331] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_332 br[331] vdd vss bl[331] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_332 br[331] vdd vss bl[331] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_333 br[332] vdd vss bl[332] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_333 br[332] vdd vss bl[332] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_333 br[332] vdd vss bl[332] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_333 br[332] vdd vss bl[332] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_333 br[332] vdd vss bl[332] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_333 br[332] vdd vss bl[332] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_333 br[332] vdd vss bl[332] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_333 br[332] vdd vss bl[332] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_333 br[332] vdd vss bl[332] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_333 br[332] vdd vss bl[332] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_333 br[332] vdd vss bl[332] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_333 br[332] vdd vss bl[332] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_333 br[332] vdd vss bl[332] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_333 br[332] vdd vss bl[332] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_333 br[332] vdd vss bl[332] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_333 br[332] vdd vss bl[332] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_333 br[332] vdd vss bl[332] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_333 br[332] vdd vss bl[332] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_333 br[332] vdd vss bl[332] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_334 br[333] vdd vss bl[333] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_334 br[333] vdd vss bl[333] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_334 br[333] vdd vss bl[333] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_334 br[333] vdd vss bl[333] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_334 br[333] vdd vss bl[333] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_334 br[333] vdd vss bl[333] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_334 br[333] vdd vss bl[333] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_334 br[333] vdd vss bl[333] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_334 br[333] vdd vss bl[333] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_334 br[333] vdd vss bl[333] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_334 br[333] vdd vss bl[333] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_334 br[333] vdd vss bl[333] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_334 br[333] vdd vss bl[333] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_334 br[333] vdd vss bl[333] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_334 br[333] vdd vss bl[333] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_334 br[333] vdd vss bl[333] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_334 br[333] vdd vss bl[333] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_334 br[333] vdd vss bl[333] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_334 br[333] vdd vss bl[333] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_335 br[334] vdd vss bl[334] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_335 br[334] vdd vss bl[334] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_335 br[334] vdd vss bl[334] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_335 br[334] vdd vss bl[334] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_335 br[334] vdd vss bl[334] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_335 br[334] vdd vss bl[334] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_335 br[334] vdd vss bl[334] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_335 br[334] vdd vss bl[334] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_335 br[334] vdd vss bl[334] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_335 br[334] vdd vss bl[334] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_335 br[334] vdd vss bl[334] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_335 br[334] vdd vss bl[334] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_335 br[334] vdd vss bl[334] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_335 br[334] vdd vss bl[334] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_335 br[334] vdd vss bl[334] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_335 br[334] vdd vss bl[334] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_335 br[334] vdd vss bl[334] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_335 br[334] vdd vss bl[334] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_335 br[334] vdd vss bl[334] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_336 br[335] vdd vss bl[335] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_336 br[335] vdd vss bl[335] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_336 br[335] vdd vss bl[335] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_336 br[335] vdd vss bl[335] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_336 br[335] vdd vss bl[335] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_336 br[335] vdd vss bl[335] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_336 br[335] vdd vss bl[335] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_336 br[335] vdd vss bl[335] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_336 br[335] vdd vss bl[335] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_336 br[335] vdd vss bl[335] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_336 br[335] vdd vss bl[335] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_336 br[335] vdd vss bl[335] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_336 br[335] vdd vss bl[335] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_336 br[335] vdd vss bl[335] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_336 br[335] vdd vss bl[335] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_336 br[335] vdd vss bl[335] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_336 br[335] vdd vss bl[335] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_336 br[335] vdd vss bl[335] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_336 br[335] vdd vss bl[335] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_337 br[336] vdd vss bl[336] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_337 br[336] vdd vss bl[336] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_337 br[336] vdd vss bl[336] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_337 br[336] vdd vss bl[336] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_337 br[336] vdd vss bl[336] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_337 br[336] vdd vss bl[336] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_337 br[336] vdd vss bl[336] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_337 br[336] vdd vss bl[336] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_337 br[336] vdd vss bl[336] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_337 br[336] vdd vss bl[336] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_337 br[336] vdd vss bl[336] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_337 br[336] vdd vss bl[336] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_337 br[336] vdd vss bl[336] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_337 br[336] vdd vss bl[336] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_337 br[336] vdd vss bl[336] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_337 br[336] vdd vss bl[336] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_337 br[336] vdd vss bl[336] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_337 br[336] vdd vss bl[336] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_337 br[336] vdd vss bl[336] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_338 br[337] vdd vss bl[337] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_338 br[337] vdd vss bl[337] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_338 br[337] vdd vss bl[337] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_338 br[337] vdd vss bl[337] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_338 br[337] vdd vss bl[337] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_338 br[337] vdd vss bl[337] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_338 br[337] vdd vss bl[337] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_338 br[337] vdd vss bl[337] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_338 br[337] vdd vss bl[337] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_338 br[337] vdd vss bl[337] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_338 br[337] vdd vss bl[337] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_338 br[337] vdd vss bl[337] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_338 br[337] vdd vss bl[337] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_338 br[337] vdd vss bl[337] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_338 br[337] vdd vss bl[337] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_338 br[337] vdd vss bl[337] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_338 br[337] vdd vss bl[337] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_338 br[337] vdd vss bl[337] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_338 br[337] vdd vss bl[337] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_339 br[338] vdd vss bl[338] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_339 br[338] vdd vss bl[338] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_339 br[338] vdd vss bl[338] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_339 br[338] vdd vss bl[338] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_339 br[338] vdd vss bl[338] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_339 br[338] vdd vss bl[338] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_339 br[338] vdd vss bl[338] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_339 br[338] vdd vss bl[338] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_339 br[338] vdd vss bl[338] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_339 br[338] vdd vss bl[338] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_339 br[338] vdd vss bl[338] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_339 br[338] vdd vss bl[338] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_339 br[338] vdd vss bl[338] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_339 br[338] vdd vss bl[338] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_339 br[338] vdd vss bl[338] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_339 br[338] vdd vss bl[338] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_339 br[338] vdd vss bl[338] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_339 br[338] vdd vss bl[338] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_339 br[338] vdd vss bl[338] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_340 br[339] vdd vss bl[339] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_340 br[339] vdd vss bl[339] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_340 br[339] vdd vss bl[339] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_340 br[339] vdd vss bl[339] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_340 br[339] vdd vss bl[339] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_340 br[339] vdd vss bl[339] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_340 br[339] vdd vss bl[339] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_340 br[339] vdd vss bl[339] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_340 br[339] vdd vss bl[339] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_340 br[339] vdd vss bl[339] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_340 br[339] vdd vss bl[339] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_340 br[339] vdd vss bl[339] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_340 br[339] vdd vss bl[339] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_340 br[339] vdd vss bl[339] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_340 br[339] vdd vss bl[339] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_340 br[339] vdd vss bl[339] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_340 br[339] vdd vss bl[339] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_340 br[339] vdd vss bl[339] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_340 br[339] vdd vss bl[339] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_341 br[340] vdd vss bl[340] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_341 br[340] vdd vss bl[340] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_341 br[340] vdd vss bl[340] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_341 br[340] vdd vss bl[340] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_341 br[340] vdd vss bl[340] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_341 br[340] vdd vss bl[340] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_341 br[340] vdd vss bl[340] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_341 br[340] vdd vss bl[340] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_341 br[340] vdd vss bl[340] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_341 br[340] vdd vss bl[340] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_341 br[340] vdd vss bl[340] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_341 br[340] vdd vss bl[340] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_341 br[340] vdd vss bl[340] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_341 br[340] vdd vss bl[340] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_341 br[340] vdd vss bl[340] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_341 br[340] vdd vss bl[340] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_341 br[340] vdd vss bl[340] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_341 br[340] vdd vss bl[340] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_341 br[340] vdd vss bl[340] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_342 br[341] vdd vss bl[341] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_342 br[341] vdd vss bl[341] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_342 br[341] vdd vss bl[341] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_342 br[341] vdd vss bl[341] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_342 br[341] vdd vss bl[341] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_342 br[341] vdd vss bl[341] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_342 br[341] vdd vss bl[341] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_342 br[341] vdd vss bl[341] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_342 br[341] vdd vss bl[341] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_342 br[341] vdd vss bl[341] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_342 br[341] vdd vss bl[341] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_342 br[341] vdd vss bl[341] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_342 br[341] vdd vss bl[341] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_342 br[341] vdd vss bl[341] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_342 br[341] vdd vss bl[341] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_342 br[341] vdd vss bl[341] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_342 br[341] vdd vss bl[341] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_342 br[341] vdd vss bl[341] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_342 br[341] vdd vss bl[341] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_343 br[342] vdd vss bl[342] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_343 br[342] vdd vss bl[342] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_343 br[342] vdd vss bl[342] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_343 br[342] vdd vss bl[342] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_343 br[342] vdd vss bl[342] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_343 br[342] vdd vss bl[342] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_343 br[342] vdd vss bl[342] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_343 br[342] vdd vss bl[342] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_343 br[342] vdd vss bl[342] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_343 br[342] vdd vss bl[342] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_343 br[342] vdd vss bl[342] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_343 br[342] vdd vss bl[342] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_343 br[342] vdd vss bl[342] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_343 br[342] vdd vss bl[342] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_343 br[342] vdd vss bl[342] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_343 br[342] vdd vss bl[342] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_343 br[342] vdd vss bl[342] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_343 br[342] vdd vss bl[342] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_343 br[342] vdd vss bl[342] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_344 br[343] vdd vss bl[343] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_344 br[343] vdd vss bl[343] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_344 br[343] vdd vss bl[343] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_344 br[343] vdd vss bl[343] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_344 br[343] vdd vss bl[343] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_344 br[343] vdd vss bl[343] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_344 br[343] vdd vss bl[343] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_344 br[343] vdd vss bl[343] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_344 br[343] vdd vss bl[343] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_344 br[343] vdd vss bl[343] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_344 br[343] vdd vss bl[343] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_344 br[343] vdd vss bl[343] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_344 br[343] vdd vss bl[343] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_344 br[343] vdd vss bl[343] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_344 br[343] vdd vss bl[343] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_344 br[343] vdd vss bl[343] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_344 br[343] vdd vss bl[343] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_344 br[343] vdd vss bl[343] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_344 br[343] vdd vss bl[343] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_345 br[344] vdd vss bl[344] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_345 br[344] vdd vss bl[344] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_345 br[344] vdd vss bl[344] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_345 br[344] vdd vss bl[344] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_345 br[344] vdd vss bl[344] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_345 br[344] vdd vss bl[344] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_345 br[344] vdd vss bl[344] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_345 br[344] vdd vss bl[344] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_345 br[344] vdd vss bl[344] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_345 br[344] vdd vss bl[344] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_345 br[344] vdd vss bl[344] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_345 br[344] vdd vss bl[344] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_345 br[344] vdd vss bl[344] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_345 br[344] vdd vss bl[344] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_345 br[344] vdd vss bl[344] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_345 br[344] vdd vss bl[344] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_345 br[344] vdd vss bl[344] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_345 br[344] vdd vss bl[344] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_345 br[344] vdd vss bl[344] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_346 br[345] vdd vss bl[345] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_346 br[345] vdd vss bl[345] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_346 br[345] vdd vss bl[345] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_346 br[345] vdd vss bl[345] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_346 br[345] vdd vss bl[345] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_346 br[345] vdd vss bl[345] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_346 br[345] vdd vss bl[345] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_346 br[345] vdd vss bl[345] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_346 br[345] vdd vss bl[345] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_346 br[345] vdd vss bl[345] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_346 br[345] vdd vss bl[345] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_346 br[345] vdd vss bl[345] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_346 br[345] vdd vss bl[345] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_346 br[345] vdd vss bl[345] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_346 br[345] vdd vss bl[345] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_346 br[345] vdd vss bl[345] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_346 br[345] vdd vss bl[345] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_346 br[345] vdd vss bl[345] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_346 br[345] vdd vss bl[345] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_347 br[346] vdd vss bl[346] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_347 br[346] vdd vss bl[346] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_347 br[346] vdd vss bl[346] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_347 br[346] vdd vss bl[346] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_347 br[346] vdd vss bl[346] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_347 br[346] vdd vss bl[346] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_347 br[346] vdd vss bl[346] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_347 br[346] vdd vss bl[346] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_347 br[346] vdd vss bl[346] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_347 br[346] vdd vss bl[346] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_347 br[346] vdd vss bl[346] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_347 br[346] vdd vss bl[346] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_347 br[346] vdd vss bl[346] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_347 br[346] vdd vss bl[346] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_347 br[346] vdd vss bl[346] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_347 br[346] vdd vss bl[346] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_347 br[346] vdd vss bl[346] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_347 br[346] vdd vss bl[346] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_347 br[346] vdd vss bl[346] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_348 br[347] vdd vss bl[347] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_348 br[347] vdd vss bl[347] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_348 br[347] vdd vss bl[347] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_348 br[347] vdd vss bl[347] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_348 br[347] vdd vss bl[347] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_348 br[347] vdd vss bl[347] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_348 br[347] vdd vss bl[347] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_348 br[347] vdd vss bl[347] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_348 br[347] vdd vss bl[347] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_348 br[347] vdd vss bl[347] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_348 br[347] vdd vss bl[347] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_348 br[347] vdd vss bl[347] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_348 br[347] vdd vss bl[347] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_348 br[347] vdd vss bl[347] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_348 br[347] vdd vss bl[347] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_348 br[347] vdd vss bl[347] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_348 br[347] vdd vss bl[347] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_348 br[347] vdd vss bl[347] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_348 br[347] vdd vss bl[347] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_349 br[348] vdd vss bl[348] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_349 br[348] vdd vss bl[348] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_349 br[348] vdd vss bl[348] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_349 br[348] vdd vss bl[348] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_349 br[348] vdd vss bl[348] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_349 br[348] vdd vss bl[348] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_349 br[348] vdd vss bl[348] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_349 br[348] vdd vss bl[348] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_349 br[348] vdd vss bl[348] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_349 br[348] vdd vss bl[348] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_349 br[348] vdd vss bl[348] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_349 br[348] vdd vss bl[348] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_349 br[348] vdd vss bl[348] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_349 br[348] vdd vss bl[348] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_349 br[348] vdd vss bl[348] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_349 br[348] vdd vss bl[348] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_349 br[348] vdd vss bl[348] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_349 br[348] vdd vss bl[348] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_349 br[348] vdd vss bl[348] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_350 br[349] vdd vss bl[349] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_350 br[349] vdd vss bl[349] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_350 br[349] vdd vss bl[349] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_350 br[349] vdd vss bl[349] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_350 br[349] vdd vss bl[349] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_350 br[349] vdd vss bl[349] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_350 br[349] vdd vss bl[349] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_350 br[349] vdd vss bl[349] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_350 br[349] vdd vss bl[349] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_350 br[349] vdd vss bl[349] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_350 br[349] vdd vss bl[349] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_350 br[349] vdd vss bl[349] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_350 br[349] vdd vss bl[349] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_350 br[349] vdd vss bl[349] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_350 br[349] vdd vss bl[349] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_350 br[349] vdd vss bl[349] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_350 br[349] vdd vss bl[349] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_350 br[349] vdd vss bl[349] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_350 br[349] vdd vss bl[349] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_351 br[350] vdd vss bl[350] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_351 br[350] vdd vss bl[350] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_351 br[350] vdd vss bl[350] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_351 br[350] vdd vss bl[350] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_351 br[350] vdd vss bl[350] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_351 br[350] vdd vss bl[350] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_351 br[350] vdd vss bl[350] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_351 br[350] vdd vss bl[350] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_351 br[350] vdd vss bl[350] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_351 br[350] vdd vss bl[350] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_351 br[350] vdd vss bl[350] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_351 br[350] vdd vss bl[350] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_351 br[350] vdd vss bl[350] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_351 br[350] vdd vss bl[350] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_351 br[350] vdd vss bl[350] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_351 br[350] vdd vss bl[350] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_351 br[350] vdd vss bl[350] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_351 br[350] vdd vss bl[350] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_351 br[350] vdd vss bl[350] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_352 br[351] vdd vss bl[351] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_352 br[351] vdd vss bl[351] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_352 br[351] vdd vss bl[351] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_352 br[351] vdd vss bl[351] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_352 br[351] vdd vss bl[351] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_352 br[351] vdd vss bl[351] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_352 br[351] vdd vss bl[351] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_352 br[351] vdd vss bl[351] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_352 br[351] vdd vss bl[351] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_352 br[351] vdd vss bl[351] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_352 br[351] vdd vss bl[351] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_352 br[351] vdd vss bl[351] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_352 br[351] vdd vss bl[351] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_352 br[351] vdd vss bl[351] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_352 br[351] vdd vss bl[351] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_352 br[351] vdd vss bl[351] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_352 br[351] vdd vss bl[351] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_352 br[351] vdd vss bl[351] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_352 br[351] vdd vss bl[351] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_353 br[352] vdd vss bl[352] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_353 br[352] vdd vss bl[352] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_353 br[352] vdd vss bl[352] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_353 br[352] vdd vss bl[352] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_353 br[352] vdd vss bl[352] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_353 br[352] vdd vss bl[352] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_353 br[352] vdd vss bl[352] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_353 br[352] vdd vss bl[352] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_353 br[352] vdd vss bl[352] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_353 br[352] vdd vss bl[352] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_353 br[352] vdd vss bl[352] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_353 br[352] vdd vss bl[352] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_353 br[352] vdd vss bl[352] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_353 br[352] vdd vss bl[352] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_353 br[352] vdd vss bl[352] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_353 br[352] vdd vss bl[352] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_353 br[352] vdd vss bl[352] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_353 br[352] vdd vss bl[352] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_353 br[352] vdd vss bl[352] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_354 br[353] vdd vss bl[353] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_354 br[353] vdd vss bl[353] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_354 br[353] vdd vss bl[353] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_354 br[353] vdd vss bl[353] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_354 br[353] vdd vss bl[353] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_354 br[353] vdd vss bl[353] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_354 br[353] vdd vss bl[353] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_354 br[353] vdd vss bl[353] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_354 br[353] vdd vss bl[353] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_354 br[353] vdd vss bl[353] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_354 br[353] vdd vss bl[353] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_354 br[353] vdd vss bl[353] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_354 br[353] vdd vss bl[353] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_354 br[353] vdd vss bl[353] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_354 br[353] vdd vss bl[353] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_354 br[353] vdd vss bl[353] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_354 br[353] vdd vss bl[353] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_354 br[353] vdd vss bl[353] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_354 br[353] vdd vss bl[353] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_355 br[354] vdd vss bl[354] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_355 br[354] vdd vss bl[354] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_355 br[354] vdd vss bl[354] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_355 br[354] vdd vss bl[354] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_355 br[354] vdd vss bl[354] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_355 br[354] vdd vss bl[354] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_355 br[354] vdd vss bl[354] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_355 br[354] vdd vss bl[354] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_355 br[354] vdd vss bl[354] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_355 br[354] vdd vss bl[354] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_355 br[354] vdd vss bl[354] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_355 br[354] vdd vss bl[354] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_355 br[354] vdd vss bl[354] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_355 br[354] vdd vss bl[354] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_355 br[354] vdd vss bl[354] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_355 br[354] vdd vss bl[354] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_355 br[354] vdd vss bl[354] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_355 br[354] vdd vss bl[354] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_355 br[354] vdd vss bl[354] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_356 br[355] vdd vss bl[355] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_356 br[355] vdd vss bl[355] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_356 br[355] vdd vss bl[355] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_356 br[355] vdd vss bl[355] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_356 br[355] vdd vss bl[355] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_356 br[355] vdd vss bl[355] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_356 br[355] vdd vss bl[355] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_356 br[355] vdd vss bl[355] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_356 br[355] vdd vss bl[355] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_356 br[355] vdd vss bl[355] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_356 br[355] vdd vss bl[355] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_356 br[355] vdd vss bl[355] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_356 br[355] vdd vss bl[355] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_356 br[355] vdd vss bl[355] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_356 br[355] vdd vss bl[355] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_356 br[355] vdd vss bl[355] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_356 br[355] vdd vss bl[355] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_356 br[355] vdd vss bl[355] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_356 br[355] vdd vss bl[355] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_357 br[356] vdd vss bl[356] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_357 br[356] vdd vss bl[356] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_357 br[356] vdd vss bl[356] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_357 br[356] vdd vss bl[356] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_357 br[356] vdd vss bl[356] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_357 br[356] vdd vss bl[356] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_357 br[356] vdd vss bl[356] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_357 br[356] vdd vss bl[356] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_357 br[356] vdd vss bl[356] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_357 br[356] vdd vss bl[356] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_357 br[356] vdd vss bl[356] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_357 br[356] vdd vss bl[356] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_357 br[356] vdd vss bl[356] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_357 br[356] vdd vss bl[356] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_357 br[356] vdd vss bl[356] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_357 br[356] vdd vss bl[356] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_357 br[356] vdd vss bl[356] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_357 br[356] vdd vss bl[356] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_357 br[356] vdd vss bl[356] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_358 br[357] vdd vss bl[357] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_358 br[357] vdd vss bl[357] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_358 br[357] vdd vss bl[357] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_358 br[357] vdd vss bl[357] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_358 br[357] vdd vss bl[357] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_358 br[357] vdd vss bl[357] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_358 br[357] vdd vss bl[357] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_358 br[357] vdd vss bl[357] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_358 br[357] vdd vss bl[357] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_358 br[357] vdd vss bl[357] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_358 br[357] vdd vss bl[357] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_358 br[357] vdd vss bl[357] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_358 br[357] vdd vss bl[357] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_358 br[357] vdd vss bl[357] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_358 br[357] vdd vss bl[357] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_358 br[357] vdd vss bl[357] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_358 br[357] vdd vss bl[357] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_358 br[357] vdd vss bl[357] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_358 br[357] vdd vss bl[357] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_359 br[358] vdd vss bl[358] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_359 br[358] vdd vss bl[358] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_359 br[358] vdd vss bl[358] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_359 br[358] vdd vss bl[358] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_359 br[358] vdd vss bl[358] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_359 br[358] vdd vss bl[358] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_359 br[358] vdd vss bl[358] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_359 br[358] vdd vss bl[358] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_359 br[358] vdd vss bl[358] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_359 br[358] vdd vss bl[358] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_359 br[358] vdd vss bl[358] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_359 br[358] vdd vss bl[358] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_359 br[358] vdd vss bl[358] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_359 br[358] vdd vss bl[358] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_359 br[358] vdd vss bl[358] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_359 br[358] vdd vss bl[358] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_359 br[358] vdd vss bl[358] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_359 br[358] vdd vss bl[358] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_359 br[358] vdd vss bl[358] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_360 br[359] vdd vss bl[359] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_360 br[359] vdd vss bl[359] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_360 br[359] vdd vss bl[359] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_360 br[359] vdd vss bl[359] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_360 br[359] vdd vss bl[359] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_360 br[359] vdd vss bl[359] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_360 br[359] vdd vss bl[359] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_360 br[359] vdd vss bl[359] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_360 br[359] vdd vss bl[359] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_360 br[359] vdd vss bl[359] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_360 br[359] vdd vss bl[359] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_360 br[359] vdd vss bl[359] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_360 br[359] vdd vss bl[359] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_360 br[359] vdd vss bl[359] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_360 br[359] vdd vss bl[359] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_360 br[359] vdd vss bl[359] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_360 br[359] vdd vss bl[359] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_360 br[359] vdd vss bl[359] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_360 br[359] vdd vss bl[359] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_361 br[360] vdd vss bl[360] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_361 br[360] vdd vss bl[360] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_361 br[360] vdd vss bl[360] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_361 br[360] vdd vss bl[360] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_361 br[360] vdd vss bl[360] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_361 br[360] vdd vss bl[360] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_361 br[360] vdd vss bl[360] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_361 br[360] vdd vss bl[360] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_361 br[360] vdd vss bl[360] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_361 br[360] vdd vss bl[360] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_361 br[360] vdd vss bl[360] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_361 br[360] vdd vss bl[360] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_361 br[360] vdd vss bl[360] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_361 br[360] vdd vss bl[360] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_361 br[360] vdd vss bl[360] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_361 br[360] vdd vss bl[360] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_361 br[360] vdd vss bl[360] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_361 br[360] vdd vss bl[360] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_361 br[360] vdd vss bl[360] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_362 br[361] vdd vss bl[361] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_362 br[361] vdd vss bl[361] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_362 br[361] vdd vss bl[361] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_362 br[361] vdd vss bl[361] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_362 br[361] vdd vss bl[361] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_362 br[361] vdd vss bl[361] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_362 br[361] vdd vss bl[361] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_362 br[361] vdd vss bl[361] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_362 br[361] vdd vss bl[361] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_362 br[361] vdd vss bl[361] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_362 br[361] vdd vss bl[361] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_362 br[361] vdd vss bl[361] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_362 br[361] vdd vss bl[361] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_362 br[361] vdd vss bl[361] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_362 br[361] vdd vss bl[361] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_362 br[361] vdd vss bl[361] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_362 br[361] vdd vss bl[361] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_362 br[361] vdd vss bl[361] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_362 br[361] vdd vss bl[361] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_363 br[362] vdd vss bl[362] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_363 br[362] vdd vss bl[362] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_363 br[362] vdd vss bl[362] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_363 br[362] vdd vss bl[362] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_363 br[362] vdd vss bl[362] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_363 br[362] vdd vss bl[362] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_363 br[362] vdd vss bl[362] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_363 br[362] vdd vss bl[362] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_363 br[362] vdd vss bl[362] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_363 br[362] vdd vss bl[362] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_363 br[362] vdd vss bl[362] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_363 br[362] vdd vss bl[362] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_363 br[362] vdd vss bl[362] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_363 br[362] vdd vss bl[362] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_363 br[362] vdd vss bl[362] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_363 br[362] vdd vss bl[362] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_363 br[362] vdd vss bl[362] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_363 br[362] vdd vss bl[362] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_363 br[362] vdd vss bl[362] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_364 br[363] vdd vss bl[363] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_364 br[363] vdd vss bl[363] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_364 br[363] vdd vss bl[363] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_364 br[363] vdd vss bl[363] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_364 br[363] vdd vss bl[363] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_364 br[363] vdd vss bl[363] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_364 br[363] vdd vss bl[363] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_364 br[363] vdd vss bl[363] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_364 br[363] vdd vss bl[363] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_364 br[363] vdd vss bl[363] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_364 br[363] vdd vss bl[363] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_364 br[363] vdd vss bl[363] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_364 br[363] vdd vss bl[363] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_364 br[363] vdd vss bl[363] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_364 br[363] vdd vss bl[363] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_364 br[363] vdd vss bl[363] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_364 br[363] vdd vss bl[363] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_364 br[363] vdd vss bl[363] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_364 br[363] vdd vss bl[363] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_365 br[364] vdd vss bl[364] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_365 br[364] vdd vss bl[364] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_365 br[364] vdd vss bl[364] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_365 br[364] vdd vss bl[364] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_365 br[364] vdd vss bl[364] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_365 br[364] vdd vss bl[364] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_365 br[364] vdd vss bl[364] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_365 br[364] vdd vss bl[364] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_365 br[364] vdd vss bl[364] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_365 br[364] vdd vss bl[364] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_365 br[364] vdd vss bl[364] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_365 br[364] vdd vss bl[364] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_365 br[364] vdd vss bl[364] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_365 br[364] vdd vss bl[364] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_365 br[364] vdd vss bl[364] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_365 br[364] vdd vss bl[364] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_365 br[364] vdd vss bl[364] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_365 br[364] vdd vss bl[364] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_365 br[364] vdd vss bl[364] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_366 br[365] vdd vss bl[365] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_366 br[365] vdd vss bl[365] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_366 br[365] vdd vss bl[365] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_366 br[365] vdd vss bl[365] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_366 br[365] vdd vss bl[365] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_366 br[365] vdd vss bl[365] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_366 br[365] vdd vss bl[365] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_366 br[365] vdd vss bl[365] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_366 br[365] vdd vss bl[365] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_366 br[365] vdd vss bl[365] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_366 br[365] vdd vss bl[365] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_366 br[365] vdd vss bl[365] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_366 br[365] vdd vss bl[365] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_366 br[365] vdd vss bl[365] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_366 br[365] vdd vss bl[365] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_366 br[365] vdd vss bl[365] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_366 br[365] vdd vss bl[365] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_366 br[365] vdd vss bl[365] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_366 br[365] vdd vss bl[365] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_367 br[366] vdd vss bl[366] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_367 br[366] vdd vss bl[366] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_367 br[366] vdd vss bl[366] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_367 br[366] vdd vss bl[366] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_367 br[366] vdd vss bl[366] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_367 br[366] vdd vss bl[366] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_367 br[366] vdd vss bl[366] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_367 br[366] vdd vss bl[366] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_367 br[366] vdd vss bl[366] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_367 br[366] vdd vss bl[366] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_367 br[366] vdd vss bl[366] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_367 br[366] vdd vss bl[366] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_367 br[366] vdd vss bl[366] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_367 br[366] vdd vss bl[366] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_367 br[366] vdd vss bl[366] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_367 br[366] vdd vss bl[366] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_367 br[366] vdd vss bl[366] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_367 br[366] vdd vss bl[366] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_367 br[366] vdd vss bl[366] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_368 br[367] vdd vss bl[367] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_368 br[367] vdd vss bl[367] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_368 br[367] vdd vss bl[367] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_368 br[367] vdd vss bl[367] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_368 br[367] vdd vss bl[367] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_368 br[367] vdd vss bl[367] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_368 br[367] vdd vss bl[367] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_368 br[367] vdd vss bl[367] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_368 br[367] vdd vss bl[367] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_368 br[367] vdd vss bl[367] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_368 br[367] vdd vss bl[367] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_368 br[367] vdd vss bl[367] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_368 br[367] vdd vss bl[367] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_368 br[367] vdd vss bl[367] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_368 br[367] vdd vss bl[367] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_368 br[367] vdd vss bl[367] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_368 br[367] vdd vss bl[367] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_368 br[367] vdd vss bl[367] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_368 br[367] vdd vss bl[367] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_369 br[368] vdd vss bl[368] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_369 br[368] vdd vss bl[368] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_369 br[368] vdd vss bl[368] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_369 br[368] vdd vss bl[368] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_369 br[368] vdd vss bl[368] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_369 br[368] vdd vss bl[368] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_369 br[368] vdd vss bl[368] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_369 br[368] vdd vss bl[368] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_369 br[368] vdd vss bl[368] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_369 br[368] vdd vss bl[368] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_369 br[368] vdd vss bl[368] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_369 br[368] vdd vss bl[368] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_369 br[368] vdd vss bl[368] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_369 br[368] vdd vss bl[368] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_369 br[368] vdd vss bl[368] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_369 br[368] vdd vss bl[368] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_369 br[368] vdd vss bl[368] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_369 br[368] vdd vss bl[368] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_369 br[368] vdd vss bl[368] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_370 br[369] vdd vss bl[369] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_370 br[369] vdd vss bl[369] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_370 br[369] vdd vss bl[369] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_370 br[369] vdd vss bl[369] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_370 br[369] vdd vss bl[369] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_370 br[369] vdd vss bl[369] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_370 br[369] vdd vss bl[369] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_370 br[369] vdd vss bl[369] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_370 br[369] vdd vss bl[369] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_370 br[369] vdd vss bl[369] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_370 br[369] vdd vss bl[369] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_370 br[369] vdd vss bl[369] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_370 br[369] vdd vss bl[369] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_370 br[369] vdd vss bl[369] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_370 br[369] vdd vss bl[369] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_370 br[369] vdd vss bl[369] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_370 br[369] vdd vss bl[369] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_370 br[369] vdd vss bl[369] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_370 br[369] vdd vss bl[369] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_371 br[370] vdd vss bl[370] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_371 br[370] vdd vss bl[370] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_371 br[370] vdd vss bl[370] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_371 br[370] vdd vss bl[370] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_371 br[370] vdd vss bl[370] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_371 br[370] vdd vss bl[370] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_371 br[370] vdd vss bl[370] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_371 br[370] vdd vss bl[370] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_371 br[370] vdd vss bl[370] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_371 br[370] vdd vss bl[370] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_371 br[370] vdd vss bl[370] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_371 br[370] vdd vss bl[370] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_371 br[370] vdd vss bl[370] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_371 br[370] vdd vss bl[370] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_371 br[370] vdd vss bl[370] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_371 br[370] vdd vss bl[370] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_371 br[370] vdd vss bl[370] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_371 br[370] vdd vss bl[370] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_371 br[370] vdd vss bl[370] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_372 br[371] vdd vss bl[371] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_372 br[371] vdd vss bl[371] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_372 br[371] vdd vss bl[371] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_372 br[371] vdd vss bl[371] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_372 br[371] vdd vss bl[371] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_372 br[371] vdd vss bl[371] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_372 br[371] vdd vss bl[371] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_372 br[371] vdd vss bl[371] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_372 br[371] vdd vss bl[371] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_372 br[371] vdd vss bl[371] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_372 br[371] vdd vss bl[371] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_372 br[371] vdd vss bl[371] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_372 br[371] vdd vss bl[371] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_372 br[371] vdd vss bl[371] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_372 br[371] vdd vss bl[371] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_372 br[371] vdd vss bl[371] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_372 br[371] vdd vss bl[371] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_372 br[371] vdd vss bl[371] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_372 br[371] vdd vss bl[371] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_373 br[372] vdd vss bl[372] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_373 br[372] vdd vss bl[372] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_373 br[372] vdd vss bl[372] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_373 br[372] vdd vss bl[372] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_373 br[372] vdd vss bl[372] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_373 br[372] vdd vss bl[372] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_373 br[372] vdd vss bl[372] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_373 br[372] vdd vss bl[372] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_373 br[372] vdd vss bl[372] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_373 br[372] vdd vss bl[372] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_373 br[372] vdd vss bl[372] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_373 br[372] vdd vss bl[372] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_373 br[372] vdd vss bl[372] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_373 br[372] vdd vss bl[372] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_373 br[372] vdd vss bl[372] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_373 br[372] vdd vss bl[372] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_373 br[372] vdd vss bl[372] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_373 br[372] vdd vss bl[372] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_373 br[372] vdd vss bl[372] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_374 br[373] vdd vss bl[373] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_374 br[373] vdd vss bl[373] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_374 br[373] vdd vss bl[373] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_374 br[373] vdd vss bl[373] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_374 br[373] vdd vss bl[373] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_374 br[373] vdd vss bl[373] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_374 br[373] vdd vss bl[373] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_374 br[373] vdd vss bl[373] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_374 br[373] vdd vss bl[373] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_374 br[373] vdd vss bl[373] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_374 br[373] vdd vss bl[373] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_374 br[373] vdd vss bl[373] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_374 br[373] vdd vss bl[373] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_374 br[373] vdd vss bl[373] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_374 br[373] vdd vss bl[373] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_374 br[373] vdd vss bl[373] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_374 br[373] vdd vss bl[373] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_374 br[373] vdd vss bl[373] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_374 br[373] vdd vss bl[373] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_375 br[374] vdd vss bl[374] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_375 br[374] vdd vss bl[374] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_375 br[374] vdd vss bl[374] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_375 br[374] vdd vss bl[374] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_375 br[374] vdd vss bl[374] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_375 br[374] vdd vss bl[374] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_375 br[374] vdd vss bl[374] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_375 br[374] vdd vss bl[374] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_375 br[374] vdd vss bl[374] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_375 br[374] vdd vss bl[374] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_375 br[374] vdd vss bl[374] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_375 br[374] vdd vss bl[374] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_375 br[374] vdd vss bl[374] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_375 br[374] vdd vss bl[374] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_375 br[374] vdd vss bl[374] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_375 br[374] vdd vss bl[374] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_375 br[374] vdd vss bl[374] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_375 br[374] vdd vss bl[374] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_375 br[374] vdd vss bl[374] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_376 br[375] vdd vss bl[375] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_376 br[375] vdd vss bl[375] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_376 br[375] vdd vss bl[375] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_376 br[375] vdd vss bl[375] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_376 br[375] vdd vss bl[375] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_376 br[375] vdd vss bl[375] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_376 br[375] vdd vss bl[375] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_376 br[375] vdd vss bl[375] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_376 br[375] vdd vss bl[375] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_376 br[375] vdd vss bl[375] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_376 br[375] vdd vss bl[375] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_376 br[375] vdd vss bl[375] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_376 br[375] vdd vss bl[375] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_376 br[375] vdd vss bl[375] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_376 br[375] vdd vss bl[375] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_376 br[375] vdd vss bl[375] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_376 br[375] vdd vss bl[375] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_376 br[375] vdd vss bl[375] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_376 br[375] vdd vss bl[375] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_377 br[376] vdd vss bl[376] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_377 br[376] vdd vss bl[376] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_377 br[376] vdd vss bl[376] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_377 br[376] vdd vss bl[376] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_377 br[376] vdd vss bl[376] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_377 br[376] vdd vss bl[376] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_377 br[376] vdd vss bl[376] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_377 br[376] vdd vss bl[376] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_377 br[376] vdd vss bl[376] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_377 br[376] vdd vss bl[376] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_377 br[376] vdd vss bl[376] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_377 br[376] vdd vss bl[376] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_377 br[376] vdd vss bl[376] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_377 br[376] vdd vss bl[376] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_377 br[376] vdd vss bl[376] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_377 br[376] vdd vss bl[376] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_377 br[376] vdd vss bl[376] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_377 br[376] vdd vss bl[376] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_377 br[376] vdd vss bl[376] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_378 br[377] vdd vss bl[377] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_378 br[377] vdd vss bl[377] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_378 br[377] vdd vss bl[377] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_378 br[377] vdd vss bl[377] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_378 br[377] vdd vss bl[377] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_378 br[377] vdd vss bl[377] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_378 br[377] vdd vss bl[377] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_378 br[377] vdd vss bl[377] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_378 br[377] vdd vss bl[377] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_378 br[377] vdd vss bl[377] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_378 br[377] vdd vss bl[377] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_378 br[377] vdd vss bl[377] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_378 br[377] vdd vss bl[377] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_378 br[377] vdd vss bl[377] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_378 br[377] vdd vss bl[377] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_378 br[377] vdd vss bl[377] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_378 br[377] vdd vss bl[377] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_378 br[377] vdd vss bl[377] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_378 br[377] vdd vss bl[377] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_379 br[378] vdd vss bl[378] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_379 br[378] vdd vss bl[378] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_379 br[378] vdd vss bl[378] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_379 br[378] vdd vss bl[378] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_379 br[378] vdd vss bl[378] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_379 br[378] vdd vss bl[378] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_379 br[378] vdd vss bl[378] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_379 br[378] vdd vss bl[378] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_379 br[378] vdd vss bl[378] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_379 br[378] vdd vss bl[378] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_379 br[378] vdd vss bl[378] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_379 br[378] vdd vss bl[378] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_379 br[378] vdd vss bl[378] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_379 br[378] vdd vss bl[378] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_379 br[378] vdd vss bl[378] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_379 br[378] vdd vss bl[378] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_379 br[378] vdd vss bl[378] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_379 br[378] vdd vss bl[378] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_379 br[378] vdd vss bl[378] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_380 br[379] vdd vss bl[379] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_380 br[379] vdd vss bl[379] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_380 br[379] vdd vss bl[379] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_380 br[379] vdd vss bl[379] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_380 br[379] vdd vss bl[379] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_380 br[379] vdd vss bl[379] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_380 br[379] vdd vss bl[379] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_380 br[379] vdd vss bl[379] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_380 br[379] vdd vss bl[379] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_380 br[379] vdd vss bl[379] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_380 br[379] vdd vss bl[379] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_380 br[379] vdd vss bl[379] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_380 br[379] vdd vss bl[379] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_380 br[379] vdd vss bl[379] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_380 br[379] vdd vss bl[379] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_380 br[379] vdd vss bl[379] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_380 br[379] vdd vss bl[379] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_380 br[379] vdd vss bl[379] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_380 br[379] vdd vss bl[379] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_381 br[380] vdd vss bl[380] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_381 br[380] vdd vss bl[380] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_381 br[380] vdd vss bl[380] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_381 br[380] vdd vss bl[380] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_381 br[380] vdd vss bl[380] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_381 br[380] vdd vss bl[380] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_381 br[380] vdd vss bl[380] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_381 br[380] vdd vss bl[380] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_381 br[380] vdd vss bl[380] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_381 br[380] vdd vss bl[380] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_381 br[380] vdd vss bl[380] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_381 br[380] vdd vss bl[380] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_381 br[380] vdd vss bl[380] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_381 br[380] vdd vss bl[380] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_381 br[380] vdd vss bl[380] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_381 br[380] vdd vss bl[380] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_381 br[380] vdd vss bl[380] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_381 br[380] vdd vss bl[380] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_381 br[380] vdd vss bl[380] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_382 br[381] vdd vss bl[381] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_382 br[381] vdd vss bl[381] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_382 br[381] vdd vss bl[381] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_382 br[381] vdd vss bl[381] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_382 br[381] vdd vss bl[381] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_382 br[381] vdd vss bl[381] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_382 br[381] vdd vss bl[381] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_382 br[381] vdd vss bl[381] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_382 br[381] vdd vss bl[381] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_382 br[381] vdd vss bl[381] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_382 br[381] vdd vss bl[381] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_382 br[381] vdd vss bl[381] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_382 br[381] vdd vss bl[381] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_382 br[381] vdd vss bl[381] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_382 br[381] vdd vss bl[381] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_382 br[381] vdd vss bl[381] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_382 br[381] vdd vss bl[381] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_382 br[381] vdd vss bl[381] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_382 br[381] vdd vss bl[381] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_383 br[382] vdd vss bl[382] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_383 br[382] vdd vss bl[382] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_383 br[382] vdd vss bl[382] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_383 br[382] vdd vss bl[382] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_383 br[382] vdd vss bl[382] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_383 br[382] vdd vss bl[382] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_383 br[382] vdd vss bl[382] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_383 br[382] vdd vss bl[382] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_383 br[382] vdd vss bl[382] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_383 br[382] vdd vss bl[382] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_383 br[382] vdd vss bl[382] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_383 br[382] vdd vss bl[382] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_383 br[382] vdd vss bl[382] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_383 br[382] vdd vss bl[382] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_383 br[382] vdd vss bl[382] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_383 br[382] vdd vss bl[382] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_383 br[382] vdd vss bl[382] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_383 br[382] vdd vss bl[382] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_383 br[382] vdd vss bl[382] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_384 br[383] vdd vss bl[383] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_384 br[383] vdd vss bl[383] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_384 br[383] vdd vss bl[383] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_384 br[383] vdd vss bl[383] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_384 br[383] vdd vss bl[383] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_384 br[383] vdd vss bl[383] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_384 br[383] vdd vss bl[383] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_384 br[383] vdd vss bl[383] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_384 br[383] vdd vss bl[383] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_384 br[383] vdd vss bl[383] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_384 br[383] vdd vss bl[383] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_384 br[383] vdd vss bl[383] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_384 br[383] vdd vss bl[383] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_384 br[383] vdd vss bl[383] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_384 br[383] vdd vss bl[383] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_384 br[383] vdd vss bl[383] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_384 br[383] vdd vss bl[383] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_384 br[383] vdd vss bl[383] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_384 br[383] vdd vss bl[383] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_385 br[384] vdd vss bl[384] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_385 br[384] vdd vss bl[384] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_385 br[384] vdd vss bl[384] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_385 br[384] vdd vss bl[384] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_385 br[384] vdd vss bl[384] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_385 br[384] vdd vss bl[384] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_385 br[384] vdd vss bl[384] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_385 br[384] vdd vss bl[384] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_385 br[384] vdd vss bl[384] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_385 br[384] vdd vss bl[384] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_385 br[384] vdd vss bl[384] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_385 br[384] vdd vss bl[384] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_385 br[384] vdd vss bl[384] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_385 br[384] vdd vss bl[384] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_385 br[384] vdd vss bl[384] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_385 br[384] vdd vss bl[384] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_385 br[384] vdd vss bl[384] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_385 br[384] vdd vss bl[384] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_385 br[384] vdd vss bl[384] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_386 br[385] vdd vss bl[385] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_386 br[385] vdd vss bl[385] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_386 br[385] vdd vss bl[385] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_386 br[385] vdd vss bl[385] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_386 br[385] vdd vss bl[385] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_386 br[385] vdd vss bl[385] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_386 br[385] vdd vss bl[385] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_386 br[385] vdd vss bl[385] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_386 br[385] vdd vss bl[385] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_386 br[385] vdd vss bl[385] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_386 br[385] vdd vss bl[385] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_386 br[385] vdd vss bl[385] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_386 br[385] vdd vss bl[385] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_386 br[385] vdd vss bl[385] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_386 br[385] vdd vss bl[385] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_386 br[385] vdd vss bl[385] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_386 br[385] vdd vss bl[385] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_386 br[385] vdd vss bl[385] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_386 br[385] vdd vss bl[385] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_387 br[386] vdd vss bl[386] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_387 br[386] vdd vss bl[386] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_387 br[386] vdd vss bl[386] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_387 br[386] vdd vss bl[386] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_387 br[386] vdd vss bl[386] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_387 br[386] vdd vss bl[386] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_387 br[386] vdd vss bl[386] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_387 br[386] vdd vss bl[386] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_387 br[386] vdd vss bl[386] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_387 br[386] vdd vss bl[386] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_387 br[386] vdd vss bl[386] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_387 br[386] vdd vss bl[386] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_387 br[386] vdd vss bl[386] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_387 br[386] vdd vss bl[386] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_387 br[386] vdd vss bl[386] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_387 br[386] vdd vss bl[386] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_387 br[386] vdd vss bl[386] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_387 br[386] vdd vss bl[386] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_387 br[386] vdd vss bl[386] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_388 br[387] vdd vss bl[387] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_388 br[387] vdd vss bl[387] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_388 br[387] vdd vss bl[387] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_388 br[387] vdd vss bl[387] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_388 br[387] vdd vss bl[387] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_388 br[387] vdd vss bl[387] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_388 br[387] vdd vss bl[387] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_388 br[387] vdd vss bl[387] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_388 br[387] vdd vss bl[387] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_388 br[387] vdd vss bl[387] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_388 br[387] vdd vss bl[387] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_388 br[387] vdd vss bl[387] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_388 br[387] vdd vss bl[387] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_388 br[387] vdd vss bl[387] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_388 br[387] vdd vss bl[387] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_388 br[387] vdd vss bl[387] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_388 br[387] vdd vss bl[387] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_388 br[387] vdd vss bl[387] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_388 br[387] vdd vss bl[387] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_389 br[388] vdd vss bl[388] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_389 br[388] vdd vss bl[388] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_389 br[388] vdd vss bl[388] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_389 br[388] vdd vss bl[388] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_389 br[388] vdd vss bl[388] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_389 br[388] vdd vss bl[388] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_389 br[388] vdd vss bl[388] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_389 br[388] vdd vss bl[388] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_389 br[388] vdd vss bl[388] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_389 br[388] vdd vss bl[388] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_389 br[388] vdd vss bl[388] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_389 br[388] vdd vss bl[388] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_389 br[388] vdd vss bl[388] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_389 br[388] vdd vss bl[388] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_389 br[388] vdd vss bl[388] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_389 br[388] vdd vss bl[388] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_389 br[388] vdd vss bl[388] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_389 br[388] vdd vss bl[388] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_389 br[388] vdd vss bl[388] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_390 br[389] vdd vss bl[389] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_390 br[389] vdd vss bl[389] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_390 br[389] vdd vss bl[389] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_390 br[389] vdd vss bl[389] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_390 br[389] vdd vss bl[389] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_390 br[389] vdd vss bl[389] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_390 br[389] vdd vss bl[389] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_390 br[389] vdd vss bl[389] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_390 br[389] vdd vss bl[389] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_390 br[389] vdd vss bl[389] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_390 br[389] vdd vss bl[389] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_390 br[389] vdd vss bl[389] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_390 br[389] vdd vss bl[389] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_390 br[389] vdd vss bl[389] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_390 br[389] vdd vss bl[389] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_390 br[389] vdd vss bl[389] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_390 br[389] vdd vss bl[389] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_390 br[389] vdd vss bl[389] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_390 br[389] vdd vss bl[389] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_391 br[390] vdd vss bl[390] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_391 br[390] vdd vss bl[390] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_391 br[390] vdd vss bl[390] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_391 br[390] vdd vss bl[390] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_391 br[390] vdd vss bl[390] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_391 br[390] vdd vss bl[390] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_391 br[390] vdd vss bl[390] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_391 br[390] vdd vss bl[390] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_391 br[390] vdd vss bl[390] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_391 br[390] vdd vss bl[390] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_391 br[390] vdd vss bl[390] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_391 br[390] vdd vss bl[390] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_391 br[390] vdd vss bl[390] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_391 br[390] vdd vss bl[390] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_391 br[390] vdd vss bl[390] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_391 br[390] vdd vss bl[390] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_391 br[390] vdd vss bl[390] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_391 br[390] vdd vss bl[390] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_391 br[390] vdd vss bl[390] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_392 br[391] vdd vss bl[391] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_392 br[391] vdd vss bl[391] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_392 br[391] vdd vss bl[391] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_392 br[391] vdd vss bl[391] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_392 br[391] vdd vss bl[391] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_392 br[391] vdd vss bl[391] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_392 br[391] vdd vss bl[391] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_392 br[391] vdd vss bl[391] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_392 br[391] vdd vss bl[391] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_392 br[391] vdd vss bl[391] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_392 br[391] vdd vss bl[391] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_392 br[391] vdd vss bl[391] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_392 br[391] vdd vss bl[391] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_392 br[391] vdd vss bl[391] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_392 br[391] vdd vss bl[391] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_392 br[391] vdd vss bl[391] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_392 br[391] vdd vss bl[391] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_392 br[391] vdd vss bl[391] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_392 br[391] vdd vss bl[391] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_393 br[392] vdd vss bl[392] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_393 br[392] vdd vss bl[392] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_393 br[392] vdd vss bl[392] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_393 br[392] vdd vss bl[392] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_393 br[392] vdd vss bl[392] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_393 br[392] vdd vss bl[392] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_393 br[392] vdd vss bl[392] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_393 br[392] vdd vss bl[392] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_393 br[392] vdd vss bl[392] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_393 br[392] vdd vss bl[392] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_393 br[392] vdd vss bl[392] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_393 br[392] vdd vss bl[392] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_393 br[392] vdd vss bl[392] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_393 br[392] vdd vss bl[392] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_393 br[392] vdd vss bl[392] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_393 br[392] vdd vss bl[392] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_393 br[392] vdd vss bl[392] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_393 br[392] vdd vss bl[392] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_393 br[392] vdd vss bl[392] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_394 br[393] vdd vss bl[393] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_394 br[393] vdd vss bl[393] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_394 br[393] vdd vss bl[393] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_394 br[393] vdd vss bl[393] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_394 br[393] vdd vss bl[393] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_394 br[393] vdd vss bl[393] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_394 br[393] vdd vss bl[393] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_394 br[393] vdd vss bl[393] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_394 br[393] vdd vss bl[393] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_394 br[393] vdd vss bl[393] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_394 br[393] vdd vss bl[393] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_394 br[393] vdd vss bl[393] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_394 br[393] vdd vss bl[393] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_394 br[393] vdd vss bl[393] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_394 br[393] vdd vss bl[393] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_394 br[393] vdd vss bl[393] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_394 br[393] vdd vss bl[393] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_394 br[393] vdd vss bl[393] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_394 br[393] vdd vss bl[393] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_395 br[394] vdd vss bl[394] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_395 br[394] vdd vss bl[394] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_395 br[394] vdd vss bl[394] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_395 br[394] vdd vss bl[394] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_395 br[394] vdd vss bl[394] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_395 br[394] vdd vss bl[394] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_395 br[394] vdd vss bl[394] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_395 br[394] vdd vss bl[394] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_395 br[394] vdd vss bl[394] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_395 br[394] vdd vss bl[394] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_395 br[394] vdd vss bl[394] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_395 br[394] vdd vss bl[394] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_395 br[394] vdd vss bl[394] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_395 br[394] vdd vss bl[394] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_395 br[394] vdd vss bl[394] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_395 br[394] vdd vss bl[394] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_395 br[394] vdd vss bl[394] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_395 br[394] vdd vss bl[394] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_395 br[394] vdd vss bl[394] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_396 br[395] vdd vss bl[395] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_396 br[395] vdd vss bl[395] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_396 br[395] vdd vss bl[395] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_396 br[395] vdd vss bl[395] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_396 br[395] vdd vss bl[395] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_396 br[395] vdd vss bl[395] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_396 br[395] vdd vss bl[395] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_396 br[395] vdd vss bl[395] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_396 br[395] vdd vss bl[395] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_396 br[395] vdd vss bl[395] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_396 br[395] vdd vss bl[395] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_396 br[395] vdd vss bl[395] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_396 br[395] vdd vss bl[395] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_396 br[395] vdd vss bl[395] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_396 br[395] vdd vss bl[395] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_396 br[395] vdd vss bl[395] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_396 br[395] vdd vss bl[395] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_396 br[395] vdd vss bl[395] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_396 br[395] vdd vss bl[395] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_397 br[396] vdd vss bl[396] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_397 br[396] vdd vss bl[396] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_397 br[396] vdd vss bl[396] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_397 br[396] vdd vss bl[396] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_397 br[396] vdd vss bl[396] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_397 br[396] vdd vss bl[396] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_397 br[396] vdd vss bl[396] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_397 br[396] vdd vss bl[396] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_397 br[396] vdd vss bl[396] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_397 br[396] vdd vss bl[396] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_397 br[396] vdd vss bl[396] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_397 br[396] vdd vss bl[396] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_397 br[396] vdd vss bl[396] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_397 br[396] vdd vss bl[396] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_397 br[396] vdd vss bl[396] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_397 br[396] vdd vss bl[396] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_397 br[396] vdd vss bl[396] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_397 br[396] vdd vss bl[396] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_397 br[396] vdd vss bl[396] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_398 br[397] vdd vss bl[397] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_398 br[397] vdd vss bl[397] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_398 br[397] vdd vss bl[397] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_398 br[397] vdd vss bl[397] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_398 br[397] vdd vss bl[397] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_398 br[397] vdd vss bl[397] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_398 br[397] vdd vss bl[397] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_398 br[397] vdd vss bl[397] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_398 br[397] vdd vss bl[397] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_398 br[397] vdd vss bl[397] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_398 br[397] vdd vss bl[397] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_398 br[397] vdd vss bl[397] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_398 br[397] vdd vss bl[397] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_398 br[397] vdd vss bl[397] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_398 br[397] vdd vss bl[397] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_398 br[397] vdd vss bl[397] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_398 br[397] vdd vss bl[397] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_398 br[397] vdd vss bl[397] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_398 br[397] vdd vss bl[397] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_399 br[398] vdd vss bl[398] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_399 br[398] vdd vss bl[398] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_399 br[398] vdd vss bl[398] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_399 br[398] vdd vss bl[398] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_399 br[398] vdd vss bl[398] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_399 br[398] vdd vss bl[398] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_399 br[398] vdd vss bl[398] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_399 br[398] vdd vss bl[398] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_399 br[398] vdd vss bl[398] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_399 br[398] vdd vss bl[398] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_399 br[398] vdd vss bl[398] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_399 br[398] vdd vss bl[398] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_399 br[398] vdd vss bl[398] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_399 br[398] vdd vss bl[398] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_399 br[398] vdd vss bl[398] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_399 br[398] vdd vss bl[398] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_399 br[398] vdd vss bl[398] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_399 br[398] vdd vss bl[398] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_399 br[398] vdd vss bl[398] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_400 br[399] vdd vss bl[399] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_400 br[399] vdd vss bl[399] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_400 br[399] vdd vss bl[399] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_400 br[399] vdd vss bl[399] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_400 br[399] vdd vss bl[399] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_400 br[399] vdd vss bl[399] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_400 br[399] vdd vss bl[399] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_400 br[399] vdd vss bl[399] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_400 br[399] vdd vss bl[399] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_400 br[399] vdd vss bl[399] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_400 br[399] vdd vss bl[399] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_400 br[399] vdd vss bl[399] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_400 br[399] vdd vss bl[399] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_400 br[399] vdd vss bl[399] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_400 br[399] vdd vss bl[399] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_400 br[399] vdd vss bl[399] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_400 br[399] vdd vss bl[399] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_400 br[399] vdd vss bl[399] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_400 br[399] vdd vss bl[399] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_401 br[400] vdd vss bl[400] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_401 br[400] vdd vss bl[400] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_401 br[400] vdd vss bl[400] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_401 br[400] vdd vss bl[400] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_401 br[400] vdd vss bl[400] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_401 br[400] vdd vss bl[400] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_401 br[400] vdd vss bl[400] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_401 br[400] vdd vss bl[400] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_401 br[400] vdd vss bl[400] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_401 br[400] vdd vss bl[400] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_401 br[400] vdd vss bl[400] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_401 br[400] vdd vss bl[400] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_401 br[400] vdd vss bl[400] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_401 br[400] vdd vss bl[400] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_401 br[400] vdd vss bl[400] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_401 br[400] vdd vss bl[400] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_401 br[400] vdd vss bl[400] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_401 br[400] vdd vss bl[400] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_401 br[400] vdd vss bl[400] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_402 br[401] vdd vss bl[401] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_402 br[401] vdd vss bl[401] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_402 br[401] vdd vss bl[401] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_402 br[401] vdd vss bl[401] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_402 br[401] vdd vss bl[401] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_402 br[401] vdd vss bl[401] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_402 br[401] vdd vss bl[401] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_402 br[401] vdd vss bl[401] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_402 br[401] vdd vss bl[401] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_402 br[401] vdd vss bl[401] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_402 br[401] vdd vss bl[401] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_402 br[401] vdd vss bl[401] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_402 br[401] vdd vss bl[401] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_402 br[401] vdd vss bl[401] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_402 br[401] vdd vss bl[401] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_402 br[401] vdd vss bl[401] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_402 br[401] vdd vss bl[401] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_402 br[401] vdd vss bl[401] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_402 br[401] vdd vss bl[401] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_403 br[402] vdd vss bl[402] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_403 br[402] vdd vss bl[402] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_403 br[402] vdd vss bl[402] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_403 br[402] vdd vss bl[402] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_403 br[402] vdd vss bl[402] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_403 br[402] vdd vss bl[402] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_403 br[402] vdd vss bl[402] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_403 br[402] vdd vss bl[402] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_403 br[402] vdd vss bl[402] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_403 br[402] vdd vss bl[402] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_403 br[402] vdd vss bl[402] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_403 br[402] vdd vss bl[402] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_403 br[402] vdd vss bl[402] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_403 br[402] vdd vss bl[402] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_403 br[402] vdd vss bl[402] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_403 br[402] vdd vss bl[402] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_403 br[402] vdd vss bl[402] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_403 br[402] vdd vss bl[402] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_403 br[402] vdd vss bl[402] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_404 br[403] vdd vss bl[403] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_404 br[403] vdd vss bl[403] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_404 br[403] vdd vss bl[403] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_404 br[403] vdd vss bl[403] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_404 br[403] vdd vss bl[403] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_404 br[403] vdd vss bl[403] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_404 br[403] vdd vss bl[403] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_404 br[403] vdd vss bl[403] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_404 br[403] vdd vss bl[403] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_404 br[403] vdd vss bl[403] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_404 br[403] vdd vss bl[403] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_404 br[403] vdd vss bl[403] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_404 br[403] vdd vss bl[403] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_404 br[403] vdd vss bl[403] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_404 br[403] vdd vss bl[403] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_404 br[403] vdd vss bl[403] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_404 br[403] vdd vss bl[403] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_404 br[403] vdd vss bl[403] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_404 br[403] vdd vss bl[403] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_405 br[404] vdd vss bl[404] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_405 br[404] vdd vss bl[404] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_405 br[404] vdd vss bl[404] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_405 br[404] vdd vss bl[404] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_405 br[404] vdd vss bl[404] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_405 br[404] vdd vss bl[404] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_405 br[404] vdd vss bl[404] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_405 br[404] vdd vss bl[404] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_405 br[404] vdd vss bl[404] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_405 br[404] vdd vss bl[404] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_405 br[404] vdd vss bl[404] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_405 br[404] vdd vss bl[404] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_405 br[404] vdd vss bl[404] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_405 br[404] vdd vss bl[404] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_405 br[404] vdd vss bl[404] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_405 br[404] vdd vss bl[404] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_405 br[404] vdd vss bl[404] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_405 br[404] vdd vss bl[404] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_405 br[404] vdd vss bl[404] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_406 br[405] vdd vss bl[405] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_406 br[405] vdd vss bl[405] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_406 br[405] vdd vss bl[405] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_406 br[405] vdd vss bl[405] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_406 br[405] vdd vss bl[405] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_406 br[405] vdd vss bl[405] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_406 br[405] vdd vss bl[405] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_406 br[405] vdd vss bl[405] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_406 br[405] vdd vss bl[405] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_406 br[405] vdd vss bl[405] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_406 br[405] vdd vss bl[405] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_406 br[405] vdd vss bl[405] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_406 br[405] vdd vss bl[405] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_406 br[405] vdd vss bl[405] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_406 br[405] vdd vss bl[405] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_406 br[405] vdd vss bl[405] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_406 br[405] vdd vss bl[405] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_406 br[405] vdd vss bl[405] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_406 br[405] vdd vss bl[405] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_407 br[406] vdd vss bl[406] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_407 br[406] vdd vss bl[406] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_407 br[406] vdd vss bl[406] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_407 br[406] vdd vss bl[406] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_407 br[406] vdd vss bl[406] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_407 br[406] vdd vss bl[406] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_407 br[406] vdd vss bl[406] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_407 br[406] vdd vss bl[406] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_407 br[406] vdd vss bl[406] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_407 br[406] vdd vss bl[406] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_407 br[406] vdd vss bl[406] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_407 br[406] vdd vss bl[406] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_407 br[406] vdd vss bl[406] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_407 br[406] vdd vss bl[406] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_407 br[406] vdd vss bl[406] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_407 br[406] vdd vss bl[406] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_407 br[406] vdd vss bl[406] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_407 br[406] vdd vss bl[406] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_407 br[406] vdd vss bl[406] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_408 br[407] vdd vss bl[407] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_408 br[407] vdd vss bl[407] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_408 br[407] vdd vss bl[407] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_408 br[407] vdd vss bl[407] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_408 br[407] vdd vss bl[407] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_408 br[407] vdd vss bl[407] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_408 br[407] vdd vss bl[407] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_408 br[407] vdd vss bl[407] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_408 br[407] vdd vss bl[407] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_408 br[407] vdd vss bl[407] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_408 br[407] vdd vss bl[407] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_408 br[407] vdd vss bl[407] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_408 br[407] vdd vss bl[407] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_408 br[407] vdd vss bl[407] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_408 br[407] vdd vss bl[407] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_408 br[407] vdd vss bl[407] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_408 br[407] vdd vss bl[407] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_408 br[407] vdd vss bl[407] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_408 br[407] vdd vss bl[407] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_409 br[408] vdd vss bl[408] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_409 br[408] vdd vss bl[408] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_409 br[408] vdd vss bl[408] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_409 br[408] vdd vss bl[408] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_409 br[408] vdd vss bl[408] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_409 br[408] vdd vss bl[408] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_409 br[408] vdd vss bl[408] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_409 br[408] vdd vss bl[408] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_409 br[408] vdd vss bl[408] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_409 br[408] vdd vss bl[408] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_409 br[408] vdd vss bl[408] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_409 br[408] vdd vss bl[408] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_409 br[408] vdd vss bl[408] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_409 br[408] vdd vss bl[408] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_409 br[408] vdd vss bl[408] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_409 br[408] vdd vss bl[408] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_409 br[408] vdd vss bl[408] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_409 br[408] vdd vss bl[408] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_409 br[408] vdd vss bl[408] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_410 br[409] vdd vss bl[409] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_410 br[409] vdd vss bl[409] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_410 br[409] vdd vss bl[409] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_410 br[409] vdd vss bl[409] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_410 br[409] vdd vss bl[409] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_410 br[409] vdd vss bl[409] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_410 br[409] vdd vss bl[409] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_410 br[409] vdd vss bl[409] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_410 br[409] vdd vss bl[409] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_410 br[409] vdd vss bl[409] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_410 br[409] vdd vss bl[409] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_410 br[409] vdd vss bl[409] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_410 br[409] vdd vss bl[409] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_410 br[409] vdd vss bl[409] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_410 br[409] vdd vss bl[409] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_410 br[409] vdd vss bl[409] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_410 br[409] vdd vss bl[409] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_410 br[409] vdd vss bl[409] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_410 br[409] vdd vss bl[409] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_411 br[410] vdd vss bl[410] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_411 br[410] vdd vss bl[410] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_411 br[410] vdd vss bl[410] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_411 br[410] vdd vss bl[410] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_411 br[410] vdd vss bl[410] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_411 br[410] vdd vss bl[410] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_411 br[410] vdd vss bl[410] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_411 br[410] vdd vss bl[410] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_411 br[410] vdd vss bl[410] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_411 br[410] vdd vss bl[410] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_411 br[410] vdd vss bl[410] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_411 br[410] vdd vss bl[410] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_411 br[410] vdd vss bl[410] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_411 br[410] vdd vss bl[410] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_411 br[410] vdd vss bl[410] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_411 br[410] vdd vss bl[410] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_411 br[410] vdd vss bl[410] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_411 br[410] vdd vss bl[410] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_411 br[410] vdd vss bl[410] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_412 br[411] vdd vss bl[411] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_412 br[411] vdd vss bl[411] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_412 br[411] vdd vss bl[411] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_412 br[411] vdd vss bl[411] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_412 br[411] vdd vss bl[411] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_412 br[411] vdd vss bl[411] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_412 br[411] vdd vss bl[411] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_412 br[411] vdd vss bl[411] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_412 br[411] vdd vss bl[411] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_412 br[411] vdd vss bl[411] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_412 br[411] vdd vss bl[411] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_412 br[411] vdd vss bl[411] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_412 br[411] vdd vss bl[411] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_412 br[411] vdd vss bl[411] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_412 br[411] vdd vss bl[411] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_412 br[411] vdd vss bl[411] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_412 br[411] vdd vss bl[411] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_412 br[411] vdd vss bl[411] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_412 br[411] vdd vss bl[411] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_413 br[412] vdd vss bl[412] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_413 br[412] vdd vss bl[412] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_413 br[412] vdd vss bl[412] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_413 br[412] vdd vss bl[412] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_413 br[412] vdd vss bl[412] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_413 br[412] vdd vss bl[412] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_413 br[412] vdd vss bl[412] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_413 br[412] vdd vss bl[412] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_413 br[412] vdd vss bl[412] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_413 br[412] vdd vss bl[412] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_413 br[412] vdd vss bl[412] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_413 br[412] vdd vss bl[412] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_413 br[412] vdd vss bl[412] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_413 br[412] vdd vss bl[412] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_413 br[412] vdd vss bl[412] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_413 br[412] vdd vss bl[412] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_413 br[412] vdd vss bl[412] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_413 br[412] vdd vss bl[412] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_413 br[412] vdd vss bl[412] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_414 br[413] vdd vss bl[413] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_414 br[413] vdd vss bl[413] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_414 br[413] vdd vss bl[413] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_414 br[413] vdd vss bl[413] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_414 br[413] vdd vss bl[413] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_414 br[413] vdd vss bl[413] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_414 br[413] vdd vss bl[413] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_414 br[413] vdd vss bl[413] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_414 br[413] vdd vss bl[413] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_414 br[413] vdd vss bl[413] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_414 br[413] vdd vss bl[413] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_414 br[413] vdd vss bl[413] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_414 br[413] vdd vss bl[413] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_414 br[413] vdd vss bl[413] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_414 br[413] vdd vss bl[413] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_414 br[413] vdd vss bl[413] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_414 br[413] vdd vss bl[413] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_414 br[413] vdd vss bl[413] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_414 br[413] vdd vss bl[413] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_415 br[414] vdd vss bl[414] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_415 br[414] vdd vss bl[414] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_415 br[414] vdd vss bl[414] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_415 br[414] vdd vss bl[414] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_415 br[414] vdd vss bl[414] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_415 br[414] vdd vss bl[414] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_415 br[414] vdd vss bl[414] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_415 br[414] vdd vss bl[414] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_415 br[414] vdd vss bl[414] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_415 br[414] vdd vss bl[414] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_415 br[414] vdd vss bl[414] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_415 br[414] vdd vss bl[414] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_415 br[414] vdd vss bl[414] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_415 br[414] vdd vss bl[414] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_415 br[414] vdd vss bl[414] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_415 br[414] vdd vss bl[414] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_415 br[414] vdd vss bl[414] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_415 br[414] vdd vss bl[414] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_415 br[414] vdd vss bl[414] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_416 br[415] vdd vss bl[415] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_416 br[415] vdd vss bl[415] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_416 br[415] vdd vss bl[415] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_416 br[415] vdd vss bl[415] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_416 br[415] vdd vss bl[415] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_416 br[415] vdd vss bl[415] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_416 br[415] vdd vss bl[415] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_416 br[415] vdd vss bl[415] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_416 br[415] vdd vss bl[415] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_416 br[415] vdd vss bl[415] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_416 br[415] vdd vss bl[415] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_416 br[415] vdd vss bl[415] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_416 br[415] vdd vss bl[415] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_416 br[415] vdd vss bl[415] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_416 br[415] vdd vss bl[415] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_416 br[415] vdd vss bl[415] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_416 br[415] vdd vss bl[415] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_416 br[415] vdd vss bl[415] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_416 br[415] vdd vss bl[415] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_417 br[416] vdd vss bl[416] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_417 br[416] vdd vss bl[416] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_417 br[416] vdd vss bl[416] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_417 br[416] vdd vss bl[416] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_417 br[416] vdd vss bl[416] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_417 br[416] vdd vss bl[416] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_417 br[416] vdd vss bl[416] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_417 br[416] vdd vss bl[416] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_417 br[416] vdd vss bl[416] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_417 br[416] vdd vss bl[416] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_417 br[416] vdd vss bl[416] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_417 br[416] vdd vss bl[416] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_417 br[416] vdd vss bl[416] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_417 br[416] vdd vss bl[416] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_417 br[416] vdd vss bl[416] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_417 br[416] vdd vss bl[416] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_417 br[416] vdd vss bl[416] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_417 br[416] vdd vss bl[416] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_417 br[416] vdd vss bl[416] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_418 br[417] vdd vss bl[417] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_418 br[417] vdd vss bl[417] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_418 br[417] vdd vss bl[417] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_418 br[417] vdd vss bl[417] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_418 br[417] vdd vss bl[417] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_418 br[417] vdd vss bl[417] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_418 br[417] vdd vss bl[417] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_418 br[417] vdd vss bl[417] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_418 br[417] vdd vss bl[417] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_418 br[417] vdd vss bl[417] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_418 br[417] vdd vss bl[417] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_418 br[417] vdd vss bl[417] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_418 br[417] vdd vss bl[417] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_418 br[417] vdd vss bl[417] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_418 br[417] vdd vss bl[417] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_418 br[417] vdd vss bl[417] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_418 br[417] vdd vss bl[417] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_418 br[417] vdd vss bl[417] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_418 br[417] vdd vss bl[417] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_419 br[418] vdd vss bl[418] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_419 br[418] vdd vss bl[418] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_419 br[418] vdd vss bl[418] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_419 br[418] vdd vss bl[418] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_419 br[418] vdd vss bl[418] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_419 br[418] vdd vss bl[418] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_419 br[418] vdd vss bl[418] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_419 br[418] vdd vss bl[418] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_419 br[418] vdd vss bl[418] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_419 br[418] vdd vss bl[418] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_419 br[418] vdd vss bl[418] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_419 br[418] vdd vss bl[418] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_419 br[418] vdd vss bl[418] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_419 br[418] vdd vss bl[418] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_419 br[418] vdd vss bl[418] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_419 br[418] vdd vss bl[418] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_419 br[418] vdd vss bl[418] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_419 br[418] vdd vss bl[418] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_419 br[418] vdd vss bl[418] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_420 br[419] vdd vss bl[419] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_420 br[419] vdd vss bl[419] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_420 br[419] vdd vss bl[419] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_420 br[419] vdd vss bl[419] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_420 br[419] vdd vss bl[419] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_420 br[419] vdd vss bl[419] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_420 br[419] vdd vss bl[419] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_420 br[419] vdd vss bl[419] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_420 br[419] vdd vss bl[419] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_420 br[419] vdd vss bl[419] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_420 br[419] vdd vss bl[419] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_420 br[419] vdd vss bl[419] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_420 br[419] vdd vss bl[419] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_420 br[419] vdd vss bl[419] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_420 br[419] vdd vss bl[419] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_420 br[419] vdd vss bl[419] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_420 br[419] vdd vss bl[419] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_420 br[419] vdd vss bl[419] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_420 br[419] vdd vss bl[419] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_421 br[420] vdd vss bl[420] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_421 br[420] vdd vss bl[420] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_421 br[420] vdd vss bl[420] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_421 br[420] vdd vss bl[420] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_421 br[420] vdd vss bl[420] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_421 br[420] vdd vss bl[420] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_421 br[420] vdd vss bl[420] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_421 br[420] vdd vss bl[420] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_421 br[420] vdd vss bl[420] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_421 br[420] vdd vss bl[420] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_421 br[420] vdd vss bl[420] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_421 br[420] vdd vss bl[420] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_421 br[420] vdd vss bl[420] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_421 br[420] vdd vss bl[420] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_421 br[420] vdd vss bl[420] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_421 br[420] vdd vss bl[420] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_421 br[420] vdd vss bl[420] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_421 br[420] vdd vss bl[420] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_421 br[420] vdd vss bl[420] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_422 br[421] vdd vss bl[421] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_422 br[421] vdd vss bl[421] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_422 br[421] vdd vss bl[421] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_422 br[421] vdd vss bl[421] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_422 br[421] vdd vss bl[421] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_422 br[421] vdd vss bl[421] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_422 br[421] vdd vss bl[421] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_422 br[421] vdd vss bl[421] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_422 br[421] vdd vss bl[421] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_422 br[421] vdd vss bl[421] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_422 br[421] vdd vss bl[421] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_422 br[421] vdd vss bl[421] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_422 br[421] vdd vss bl[421] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_422 br[421] vdd vss bl[421] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_422 br[421] vdd vss bl[421] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_422 br[421] vdd vss bl[421] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_422 br[421] vdd vss bl[421] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_422 br[421] vdd vss bl[421] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_422 br[421] vdd vss bl[421] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_423 br[422] vdd vss bl[422] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_423 br[422] vdd vss bl[422] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_423 br[422] vdd vss bl[422] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_423 br[422] vdd vss bl[422] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_423 br[422] vdd vss bl[422] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_423 br[422] vdd vss bl[422] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_423 br[422] vdd vss bl[422] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_423 br[422] vdd vss bl[422] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_423 br[422] vdd vss bl[422] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_423 br[422] vdd vss bl[422] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_423 br[422] vdd vss bl[422] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_423 br[422] vdd vss bl[422] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_423 br[422] vdd vss bl[422] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_423 br[422] vdd vss bl[422] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_423 br[422] vdd vss bl[422] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_423 br[422] vdd vss bl[422] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_423 br[422] vdd vss bl[422] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_423 br[422] vdd vss bl[422] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_423 br[422] vdd vss bl[422] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_424 br[423] vdd vss bl[423] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_424 br[423] vdd vss bl[423] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_424 br[423] vdd vss bl[423] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_424 br[423] vdd vss bl[423] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_424 br[423] vdd vss bl[423] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_424 br[423] vdd vss bl[423] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_424 br[423] vdd vss bl[423] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_424 br[423] vdd vss bl[423] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_424 br[423] vdd vss bl[423] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_424 br[423] vdd vss bl[423] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_424 br[423] vdd vss bl[423] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_424 br[423] vdd vss bl[423] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_424 br[423] vdd vss bl[423] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_424 br[423] vdd vss bl[423] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_424 br[423] vdd vss bl[423] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_424 br[423] vdd vss bl[423] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_424 br[423] vdd vss bl[423] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_424 br[423] vdd vss bl[423] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_424 br[423] vdd vss bl[423] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_425 br[424] vdd vss bl[424] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_425 br[424] vdd vss bl[424] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_425 br[424] vdd vss bl[424] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_425 br[424] vdd vss bl[424] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_425 br[424] vdd vss bl[424] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_425 br[424] vdd vss bl[424] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_425 br[424] vdd vss bl[424] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_425 br[424] vdd vss bl[424] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_425 br[424] vdd vss bl[424] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_425 br[424] vdd vss bl[424] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_425 br[424] vdd vss bl[424] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_425 br[424] vdd vss bl[424] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_425 br[424] vdd vss bl[424] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_425 br[424] vdd vss bl[424] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_425 br[424] vdd vss bl[424] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_425 br[424] vdd vss bl[424] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_425 br[424] vdd vss bl[424] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_425 br[424] vdd vss bl[424] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_425 br[424] vdd vss bl[424] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_426 br[425] vdd vss bl[425] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_426 br[425] vdd vss bl[425] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_426 br[425] vdd vss bl[425] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_426 br[425] vdd vss bl[425] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_426 br[425] vdd vss bl[425] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_426 br[425] vdd vss bl[425] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_426 br[425] vdd vss bl[425] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_426 br[425] vdd vss bl[425] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_426 br[425] vdd vss bl[425] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_426 br[425] vdd vss bl[425] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_426 br[425] vdd vss bl[425] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_426 br[425] vdd vss bl[425] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_426 br[425] vdd vss bl[425] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_426 br[425] vdd vss bl[425] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_426 br[425] vdd vss bl[425] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_426 br[425] vdd vss bl[425] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_426 br[425] vdd vss bl[425] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_426 br[425] vdd vss bl[425] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_426 br[425] vdd vss bl[425] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_427 br[426] vdd vss bl[426] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_427 br[426] vdd vss bl[426] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_427 br[426] vdd vss bl[426] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_427 br[426] vdd vss bl[426] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_427 br[426] vdd vss bl[426] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_427 br[426] vdd vss bl[426] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_427 br[426] vdd vss bl[426] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_427 br[426] vdd vss bl[426] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_427 br[426] vdd vss bl[426] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_427 br[426] vdd vss bl[426] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_427 br[426] vdd vss bl[426] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_427 br[426] vdd vss bl[426] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_427 br[426] vdd vss bl[426] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_427 br[426] vdd vss bl[426] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_427 br[426] vdd vss bl[426] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_427 br[426] vdd vss bl[426] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_427 br[426] vdd vss bl[426] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_427 br[426] vdd vss bl[426] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_427 br[426] vdd vss bl[426] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_428 br[427] vdd vss bl[427] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_428 br[427] vdd vss bl[427] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_428 br[427] vdd vss bl[427] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_428 br[427] vdd vss bl[427] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_428 br[427] vdd vss bl[427] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_428 br[427] vdd vss bl[427] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_428 br[427] vdd vss bl[427] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_428 br[427] vdd vss bl[427] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_428 br[427] vdd vss bl[427] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_428 br[427] vdd vss bl[427] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_428 br[427] vdd vss bl[427] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_428 br[427] vdd vss bl[427] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_428 br[427] vdd vss bl[427] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_428 br[427] vdd vss bl[427] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_428 br[427] vdd vss bl[427] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_428 br[427] vdd vss bl[427] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_428 br[427] vdd vss bl[427] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_428 br[427] vdd vss bl[427] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_428 br[427] vdd vss bl[427] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_429 br[428] vdd vss bl[428] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_429 br[428] vdd vss bl[428] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_429 br[428] vdd vss bl[428] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_429 br[428] vdd vss bl[428] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_429 br[428] vdd vss bl[428] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_429 br[428] vdd vss bl[428] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_429 br[428] vdd vss bl[428] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_429 br[428] vdd vss bl[428] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_429 br[428] vdd vss bl[428] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_429 br[428] vdd vss bl[428] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_429 br[428] vdd vss bl[428] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_429 br[428] vdd vss bl[428] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_429 br[428] vdd vss bl[428] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_429 br[428] vdd vss bl[428] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_429 br[428] vdd vss bl[428] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_429 br[428] vdd vss bl[428] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_429 br[428] vdd vss bl[428] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_429 br[428] vdd vss bl[428] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_429 br[428] vdd vss bl[428] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_430 br[429] vdd vss bl[429] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_430 br[429] vdd vss bl[429] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_430 br[429] vdd vss bl[429] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_430 br[429] vdd vss bl[429] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_430 br[429] vdd vss bl[429] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_430 br[429] vdd vss bl[429] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_430 br[429] vdd vss bl[429] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_430 br[429] vdd vss bl[429] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_430 br[429] vdd vss bl[429] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_430 br[429] vdd vss bl[429] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_430 br[429] vdd vss bl[429] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_430 br[429] vdd vss bl[429] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_430 br[429] vdd vss bl[429] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_430 br[429] vdd vss bl[429] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_430 br[429] vdd vss bl[429] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_430 br[429] vdd vss bl[429] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_430 br[429] vdd vss bl[429] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_430 br[429] vdd vss bl[429] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_430 br[429] vdd vss bl[429] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_431 br[430] vdd vss bl[430] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_431 br[430] vdd vss bl[430] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_431 br[430] vdd vss bl[430] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_431 br[430] vdd vss bl[430] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_431 br[430] vdd vss bl[430] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_431 br[430] vdd vss bl[430] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_431 br[430] vdd vss bl[430] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_431 br[430] vdd vss bl[430] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_431 br[430] vdd vss bl[430] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_431 br[430] vdd vss bl[430] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_431 br[430] vdd vss bl[430] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_431 br[430] vdd vss bl[430] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_431 br[430] vdd vss bl[430] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_431 br[430] vdd vss bl[430] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_431 br[430] vdd vss bl[430] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_431 br[430] vdd vss bl[430] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_431 br[430] vdd vss bl[430] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_431 br[430] vdd vss bl[430] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_431 br[430] vdd vss bl[430] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_432 br[431] vdd vss bl[431] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_432 br[431] vdd vss bl[431] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_432 br[431] vdd vss bl[431] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_432 br[431] vdd vss bl[431] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_432 br[431] vdd vss bl[431] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_432 br[431] vdd vss bl[431] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_432 br[431] vdd vss bl[431] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_432 br[431] vdd vss bl[431] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_432 br[431] vdd vss bl[431] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_432 br[431] vdd vss bl[431] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_432 br[431] vdd vss bl[431] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_432 br[431] vdd vss bl[431] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_432 br[431] vdd vss bl[431] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_432 br[431] vdd vss bl[431] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_432 br[431] vdd vss bl[431] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_432 br[431] vdd vss bl[431] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_432 br[431] vdd vss bl[431] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_432 br[431] vdd vss bl[431] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_432 br[431] vdd vss bl[431] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_433 br[432] vdd vss bl[432] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_433 br[432] vdd vss bl[432] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_433 br[432] vdd vss bl[432] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_433 br[432] vdd vss bl[432] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_433 br[432] vdd vss bl[432] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_433 br[432] vdd vss bl[432] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_433 br[432] vdd vss bl[432] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_433 br[432] vdd vss bl[432] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_433 br[432] vdd vss bl[432] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_433 br[432] vdd vss bl[432] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_433 br[432] vdd vss bl[432] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_433 br[432] vdd vss bl[432] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_433 br[432] vdd vss bl[432] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_433 br[432] vdd vss bl[432] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_433 br[432] vdd vss bl[432] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_433 br[432] vdd vss bl[432] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_433 br[432] vdd vss bl[432] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_433 br[432] vdd vss bl[432] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_433 br[432] vdd vss bl[432] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_434 br[433] vdd vss bl[433] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_434 br[433] vdd vss bl[433] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_434 br[433] vdd vss bl[433] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_434 br[433] vdd vss bl[433] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_434 br[433] vdd vss bl[433] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_434 br[433] vdd vss bl[433] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_434 br[433] vdd vss bl[433] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_434 br[433] vdd vss bl[433] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_434 br[433] vdd vss bl[433] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_434 br[433] vdd vss bl[433] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_434 br[433] vdd vss bl[433] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_434 br[433] vdd vss bl[433] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_434 br[433] vdd vss bl[433] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_434 br[433] vdd vss bl[433] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_434 br[433] vdd vss bl[433] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_434 br[433] vdd vss bl[433] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_434 br[433] vdd vss bl[433] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_434 br[433] vdd vss bl[433] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_434 br[433] vdd vss bl[433] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_435 br[434] vdd vss bl[434] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_435 br[434] vdd vss bl[434] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_435 br[434] vdd vss bl[434] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_435 br[434] vdd vss bl[434] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_435 br[434] vdd vss bl[434] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_435 br[434] vdd vss bl[434] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_435 br[434] vdd vss bl[434] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_435 br[434] vdd vss bl[434] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_435 br[434] vdd vss bl[434] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_435 br[434] vdd vss bl[434] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_435 br[434] vdd vss bl[434] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_435 br[434] vdd vss bl[434] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_435 br[434] vdd vss bl[434] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_435 br[434] vdd vss bl[434] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_435 br[434] vdd vss bl[434] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_435 br[434] vdd vss bl[434] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_435 br[434] vdd vss bl[434] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_435 br[434] vdd vss bl[434] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_435 br[434] vdd vss bl[434] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_436 br[435] vdd vss bl[435] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_436 br[435] vdd vss bl[435] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_436 br[435] vdd vss bl[435] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_436 br[435] vdd vss bl[435] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_436 br[435] vdd vss bl[435] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_436 br[435] vdd vss bl[435] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_436 br[435] vdd vss bl[435] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_436 br[435] vdd vss bl[435] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_436 br[435] vdd vss bl[435] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_436 br[435] vdd vss bl[435] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_436 br[435] vdd vss bl[435] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_436 br[435] vdd vss bl[435] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_436 br[435] vdd vss bl[435] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_436 br[435] vdd vss bl[435] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_436 br[435] vdd vss bl[435] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_436 br[435] vdd vss bl[435] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_436 br[435] vdd vss bl[435] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_436 br[435] vdd vss bl[435] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_436 br[435] vdd vss bl[435] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_437 br[436] vdd vss bl[436] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_437 br[436] vdd vss bl[436] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_437 br[436] vdd vss bl[436] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_437 br[436] vdd vss bl[436] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_437 br[436] vdd vss bl[436] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_437 br[436] vdd vss bl[436] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_437 br[436] vdd vss bl[436] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_437 br[436] vdd vss bl[436] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_437 br[436] vdd vss bl[436] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_437 br[436] vdd vss bl[436] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_437 br[436] vdd vss bl[436] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_437 br[436] vdd vss bl[436] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_437 br[436] vdd vss bl[436] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_437 br[436] vdd vss bl[436] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_437 br[436] vdd vss bl[436] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_437 br[436] vdd vss bl[436] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_437 br[436] vdd vss bl[436] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_437 br[436] vdd vss bl[436] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_437 br[436] vdd vss bl[436] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_438 br[437] vdd vss bl[437] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_438 br[437] vdd vss bl[437] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_438 br[437] vdd vss bl[437] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_438 br[437] vdd vss bl[437] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_438 br[437] vdd vss bl[437] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_438 br[437] vdd vss bl[437] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_438 br[437] vdd vss bl[437] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_438 br[437] vdd vss bl[437] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_438 br[437] vdd vss bl[437] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_438 br[437] vdd vss bl[437] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_438 br[437] vdd vss bl[437] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_438 br[437] vdd vss bl[437] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_438 br[437] vdd vss bl[437] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_438 br[437] vdd vss bl[437] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_438 br[437] vdd vss bl[437] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_438 br[437] vdd vss bl[437] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_438 br[437] vdd vss bl[437] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_438 br[437] vdd vss bl[437] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_438 br[437] vdd vss bl[437] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_439 br[438] vdd vss bl[438] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_439 br[438] vdd vss bl[438] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_439 br[438] vdd vss bl[438] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_439 br[438] vdd vss bl[438] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_439 br[438] vdd vss bl[438] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_439 br[438] vdd vss bl[438] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_439 br[438] vdd vss bl[438] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_439 br[438] vdd vss bl[438] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_439 br[438] vdd vss bl[438] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_439 br[438] vdd vss bl[438] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_439 br[438] vdd vss bl[438] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_439 br[438] vdd vss bl[438] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_439 br[438] vdd vss bl[438] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_439 br[438] vdd vss bl[438] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_439 br[438] vdd vss bl[438] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_439 br[438] vdd vss bl[438] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_439 br[438] vdd vss bl[438] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_439 br[438] vdd vss bl[438] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_439 br[438] vdd vss bl[438] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_440 br[439] vdd vss bl[439] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_440 br[439] vdd vss bl[439] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_440 br[439] vdd vss bl[439] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_440 br[439] vdd vss bl[439] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_440 br[439] vdd vss bl[439] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_440 br[439] vdd vss bl[439] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_440 br[439] vdd vss bl[439] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_440 br[439] vdd vss bl[439] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_440 br[439] vdd vss bl[439] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_440 br[439] vdd vss bl[439] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_440 br[439] vdd vss bl[439] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_440 br[439] vdd vss bl[439] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_440 br[439] vdd vss bl[439] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_440 br[439] vdd vss bl[439] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_440 br[439] vdd vss bl[439] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_440 br[439] vdd vss bl[439] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_440 br[439] vdd vss bl[439] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_440 br[439] vdd vss bl[439] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_440 br[439] vdd vss bl[439] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_441 br[440] vdd vss bl[440] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_441 br[440] vdd vss bl[440] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_441 br[440] vdd vss bl[440] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_441 br[440] vdd vss bl[440] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_441 br[440] vdd vss bl[440] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_441 br[440] vdd vss bl[440] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_441 br[440] vdd vss bl[440] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_441 br[440] vdd vss bl[440] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_441 br[440] vdd vss bl[440] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_441 br[440] vdd vss bl[440] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_441 br[440] vdd vss bl[440] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_441 br[440] vdd vss bl[440] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_441 br[440] vdd vss bl[440] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_441 br[440] vdd vss bl[440] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_441 br[440] vdd vss bl[440] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_441 br[440] vdd vss bl[440] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_441 br[440] vdd vss bl[440] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_441 br[440] vdd vss bl[440] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_441 br[440] vdd vss bl[440] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_442 br[441] vdd vss bl[441] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_442 br[441] vdd vss bl[441] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_442 br[441] vdd vss bl[441] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_442 br[441] vdd vss bl[441] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_442 br[441] vdd vss bl[441] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_442 br[441] vdd vss bl[441] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_442 br[441] vdd vss bl[441] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_442 br[441] vdd vss bl[441] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_442 br[441] vdd vss bl[441] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_442 br[441] vdd vss bl[441] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_442 br[441] vdd vss bl[441] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_442 br[441] vdd vss bl[441] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_442 br[441] vdd vss bl[441] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_442 br[441] vdd vss bl[441] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_442 br[441] vdd vss bl[441] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_442 br[441] vdd vss bl[441] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_442 br[441] vdd vss bl[441] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_442 br[441] vdd vss bl[441] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_442 br[441] vdd vss bl[441] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_443 br[442] vdd vss bl[442] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_443 br[442] vdd vss bl[442] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_443 br[442] vdd vss bl[442] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_443 br[442] vdd vss bl[442] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_443 br[442] vdd vss bl[442] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_443 br[442] vdd vss bl[442] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_443 br[442] vdd vss bl[442] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_443 br[442] vdd vss bl[442] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_443 br[442] vdd vss bl[442] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_443 br[442] vdd vss bl[442] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_443 br[442] vdd vss bl[442] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_443 br[442] vdd vss bl[442] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_443 br[442] vdd vss bl[442] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_443 br[442] vdd vss bl[442] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_443 br[442] vdd vss bl[442] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_443 br[442] vdd vss bl[442] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_443 br[442] vdd vss bl[442] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_443 br[442] vdd vss bl[442] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_443 br[442] vdd vss bl[442] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_444 br[443] vdd vss bl[443] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_444 br[443] vdd vss bl[443] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_444 br[443] vdd vss bl[443] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_444 br[443] vdd vss bl[443] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_444 br[443] vdd vss bl[443] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_444 br[443] vdd vss bl[443] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_444 br[443] vdd vss bl[443] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_444 br[443] vdd vss bl[443] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_444 br[443] vdd vss bl[443] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_444 br[443] vdd vss bl[443] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_444 br[443] vdd vss bl[443] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_444 br[443] vdd vss bl[443] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_444 br[443] vdd vss bl[443] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_444 br[443] vdd vss bl[443] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_444 br[443] vdd vss bl[443] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_444 br[443] vdd vss bl[443] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_444 br[443] vdd vss bl[443] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_444 br[443] vdd vss bl[443] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_444 br[443] vdd vss bl[443] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_445 br[444] vdd vss bl[444] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_445 br[444] vdd vss bl[444] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_445 br[444] vdd vss bl[444] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_445 br[444] vdd vss bl[444] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_445 br[444] vdd vss bl[444] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_445 br[444] vdd vss bl[444] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_445 br[444] vdd vss bl[444] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_445 br[444] vdd vss bl[444] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_445 br[444] vdd vss bl[444] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_445 br[444] vdd vss bl[444] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_445 br[444] vdd vss bl[444] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_445 br[444] vdd vss bl[444] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_445 br[444] vdd vss bl[444] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_445 br[444] vdd vss bl[444] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_445 br[444] vdd vss bl[444] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_445 br[444] vdd vss bl[444] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_445 br[444] vdd vss bl[444] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_445 br[444] vdd vss bl[444] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_445 br[444] vdd vss bl[444] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_446 br[445] vdd vss bl[445] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_446 br[445] vdd vss bl[445] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_446 br[445] vdd vss bl[445] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_446 br[445] vdd vss bl[445] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_446 br[445] vdd vss bl[445] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_446 br[445] vdd vss bl[445] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_446 br[445] vdd vss bl[445] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_446 br[445] vdd vss bl[445] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_446 br[445] vdd vss bl[445] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_446 br[445] vdd vss bl[445] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_446 br[445] vdd vss bl[445] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_446 br[445] vdd vss bl[445] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_446 br[445] vdd vss bl[445] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_446 br[445] vdd vss bl[445] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_446 br[445] vdd vss bl[445] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_446 br[445] vdd vss bl[445] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_446 br[445] vdd vss bl[445] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_446 br[445] vdd vss bl[445] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_446 br[445] vdd vss bl[445] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_447 br[446] vdd vss bl[446] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_447 br[446] vdd vss bl[446] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_447 br[446] vdd vss bl[446] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_447 br[446] vdd vss bl[446] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_447 br[446] vdd vss bl[446] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_447 br[446] vdd vss bl[446] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_447 br[446] vdd vss bl[446] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_447 br[446] vdd vss bl[446] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_447 br[446] vdd vss bl[446] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_447 br[446] vdd vss bl[446] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_447 br[446] vdd vss bl[446] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_447 br[446] vdd vss bl[446] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_447 br[446] vdd vss bl[446] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_447 br[446] vdd vss bl[446] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_447 br[446] vdd vss bl[446] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_447 br[446] vdd vss bl[446] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_447 br[446] vdd vss bl[446] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_447 br[446] vdd vss bl[446] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_447 br[446] vdd vss bl[446] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_448 br[447] vdd vss bl[447] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_448 br[447] vdd vss bl[447] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_448 br[447] vdd vss bl[447] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_448 br[447] vdd vss bl[447] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_448 br[447] vdd vss bl[447] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_448 br[447] vdd vss bl[447] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_448 br[447] vdd vss bl[447] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_448 br[447] vdd vss bl[447] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_448 br[447] vdd vss bl[447] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_448 br[447] vdd vss bl[447] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_448 br[447] vdd vss bl[447] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_448 br[447] vdd vss bl[447] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_448 br[447] vdd vss bl[447] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_448 br[447] vdd vss bl[447] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_448 br[447] vdd vss bl[447] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_448 br[447] vdd vss bl[447] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_448 br[447] vdd vss bl[447] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_448 br[447] vdd vss bl[447] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_448 br[447] vdd vss bl[447] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_449 br[448] vdd vss bl[448] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_449 br[448] vdd vss bl[448] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_449 br[448] vdd vss bl[448] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_449 br[448] vdd vss bl[448] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_449 br[448] vdd vss bl[448] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_449 br[448] vdd vss bl[448] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_449 br[448] vdd vss bl[448] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_449 br[448] vdd vss bl[448] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_449 br[448] vdd vss bl[448] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_449 br[448] vdd vss bl[448] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_449 br[448] vdd vss bl[448] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_449 br[448] vdd vss bl[448] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_449 br[448] vdd vss bl[448] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_449 br[448] vdd vss bl[448] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_449 br[448] vdd vss bl[448] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_449 br[448] vdd vss bl[448] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_449 br[448] vdd vss bl[448] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_449 br[448] vdd vss bl[448] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_449 br[448] vdd vss bl[448] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_450 br[449] vdd vss bl[449] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_450 br[449] vdd vss bl[449] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_450 br[449] vdd vss bl[449] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_450 br[449] vdd vss bl[449] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_450 br[449] vdd vss bl[449] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_450 br[449] vdd vss bl[449] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_450 br[449] vdd vss bl[449] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_450 br[449] vdd vss bl[449] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_450 br[449] vdd vss bl[449] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_450 br[449] vdd vss bl[449] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_450 br[449] vdd vss bl[449] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_450 br[449] vdd vss bl[449] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_450 br[449] vdd vss bl[449] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_450 br[449] vdd vss bl[449] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_450 br[449] vdd vss bl[449] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_450 br[449] vdd vss bl[449] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_450 br[449] vdd vss bl[449] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_450 br[449] vdd vss bl[449] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_450 br[449] vdd vss bl[449] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_451 br[450] vdd vss bl[450] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_451 br[450] vdd vss bl[450] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_451 br[450] vdd vss bl[450] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_451 br[450] vdd vss bl[450] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_451 br[450] vdd vss bl[450] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_451 br[450] vdd vss bl[450] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_451 br[450] vdd vss bl[450] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_451 br[450] vdd vss bl[450] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_451 br[450] vdd vss bl[450] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_451 br[450] vdd vss bl[450] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_451 br[450] vdd vss bl[450] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_451 br[450] vdd vss bl[450] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_451 br[450] vdd vss bl[450] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_451 br[450] vdd vss bl[450] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_451 br[450] vdd vss bl[450] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_451 br[450] vdd vss bl[450] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_451 br[450] vdd vss bl[450] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_451 br[450] vdd vss bl[450] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_451 br[450] vdd vss bl[450] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_452 br[451] vdd vss bl[451] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_452 br[451] vdd vss bl[451] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_452 br[451] vdd vss bl[451] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_452 br[451] vdd vss bl[451] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_452 br[451] vdd vss bl[451] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_452 br[451] vdd vss bl[451] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_452 br[451] vdd vss bl[451] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_452 br[451] vdd vss bl[451] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_452 br[451] vdd vss bl[451] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_452 br[451] vdd vss bl[451] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_452 br[451] vdd vss bl[451] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_452 br[451] vdd vss bl[451] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_452 br[451] vdd vss bl[451] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_452 br[451] vdd vss bl[451] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_452 br[451] vdd vss bl[451] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_452 br[451] vdd vss bl[451] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_452 br[451] vdd vss bl[451] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_452 br[451] vdd vss bl[451] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_452 br[451] vdd vss bl[451] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_453 br[452] vdd vss bl[452] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_453 br[452] vdd vss bl[452] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_453 br[452] vdd vss bl[452] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_453 br[452] vdd vss bl[452] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_453 br[452] vdd vss bl[452] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_453 br[452] vdd vss bl[452] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_453 br[452] vdd vss bl[452] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_453 br[452] vdd vss bl[452] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_453 br[452] vdd vss bl[452] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_453 br[452] vdd vss bl[452] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_453 br[452] vdd vss bl[452] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_453 br[452] vdd vss bl[452] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_453 br[452] vdd vss bl[452] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_453 br[452] vdd vss bl[452] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_453 br[452] vdd vss bl[452] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_453 br[452] vdd vss bl[452] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_453 br[452] vdd vss bl[452] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_453 br[452] vdd vss bl[452] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_453 br[452] vdd vss bl[452] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_454 br[453] vdd vss bl[453] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_454 br[453] vdd vss bl[453] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_454 br[453] vdd vss bl[453] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_454 br[453] vdd vss bl[453] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_454 br[453] vdd vss bl[453] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_454 br[453] vdd vss bl[453] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_454 br[453] vdd vss bl[453] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_454 br[453] vdd vss bl[453] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_454 br[453] vdd vss bl[453] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_454 br[453] vdd vss bl[453] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_454 br[453] vdd vss bl[453] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_454 br[453] vdd vss bl[453] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_454 br[453] vdd vss bl[453] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_454 br[453] vdd vss bl[453] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_454 br[453] vdd vss bl[453] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_454 br[453] vdd vss bl[453] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_454 br[453] vdd vss bl[453] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_454 br[453] vdd vss bl[453] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_454 br[453] vdd vss bl[453] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_455 br[454] vdd vss bl[454] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_455 br[454] vdd vss bl[454] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_455 br[454] vdd vss bl[454] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_455 br[454] vdd vss bl[454] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_455 br[454] vdd vss bl[454] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_455 br[454] vdd vss bl[454] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_455 br[454] vdd vss bl[454] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_455 br[454] vdd vss bl[454] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_455 br[454] vdd vss bl[454] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_455 br[454] vdd vss bl[454] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_455 br[454] vdd vss bl[454] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_455 br[454] vdd vss bl[454] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_455 br[454] vdd vss bl[454] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_455 br[454] vdd vss bl[454] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_455 br[454] vdd vss bl[454] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_455 br[454] vdd vss bl[454] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_455 br[454] vdd vss bl[454] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_455 br[454] vdd vss bl[454] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_455 br[454] vdd vss bl[454] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_456 br[455] vdd vss bl[455] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_456 br[455] vdd vss bl[455] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_456 br[455] vdd vss bl[455] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_456 br[455] vdd vss bl[455] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_456 br[455] vdd vss bl[455] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_456 br[455] vdd vss bl[455] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_456 br[455] vdd vss bl[455] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_456 br[455] vdd vss bl[455] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_456 br[455] vdd vss bl[455] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_456 br[455] vdd vss bl[455] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_456 br[455] vdd vss bl[455] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_456 br[455] vdd vss bl[455] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_456 br[455] vdd vss bl[455] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_456 br[455] vdd vss bl[455] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_456 br[455] vdd vss bl[455] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_456 br[455] vdd vss bl[455] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_456 br[455] vdd vss bl[455] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_456 br[455] vdd vss bl[455] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_456 br[455] vdd vss bl[455] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_457 br[456] vdd vss bl[456] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_457 br[456] vdd vss bl[456] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_457 br[456] vdd vss bl[456] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_457 br[456] vdd vss bl[456] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_457 br[456] vdd vss bl[456] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_457 br[456] vdd vss bl[456] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_457 br[456] vdd vss bl[456] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_457 br[456] vdd vss bl[456] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_457 br[456] vdd vss bl[456] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_457 br[456] vdd vss bl[456] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_457 br[456] vdd vss bl[456] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_457 br[456] vdd vss bl[456] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_457 br[456] vdd vss bl[456] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_457 br[456] vdd vss bl[456] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_457 br[456] vdd vss bl[456] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_457 br[456] vdd vss bl[456] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_457 br[456] vdd vss bl[456] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_457 br[456] vdd vss bl[456] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_457 br[456] vdd vss bl[456] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_458 br[457] vdd vss bl[457] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_458 br[457] vdd vss bl[457] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_458 br[457] vdd vss bl[457] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_458 br[457] vdd vss bl[457] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_458 br[457] vdd vss bl[457] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_458 br[457] vdd vss bl[457] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_458 br[457] vdd vss bl[457] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_458 br[457] vdd vss bl[457] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_458 br[457] vdd vss bl[457] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_458 br[457] vdd vss bl[457] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_458 br[457] vdd vss bl[457] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_458 br[457] vdd vss bl[457] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_458 br[457] vdd vss bl[457] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_458 br[457] vdd vss bl[457] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_458 br[457] vdd vss bl[457] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_458 br[457] vdd vss bl[457] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_458 br[457] vdd vss bl[457] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_458 br[457] vdd vss bl[457] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_458 br[457] vdd vss bl[457] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_459 br[458] vdd vss bl[458] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_459 br[458] vdd vss bl[458] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_459 br[458] vdd vss bl[458] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_459 br[458] vdd vss bl[458] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_459 br[458] vdd vss bl[458] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_459 br[458] vdd vss bl[458] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_459 br[458] vdd vss bl[458] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_459 br[458] vdd vss bl[458] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_459 br[458] vdd vss bl[458] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_459 br[458] vdd vss bl[458] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_459 br[458] vdd vss bl[458] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_459 br[458] vdd vss bl[458] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_459 br[458] vdd vss bl[458] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_459 br[458] vdd vss bl[458] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_459 br[458] vdd vss bl[458] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_459 br[458] vdd vss bl[458] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_459 br[458] vdd vss bl[458] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_459 br[458] vdd vss bl[458] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_459 br[458] vdd vss bl[458] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_460 br[459] vdd vss bl[459] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_460 br[459] vdd vss bl[459] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_460 br[459] vdd vss bl[459] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_460 br[459] vdd vss bl[459] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_460 br[459] vdd vss bl[459] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_460 br[459] vdd vss bl[459] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_460 br[459] vdd vss bl[459] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_460 br[459] vdd vss bl[459] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_460 br[459] vdd vss bl[459] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_460 br[459] vdd vss bl[459] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_460 br[459] vdd vss bl[459] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_460 br[459] vdd vss bl[459] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_460 br[459] vdd vss bl[459] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_460 br[459] vdd vss bl[459] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_460 br[459] vdd vss bl[459] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_460 br[459] vdd vss bl[459] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_460 br[459] vdd vss bl[459] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_460 br[459] vdd vss bl[459] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_460 br[459] vdd vss bl[459] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_461 br[460] vdd vss bl[460] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_461 br[460] vdd vss bl[460] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_461 br[460] vdd vss bl[460] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_461 br[460] vdd vss bl[460] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_461 br[460] vdd vss bl[460] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_461 br[460] vdd vss bl[460] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_461 br[460] vdd vss bl[460] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_461 br[460] vdd vss bl[460] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_461 br[460] vdd vss bl[460] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_461 br[460] vdd vss bl[460] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_461 br[460] vdd vss bl[460] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_461 br[460] vdd vss bl[460] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_461 br[460] vdd vss bl[460] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_461 br[460] vdd vss bl[460] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_461 br[460] vdd vss bl[460] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_461 br[460] vdd vss bl[460] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_461 br[460] vdd vss bl[460] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_461 br[460] vdd vss bl[460] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_461 br[460] vdd vss bl[460] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_462 br[461] vdd vss bl[461] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_462 br[461] vdd vss bl[461] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_462 br[461] vdd vss bl[461] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_462 br[461] vdd vss bl[461] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_462 br[461] vdd vss bl[461] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_462 br[461] vdd vss bl[461] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_462 br[461] vdd vss bl[461] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_462 br[461] vdd vss bl[461] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_462 br[461] vdd vss bl[461] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_462 br[461] vdd vss bl[461] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_462 br[461] vdd vss bl[461] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_462 br[461] vdd vss bl[461] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_462 br[461] vdd vss bl[461] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_462 br[461] vdd vss bl[461] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_462 br[461] vdd vss bl[461] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_462 br[461] vdd vss bl[461] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_462 br[461] vdd vss bl[461] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_462 br[461] vdd vss bl[461] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_462 br[461] vdd vss bl[461] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_463 br[462] vdd vss bl[462] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_463 br[462] vdd vss bl[462] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_463 br[462] vdd vss bl[462] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_463 br[462] vdd vss bl[462] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_463 br[462] vdd vss bl[462] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_463 br[462] vdd vss bl[462] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_463 br[462] vdd vss bl[462] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_463 br[462] vdd vss bl[462] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_463 br[462] vdd vss bl[462] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_463 br[462] vdd vss bl[462] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_463 br[462] vdd vss bl[462] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_463 br[462] vdd vss bl[462] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_463 br[462] vdd vss bl[462] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_463 br[462] vdd vss bl[462] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_463 br[462] vdd vss bl[462] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_463 br[462] vdd vss bl[462] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_463 br[462] vdd vss bl[462] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_463 br[462] vdd vss bl[462] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_463 br[462] vdd vss bl[462] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_464 br[463] vdd vss bl[463] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_464 br[463] vdd vss bl[463] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_464 br[463] vdd vss bl[463] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_464 br[463] vdd vss bl[463] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_464 br[463] vdd vss bl[463] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_464 br[463] vdd vss bl[463] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_464 br[463] vdd vss bl[463] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_464 br[463] vdd vss bl[463] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_464 br[463] vdd vss bl[463] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_464 br[463] vdd vss bl[463] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_464 br[463] vdd vss bl[463] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_464 br[463] vdd vss bl[463] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_464 br[463] vdd vss bl[463] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_464 br[463] vdd vss bl[463] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_464 br[463] vdd vss bl[463] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_464 br[463] vdd vss bl[463] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_464 br[463] vdd vss bl[463] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_464 br[463] vdd vss bl[463] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_464 br[463] vdd vss bl[463] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_465 br[464] vdd vss bl[464] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_465 br[464] vdd vss bl[464] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_465 br[464] vdd vss bl[464] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_465 br[464] vdd vss bl[464] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_465 br[464] vdd vss bl[464] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_465 br[464] vdd vss bl[464] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_465 br[464] vdd vss bl[464] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_465 br[464] vdd vss bl[464] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_465 br[464] vdd vss bl[464] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_465 br[464] vdd vss bl[464] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_465 br[464] vdd vss bl[464] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_465 br[464] vdd vss bl[464] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_465 br[464] vdd vss bl[464] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_465 br[464] vdd vss bl[464] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_465 br[464] vdd vss bl[464] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_465 br[464] vdd vss bl[464] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_465 br[464] vdd vss bl[464] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_465 br[464] vdd vss bl[464] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_465 br[464] vdd vss bl[464] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_466 br[465] vdd vss bl[465] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_466 br[465] vdd vss bl[465] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_466 br[465] vdd vss bl[465] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_466 br[465] vdd vss bl[465] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_466 br[465] vdd vss bl[465] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_466 br[465] vdd vss bl[465] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_466 br[465] vdd vss bl[465] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_466 br[465] vdd vss bl[465] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_466 br[465] vdd vss bl[465] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_466 br[465] vdd vss bl[465] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_466 br[465] vdd vss bl[465] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_466 br[465] vdd vss bl[465] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_466 br[465] vdd vss bl[465] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_466 br[465] vdd vss bl[465] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_466 br[465] vdd vss bl[465] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_466 br[465] vdd vss bl[465] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_466 br[465] vdd vss bl[465] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_466 br[465] vdd vss bl[465] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_466 br[465] vdd vss bl[465] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_467 br[466] vdd vss bl[466] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_467 br[466] vdd vss bl[466] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_467 br[466] vdd vss bl[466] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_467 br[466] vdd vss bl[466] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_467 br[466] vdd vss bl[466] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_467 br[466] vdd vss bl[466] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_467 br[466] vdd vss bl[466] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_467 br[466] vdd vss bl[466] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_467 br[466] vdd vss bl[466] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_467 br[466] vdd vss bl[466] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_467 br[466] vdd vss bl[466] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_467 br[466] vdd vss bl[466] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_467 br[466] vdd vss bl[466] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_467 br[466] vdd vss bl[466] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_467 br[466] vdd vss bl[466] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_467 br[466] vdd vss bl[466] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_467 br[466] vdd vss bl[466] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_467 br[466] vdd vss bl[466] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_467 br[466] vdd vss bl[466] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_468 br[467] vdd vss bl[467] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_468 br[467] vdd vss bl[467] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_468 br[467] vdd vss bl[467] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_468 br[467] vdd vss bl[467] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_468 br[467] vdd vss bl[467] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_468 br[467] vdd vss bl[467] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_468 br[467] vdd vss bl[467] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_468 br[467] vdd vss bl[467] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_468 br[467] vdd vss bl[467] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_468 br[467] vdd vss bl[467] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_468 br[467] vdd vss bl[467] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_468 br[467] vdd vss bl[467] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_468 br[467] vdd vss bl[467] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_468 br[467] vdd vss bl[467] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_468 br[467] vdd vss bl[467] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_468 br[467] vdd vss bl[467] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_468 br[467] vdd vss bl[467] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_468 br[467] vdd vss bl[467] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_468 br[467] vdd vss bl[467] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_469 br[468] vdd vss bl[468] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_469 br[468] vdd vss bl[468] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_469 br[468] vdd vss bl[468] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_469 br[468] vdd vss bl[468] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_469 br[468] vdd vss bl[468] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_469 br[468] vdd vss bl[468] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_469 br[468] vdd vss bl[468] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_469 br[468] vdd vss bl[468] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_469 br[468] vdd vss bl[468] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_469 br[468] vdd vss bl[468] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_469 br[468] vdd vss bl[468] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_469 br[468] vdd vss bl[468] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_469 br[468] vdd vss bl[468] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_469 br[468] vdd vss bl[468] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_469 br[468] vdd vss bl[468] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_469 br[468] vdd vss bl[468] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_469 br[468] vdd vss bl[468] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_469 br[468] vdd vss bl[468] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_469 br[468] vdd vss bl[468] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_470 br[469] vdd vss bl[469] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_470 br[469] vdd vss bl[469] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_470 br[469] vdd vss bl[469] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_470 br[469] vdd vss bl[469] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_470 br[469] vdd vss bl[469] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_470 br[469] vdd vss bl[469] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_470 br[469] vdd vss bl[469] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_470 br[469] vdd vss bl[469] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_470 br[469] vdd vss bl[469] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_470 br[469] vdd vss bl[469] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_470 br[469] vdd vss bl[469] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_470 br[469] vdd vss bl[469] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_470 br[469] vdd vss bl[469] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_470 br[469] vdd vss bl[469] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_470 br[469] vdd vss bl[469] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_470 br[469] vdd vss bl[469] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_470 br[469] vdd vss bl[469] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_470 br[469] vdd vss bl[469] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_470 br[469] vdd vss bl[469] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_471 br[470] vdd vss bl[470] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_471 br[470] vdd vss bl[470] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_471 br[470] vdd vss bl[470] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_471 br[470] vdd vss bl[470] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_471 br[470] vdd vss bl[470] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_471 br[470] vdd vss bl[470] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_471 br[470] vdd vss bl[470] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_471 br[470] vdd vss bl[470] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_471 br[470] vdd vss bl[470] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_471 br[470] vdd vss bl[470] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_471 br[470] vdd vss bl[470] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_471 br[470] vdd vss bl[470] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_471 br[470] vdd vss bl[470] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_471 br[470] vdd vss bl[470] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_471 br[470] vdd vss bl[470] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_471 br[470] vdd vss bl[470] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_471 br[470] vdd vss bl[470] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_471 br[470] vdd vss bl[470] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_471 br[470] vdd vss bl[470] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_472 br[471] vdd vss bl[471] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_472 br[471] vdd vss bl[471] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_472 br[471] vdd vss bl[471] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_472 br[471] vdd vss bl[471] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_472 br[471] vdd vss bl[471] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_472 br[471] vdd vss bl[471] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_472 br[471] vdd vss bl[471] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_472 br[471] vdd vss bl[471] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_472 br[471] vdd vss bl[471] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_472 br[471] vdd vss bl[471] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_472 br[471] vdd vss bl[471] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_472 br[471] vdd vss bl[471] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_472 br[471] vdd vss bl[471] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_472 br[471] vdd vss bl[471] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_472 br[471] vdd vss bl[471] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_472 br[471] vdd vss bl[471] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_472 br[471] vdd vss bl[471] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_472 br[471] vdd vss bl[471] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_472 br[471] vdd vss bl[471] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_473 br[472] vdd vss bl[472] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_473 br[472] vdd vss bl[472] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_473 br[472] vdd vss bl[472] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_473 br[472] vdd vss bl[472] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_473 br[472] vdd vss bl[472] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_473 br[472] vdd vss bl[472] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_473 br[472] vdd vss bl[472] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_473 br[472] vdd vss bl[472] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_473 br[472] vdd vss bl[472] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_473 br[472] vdd vss bl[472] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_473 br[472] vdd vss bl[472] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_473 br[472] vdd vss bl[472] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_473 br[472] vdd vss bl[472] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_473 br[472] vdd vss bl[472] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_473 br[472] vdd vss bl[472] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_473 br[472] vdd vss bl[472] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_473 br[472] vdd vss bl[472] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_473 br[472] vdd vss bl[472] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_473 br[472] vdd vss bl[472] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_474 br[473] vdd vss bl[473] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_474 br[473] vdd vss bl[473] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_474 br[473] vdd vss bl[473] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_474 br[473] vdd vss bl[473] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_474 br[473] vdd vss bl[473] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_474 br[473] vdd vss bl[473] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_474 br[473] vdd vss bl[473] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_474 br[473] vdd vss bl[473] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_474 br[473] vdd vss bl[473] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_474 br[473] vdd vss bl[473] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_474 br[473] vdd vss bl[473] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_474 br[473] vdd vss bl[473] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_474 br[473] vdd vss bl[473] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_474 br[473] vdd vss bl[473] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_474 br[473] vdd vss bl[473] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_474 br[473] vdd vss bl[473] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_474 br[473] vdd vss bl[473] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_474 br[473] vdd vss bl[473] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_474 br[473] vdd vss bl[473] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_475 br[474] vdd vss bl[474] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_475 br[474] vdd vss bl[474] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_475 br[474] vdd vss bl[474] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_475 br[474] vdd vss bl[474] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_475 br[474] vdd vss bl[474] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_475 br[474] vdd vss bl[474] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_475 br[474] vdd vss bl[474] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_475 br[474] vdd vss bl[474] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_475 br[474] vdd vss bl[474] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_475 br[474] vdd vss bl[474] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_475 br[474] vdd vss bl[474] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_475 br[474] vdd vss bl[474] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_475 br[474] vdd vss bl[474] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_475 br[474] vdd vss bl[474] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_475 br[474] vdd vss bl[474] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_475 br[474] vdd vss bl[474] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_475 br[474] vdd vss bl[474] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_475 br[474] vdd vss bl[474] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_475 br[474] vdd vss bl[474] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_476 br[475] vdd vss bl[475] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_476 br[475] vdd vss bl[475] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_476 br[475] vdd vss bl[475] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_476 br[475] vdd vss bl[475] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_476 br[475] vdd vss bl[475] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_476 br[475] vdd vss bl[475] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_476 br[475] vdd vss bl[475] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_476 br[475] vdd vss bl[475] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_476 br[475] vdd vss bl[475] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_476 br[475] vdd vss bl[475] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_476 br[475] vdd vss bl[475] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_476 br[475] vdd vss bl[475] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_476 br[475] vdd vss bl[475] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_476 br[475] vdd vss bl[475] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_476 br[475] vdd vss bl[475] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_476 br[475] vdd vss bl[475] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_476 br[475] vdd vss bl[475] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_476 br[475] vdd vss bl[475] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_476 br[475] vdd vss bl[475] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_477 br[476] vdd vss bl[476] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_477 br[476] vdd vss bl[476] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_477 br[476] vdd vss bl[476] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_477 br[476] vdd vss bl[476] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_477 br[476] vdd vss bl[476] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_477 br[476] vdd vss bl[476] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_477 br[476] vdd vss bl[476] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_477 br[476] vdd vss bl[476] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_477 br[476] vdd vss bl[476] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_477 br[476] vdd vss bl[476] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_477 br[476] vdd vss bl[476] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_477 br[476] vdd vss bl[476] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_477 br[476] vdd vss bl[476] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_477 br[476] vdd vss bl[476] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_477 br[476] vdd vss bl[476] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_477 br[476] vdd vss bl[476] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_477 br[476] vdd vss bl[476] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_477 br[476] vdd vss bl[476] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_477 br[476] vdd vss bl[476] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_478 br[477] vdd vss bl[477] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_478 br[477] vdd vss bl[477] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_478 br[477] vdd vss bl[477] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_478 br[477] vdd vss bl[477] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_478 br[477] vdd vss bl[477] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_478 br[477] vdd vss bl[477] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_478 br[477] vdd vss bl[477] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_478 br[477] vdd vss bl[477] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_478 br[477] vdd vss bl[477] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_478 br[477] vdd vss bl[477] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_478 br[477] vdd vss bl[477] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_478 br[477] vdd vss bl[477] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_478 br[477] vdd vss bl[477] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_478 br[477] vdd vss bl[477] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_478 br[477] vdd vss bl[477] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_478 br[477] vdd vss bl[477] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_478 br[477] vdd vss bl[477] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_478 br[477] vdd vss bl[477] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_478 br[477] vdd vss bl[477] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_479 br[478] vdd vss bl[478] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_479 br[478] vdd vss bl[478] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_479 br[478] vdd vss bl[478] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_479 br[478] vdd vss bl[478] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_479 br[478] vdd vss bl[478] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_479 br[478] vdd vss bl[478] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_479 br[478] vdd vss bl[478] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_479 br[478] vdd vss bl[478] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_479 br[478] vdd vss bl[478] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_479 br[478] vdd vss bl[478] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_479 br[478] vdd vss bl[478] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_479 br[478] vdd vss bl[478] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_479 br[478] vdd vss bl[478] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_479 br[478] vdd vss bl[478] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_479 br[478] vdd vss bl[478] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_479 br[478] vdd vss bl[478] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_479 br[478] vdd vss bl[478] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_479 br[478] vdd vss bl[478] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_479 br[478] vdd vss bl[478] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_480 br[479] vdd vss bl[479] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_480 br[479] vdd vss bl[479] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_480 br[479] vdd vss bl[479] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_480 br[479] vdd vss bl[479] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_480 br[479] vdd vss bl[479] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_480 br[479] vdd vss bl[479] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_480 br[479] vdd vss bl[479] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_480 br[479] vdd vss bl[479] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_480 br[479] vdd vss bl[479] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_480 br[479] vdd vss bl[479] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_480 br[479] vdd vss bl[479] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_480 br[479] vdd vss bl[479] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_480 br[479] vdd vss bl[479] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_480 br[479] vdd vss bl[479] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_480 br[479] vdd vss bl[479] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_480 br[479] vdd vss bl[479] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_480 br[479] vdd vss bl[479] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_480 br[479] vdd vss bl[479] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_480 br[479] vdd vss bl[479] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_481 br[480] vdd vss bl[480] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_481 br[480] vdd vss bl[480] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_481 br[480] vdd vss bl[480] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_481 br[480] vdd vss bl[480] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_481 br[480] vdd vss bl[480] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_481 br[480] vdd vss bl[480] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_481 br[480] vdd vss bl[480] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_481 br[480] vdd vss bl[480] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_481 br[480] vdd vss bl[480] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_481 br[480] vdd vss bl[480] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_481 br[480] vdd vss bl[480] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_481 br[480] vdd vss bl[480] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_481 br[480] vdd vss bl[480] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_481 br[480] vdd vss bl[480] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_481 br[480] vdd vss bl[480] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_481 br[480] vdd vss bl[480] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_481 br[480] vdd vss bl[480] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_481 br[480] vdd vss bl[480] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_481 br[480] vdd vss bl[480] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_482 br[481] vdd vss bl[481] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_482 br[481] vdd vss bl[481] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_482 br[481] vdd vss bl[481] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_482 br[481] vdd vss bl[481] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_482 br[481] vdd vss bl[481] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_482 br[481] vdd vss bl[481] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_482 br[481] vdd vss bl[481] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_482 br[481] vdd vss bl[481] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_482 br[481] vdd vss bl[481] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_482 br[481] vdd vss bl[481] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_482 br[481] vdd vss bl[481] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_482 br[481] vdd vss bl[481] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_482 br[481] vdd vss bl[481] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_482 br[481] vdd vss bl[481] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_482 br[481] vdd vss bl[481] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_482 br[481] vdd vss bl[481] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_482 br[481] vdd vss bl[481] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_482 br[481] vdd vss bl[481] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_482 br[481] vdd vss bl[481] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_483 br[482] vdd vss bl[482] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_483 br[482] vdd vss bl[482] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_483 br[482] vdd vss bl[482] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_483 br[482] vdd vss bl[482] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_483 br[482] vdd vss bl[482] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_483 br[482] vdd vss bl[482] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_483 br[482] vdd vss bl[482] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_483 br[482] vdd vss bl[482] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_483 br[482] vdd vss bl[482] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_483 br[482] vdd vss bl[482] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_483 br[482] vdd vss bl[482] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_483 br[482] vdd vss bl[482] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_483 br[482] vdd vss bl[482] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_483 br[482] vdd vss bl[482] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_483 br[482] vdd vss bl[482] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_483 br[482] vdd vss bl[482] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_483 br[482] vdd vss bl[482] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_483 br[482] vdd vss bl[482] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_483 br[482] vdd vss bl[482] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_484 br[483] vdd vss bl[483] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_484 br[483] vdd vss bl[483] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_484 br[483] vdd vss bl[483] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_484 br[483] vdd vss bl[483] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_484 br[483] vdd vss bl[483] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_484 br[483] vdd vss bl[483] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_484 br[483] vdd vss bl[483] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_484 br[483] vdd vss bl[483] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_484 br[483] vdd vss bl[483] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_484 br[483] vdd vss bl[483] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_484 br[483] vdd vss bl[483] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_484 br[483] vdd vss bl[483] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_484 br[483] vdd vss bl[483] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_484 br[483] vdd vss bl[483] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_484 br[483] vdd vss bl[483] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_484 br[483] vdd vss bl[483] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_484 br[483] vdd vss bl[483] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_484 br[483] vdd vss bl[483] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_484 br[483] vdd vss bl[483] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_485 br[484] vdd vss bl[484] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_485 br[484] vdd vss bl[484] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_485 br[484] vdd vss bl[484] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_485 br[484] vdd vss bl[484] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_485 br[484] vdd vss bl[484] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_485 br[484] vdd vss bl[484] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_485 br[484] vdd vss bl[484] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_485 br[484] vdd vss bl[484] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_485 br[484] vdd vss bl[484] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_485 br[484] vdd vss bl[484] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_485 br[484] vdd vss bl[484] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_485 br[484] vdd vss bl[484] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_485 br[484] vdd vss bl[484] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_485 br[484] vdd vss bl[484] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_485 br[484] vdd vss bl[484] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_485 br[484] vdd vss bl[484] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_485 br[484] vdd vss bl[484] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_485 br[484] vdd vss bl[484] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_485 br[484] vdd vss bl[484] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_486 br[485] vdd vss bl[485] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_486 br[485] vdd vss bl[485] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_486 br[485] vdd vss bl[485] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_486 br[485] vdd vss bl[485] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_486 br[485] vdd vss bl[485] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_486 br[485] vdd vss bl[485] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_486 br[485] vdd vss bl[485] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_486 br[485] vdd vss bl[485] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_486 br[485] vdd vss bl[485] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_486 br[485] vdd vss bl[485] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_486 br[485] vdd vss bl[485] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_486 br[485] vdd vss bl[485] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_486 br[485] vdd vss bl[485] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_486 br[485] vdd vss bl[485] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_486 br[485] vdd vss bl[485] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_486 br[485] vdd vss bl[485] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_486 br[485] vdd vss bl[485] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_486 br[485] vdd vss bl[485] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_486 br[485] vdd vss bl[485] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_487 br[486] vdd vss bl[486] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_487 br[486] vdd vss bl[486] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_487 br[486] vdd vss bl[486] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_487 br[486] vdd vss bl[486] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_487 br[486] vdd vss bl[486] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_487 br[486] vdd vss bl[486] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_487 br[486] vdd vss bl[486] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_487 br[486] vdd vss bl[486] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_487 br[486] vdd vss bl[486] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_487 br[486] vdd vss bl[486] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_487 br[486] vdd vss bl[486] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_487 br[486] vdd vss bl[486] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_487 br[486] vdd vss bl[486] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_487 br[486] vdd vss bl[486] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_487 br[486] vdd vss bl[486] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_487 br[486] vdd vss bl[486] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_487 br[486] vdd vss bl[486] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_487 br[486] vdd vss bl[486] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_487 br[486] vdd vss bl[486] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_488 br[487] vdd vss bl[487] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_488 br[487] vdd vss bl[487] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_488 br[487] vdd vss bl[487] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_488 br[487] vdd vss bl[487] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_488 br[487] vdd vss bl[487] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_488 br[487] vdd vss bl[487] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_488 br[487] vdd vss bl[487] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_488 br[487] vdd vss bl[487] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_488 br[487] vdd vss bl[487] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_488 br[487] vdd vss bl[487] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_488 br[487] vdd vss bl[487] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_488 br[487] vdd vss bl[487] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_488 br[487] vdd vss bl[487] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_488 br[487] vdd vss bl[487] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_488 br[487] vdd vss bl[487] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_488 br[487] vdd vss bl[487] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_488 br[487] vdd vss bl[487] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_488 br[487] vdd vss bl[487] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_488 br[487] vdd vss bl[487] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_489 br[488] vdd vss bl[488] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_489 br[488] vdd vss bl[488] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_489 br[488] vdd vss bl[488] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_489 br[488] vdd vss bl[488] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_489 br[488] vdd vss bl[488] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_489 br[488] vdd vss bl[488] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_489 br[488] vdd vss bl[488] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_489 br[488] vdd vss bl[488] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_489 br[488] vdd vss bl[488] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_489 br[488] vdd vss bl[488] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_489 br[488] vdd vss bl[488] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_489 br[488] vdd vss bl[488] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_489 br[488] vdd vss bl[488] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_489 br[488] vdd vss bl[488] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_489 br[488] vdd vss bl[488] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_489 br[488] vdd vss bl[488] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_489 br[488] vdd vss bl[488] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_489 br[488] vdd vss bl[488] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_489 br[488] vdd vss bl[488] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_490 br[489] vdd vss bl[489] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_490 br[489] vdd vss bl[489] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_490 br[489] vdd vss bl[489] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_490 br[489] vdd vss bl[489] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_490 br[489] vdd vss bl[489] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_490 br[489] vdd vss bl[489] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_490 br[489] vdd vss bl[489] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_490 br[489] vdd vss bl[489] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_490 br[489] vdd vss bl[489] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_490 br[489] vdd vss bl[489] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_490 br[489] vdd vss bl[489] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_490 br[489] vdd vss bl[489] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_490 br[489] vdd vss bl[489] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_490 br[489] vdd vss bl[489] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_490 br[489] vdd vss bl[489] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_490 br[489] vdd vss bl[489] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_490 br[489] vdd vss bl[489] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_490 br[489] vdd vss bl[489] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_490 br[489] vdd vss bl[489] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_491 br[490] vdd vss bl[490] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_491 br[490] vdd vss bl[490] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_491 br[490] vdd vss bl[490] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_491 br[490] vdd vss bl[490] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_491 br[490] vdd vss bl[490] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_491 br[490] vdd vss bl[490] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_491 br[490] vdd vss bl[490] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_491 br[490] vdd vss bl[490] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_491 br[490] vdd vss bl[490] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_491 br[490] vdd vss bl[490] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_491 br[490] vdd vss bl[490] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_491 br[490] vdd vss bl[490] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_491 br[490] vdd vss bl[490] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_491 br[490] vdd vss bl[490] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_491 br[490] vdd vss bl[490] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_491 br[490] vdd vss bl[490] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_491 br[490] vdd vss bl[490] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_491 br[490] vdd vss bl[490] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_491 br[490] vdd vss bl[490] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_492 br[491] vdd vss bl[491] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_492 br[491] vdd vss bl[491] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_492 br[491] vdd vss bl[491] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_492 br[491] vdd vss bl[491] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_492 br[491] vdd vss bl[491] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_492 br[491] vdd vss bl[491] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_492 br[491] vdd vss bl[491] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_492 br[491] vdd vss bl[491] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_492 br[491] vdd vss bl[491] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_492 br[491] vdd vss bl[491] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_492 br[491] vdd vss bl[491] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_492 br[491] vdd vss bl[491] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_492 br[491] vdd vss bl[491] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_492 br[491] vdd vss bl[491] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_492 br[491] vdd vss bl[491] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_492 br[491] vdd vss bl[491] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_492 br[491] vdd vss bl[491] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_492 br[491] vdd vss bl[491] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_492 br[491] vdd vss bl[491] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_493 br[492] vdd vss bl[492] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_493 br[492] vdd vss bl[492] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_493 br[492] vdd vss bl[492] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_493 br[492] vdd vss bl[492] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_493 br[492] vdd vss bl[492] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_493 br[492] vdd vss bl[492] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_493 br[492] vdd vss bl[492] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_493 br[492] vdd vss bl[492] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_493 br[492] vdd vss bl[492] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_493 br[492] vdd vss bl[492] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_493 br[492] vdd vss bl[492] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_493 br[492] vdd vss bl[492] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_493 br[492] vdd vss bl[492] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_493 br[492] vdd vss bl[492] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_493 br[492] vdd vss bl[492] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_493 br[492] vdd vss bl[492] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_493 br[492] vdd vss bl[492] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_493 br[492] vdd vss bl[492] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_493 br[492] vdd vss bl[492] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_494 br[493] vdd vss bl[493] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_494 br[493] vdd vss bl[493] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_494 br[493] vdd vss bl[493] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_494 br[493] vdd vss bl[493] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_494 br[493] vdd vss bl[493] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_494 br[493] vdd vss bl[493] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_494 br[493] vdd vss bl[493] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_494 br[493] vdd vss bl[493] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_494 br[493] vdd vss bl[493] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_494 br[493] vdd vss bl[493] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_494 br[493] vdd vss bl[493] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_494 br[493] vdd vss bl[493] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_494 br[493] vdd vss bl[493] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_494 br[493] vdd vss bl[493] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_494 br[493] vdd vss bl[493] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_494 br[493] vdd vss bl[493] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_494 br[493] vdd vss bl[493] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_494 br[493] vdd vss bl[493] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_494 br[493] vdd vss bl[493] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_495 br[494] vdd vss bl[494] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_495 br[494] vdd vss bl[494] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_495 br[494] vdd vss bl[494] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_495 br[494] vdd vss bl[494] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_495 br[494] vdd vss bl[494] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_495 br[494] vdd vss bl[494] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_495 br[494] vdd vss bl[494] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_495 br[494] vdd vss bl[494] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_495 br[494] vdd vss bl[494] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_495 br[494] vdd vss bl[494] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_495 br[494] vdd vss bl[494] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_495 br[494] vdd vss bl[494] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_495 br[494] vdd vss bl[494] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_495 br[494] vdd vss bl[494] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_495 br[494] vdd vss bl[494] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_495 br[494] vdd vss bl[494] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_495 br[494] vdd vss bl[494] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_495 br[494] vdd vss bl[494] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_495 br[494] vdd vss bl[494] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_496 br[495] vdd vss bl[495] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_496 br[495] vdd vss bl[495] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_496 br[495] vdd vss bl[495] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_496 br[495] vdd vss bl[495] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_496 br[495] vdd vss bl[495] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_496 br[495] vdd vss bl[495] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_496 br[495] vdd vss bl[495] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_496 br[495] vdd vss bl[495] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_496 br[495] vdd vss bl[495] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_496 br[495] vdd vss bl[495] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_496 br[495] vdd vss bl[495] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_496 br[495] vdd vss bl[495] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_496 br[495] vdd vss bl[495] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_496 br[495] vdd vss bl[495] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_496 br[495] vdd vss bl[495] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_496 br[495] vdd vss bl[495] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_496 br[495] vdd vss bl[495] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_496 br[495] vdd vss bl[495] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_496 br[495] vdd vss bl[495] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_497 br[496] vdd vss bl[496] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_497 br[496] vdd vss bl[496] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_497 br[496] vdd vss bl[496] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_497 br[496] vdd vss bl[496] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_497 br[496] vdd vss bl[496] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_497 br[496] vdd vss bl[496] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_497 br[496] vdd vss bl[496] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_497 br[496] vdd vss bl[496] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_497 br[496] vdd vss bl[496] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_497 br[496] vdd vss bl[496] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_497 br[496] vdd vss bl[496] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_497 br[496] vdd vss bl[496] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_497 br[496] vdd vss bl[496] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_497 br[496] vdd vss bl[496] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_497 br[496] vdd vss bl[496] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_497 br[496] vdd vss bl[496] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_497 br[496] vdd vss bl[496] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_497 br[496] vdd vss bl[496] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_497 br[496] vdd vss bl[496] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_498 br[497] vdd vss bl[497] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_498 br[497] vdd vss bl[497] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_498 br[497] vdd vss bl[497] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_498 br[497] vdd vss bl[497] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_498 br[497] vdd vss bl[497] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_498 br[497] vdd vss bl[497] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_498 br[497] vdd vss bl[497] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_498 br[497] vdd vss bl[497] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_498 br[497] vdd vss bl[497] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_498 br[497] vdd vss bl[497] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_498 br[497] vdd vss bl[497] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_498 br[497] vdd vss bl[497] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_498 br[497] vdd vss bl[497] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_498 br[497] vdd vss bl[497] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_498 br[497] vdd vss bl[497] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_498 br[497] vdd vss bl[497] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_498 br[497] vdd vss bl[497] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_498 br[497] vdd vss bl[497] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_498 br[497] vdd vss bl[497] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_499 br[498] vdd vss bl[498] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_499 br[498] vdd vss bl[498] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_499 br[498] vdd vss bl[498] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_499 br[498] vdd vss bl[498] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_499 br[498] vdd vss bl[498] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_499 br[498] vdd vss bl[498] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_499 br[498] vdd vss bl[498] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_499 br[498] vdd vss bl[498] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_499 br[498] vdd vss bl[498] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_499 br[498] vdd vss bl[498] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_499 br[498] vdd vss bl[498] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_499 br[498] vdd vss bl[498] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_499 br[498] vdd vss bl[498] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_499 br[498] vdd vss bl[498] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_499 br[498] vdd vss bl[498] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_499 br[498] vdd vss bl[498] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_499 br[498] vdd vss bl[498] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_499 br[498] vdd vss bl[498] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_499 br[498] vdd vss bl[498] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_500 br[499] vdd vss bl[499] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_500 br[499] vdd vss bl[499] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_500 br[499] vdd vss bl[499] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_500 br[499] vdd vss bl[499] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_500 br[499] vdd vss bl[499] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_500 br[499] vdd vss bl[499] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_500 br[499] vdd vss bl[499] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_500 br[499] vdd vss bl[499] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_500 br[499] vdd vss bl[499] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_500 br[499] vdd vss bl[499] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_500 br[499] vdd vss bl[499] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_500 br[499] vdd vss bl[499] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_500 br[499] vdd vss bl[499] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_500 br[499] vdd vss bl[499] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_500 br[499] vdd vss bl[499] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_500 br[499] vdd vss bl[499] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_500 br[499] vdd vss bl[499] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_500 br[499] vdd vss bl[499] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_500 br[499] vdd vss bl[499] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_501 br[500] vdd vss bl[500] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_501 br[500] vdd vss bl[500] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_501 br[500] vdd vss bl[500] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_501 br[500] vdd vss bl[500] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_501 br[500] vdd vss bl[500] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_501 br[500] vdd vss bl[500] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_501 br[500] vdd vss bl[500] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_501 br[500] vdd vss bl[500] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_501 br[500] vdd vss bl[500] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_501 br[500] vdd vss bl[500] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_501 br[500] vdd vss bl[500] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_501 br[500] vdd vss bl[500] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_501 br[500] vdd vss bl[500] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_501 br[500] vdd vss bl[500] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_501 br[500] vdd vss bl[500] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_501 br[500] vdd vss bl[500] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_501 br[500] vdd vss bl[500] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_501 br[500] vdd vss bl[500] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_501 br[500] vdd vss bl[500] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_502 br[501] vdd vss bl[501] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_502 br[501] vdd vss bl[501] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_502 br[501] vdd vss bl[501] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_502 br[501] vdd vss bl[501] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_502 br[501] vdd vss bl[501] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_502 br[501] vdd vss bl[501] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_502 br[501] vdd vss bl[501] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_502 br[501] vdd vss bl[501] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_502 br[501] vdd vss bl[501] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_502 br[501] vdd vss bl[501] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_502 br[501] vdd vss bl[501] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_502 br[501] vdd vss bl[501] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_502 br[501] vdd vss bl[501] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_502 br[501] vdd vss bl[501] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_502 br[501] vdd vss bl[501] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_502 br[501] vdd vss bl[501] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_502 br[501] vdd vss bl[501] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_502 br[501] vdd vss bl[501] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_502 br[501] vdd vss bl[501] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_503 br[502] vdd vss bl[502] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_503 br[502] vdd vss bl[502] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_503 br[502] vdd vss bl[502] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_503 br[502] vdd vss bl[502] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_503 br[502] vdd vss bl[502] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_503 br[502] vdd vss bl[502] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_503 br[502] vdd vss bl[502] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_503 br[502] vdd vss bl[502] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_503 br[502] vdd vss bl[502] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_503 br[502] vdd vss bl[502] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_503 br[502] vdd vss bl[502] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_503 br[502] vdd vss bl[502] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_503 br[502] vdd vss bl[502] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_503 br[502] vdd vss bl[502] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_503 br[502] vdd vss bl[502] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_503 br[502] vdd vss bl[502] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_503 br[502] vdd vss bl[502] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_503 br[502] vdd vss bl[502] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_503 br[502] vdd vss bl[502] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_504 br[503] vdd vss bl[503] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_504 br[503] vdd vss bl[503] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_504 br[503] vdd vss bl[503] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_504 br[503] vdd vss bl[503] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_504 br[503] vdd vss bl[503] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_504 br[503] vdd vss bl[503] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_504 br[503] vdd vss bl[503] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_504 br[503] vdd vss bl[503] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_504 br[503] vdd vss bl[503] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_504 br[503] vdd vss bl[503] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_504 br[503] vdd vss bl[503] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_504 br[503] vdd vss bl[503] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_504 br[503] vdd vss bl[503] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_504 br[503] vdd vss bl[503] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_504 br[503] vdd vss bl[503] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_504 br[503] vdd vss bl[503] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_504 br[503] vdd vss bl[503] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_504 br[503] vdd vss bl[503] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_504 br[503] vdd vss bl[503] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_505 br[504] vdd vss bl[504] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_505 br[504] vdd vss bl[504] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_505 br[504] vdd vss bl[504] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_505 br[504] vdd vss bl[504] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_505 br[504] vdd vss bl[504] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_505 br[504] vdd vss bl[504] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_505 br[504] vdd vss bl[504] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_505 br[504] vdd vss bl[504] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_505 br[504] vdd vss bl[504] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_505 br[504] vdd vss bl[504] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_505 br[504] vdd vss bl[504] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_505 br[504] vdd vss bl[504] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_505 br[504] vdd vss bl[504] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_505 br[504] vdd vss bl[504] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_505 br[504] vdd vss bl[504] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_505 br[504] vdd vss bl[504] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_505 br[504] vdd vss bl[504] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_505 br[504] vdd vss bl[504] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_505 br[504] vdd vss bl[504] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_506 br[505] vdd vss bl[505] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_506 br[505] vdd vss bl[505] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_506 br[505] vdd vss bl[505] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_506 br[505] vdd vss bl[505] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_506 br[505] vdd vss bl[505] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_506 br[505] vdd vss bl[505] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_506 br[505] vdd vss bl[505] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_506 br[505] vdd vss bl[505] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_506 br[505] vdd vss bl[505] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_506 br[505] vdd vss bl[505] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_506 br[505] vdd vss bl[505] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_506 br[505] vdd vss bl[505] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_506 br[505] vdd vss bl[505] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_506 br[505] vdd vss bl[505] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_506 br[505] vdd vss bl[505] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_506 br[505] vdd vss bl[505] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_506 br[505] vdd vss bl[505] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_506 br[505] vdd vss bl[505] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_506 br[505] vdd vss bl[505] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_507 br[506] vdd vss bl[506] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_507 br[506] vdd vss bl[506] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_507 br[506] vdd vss bl[506] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_507 br[506] vdd vss bl[506] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_507 br[506] vdd vss bl[506] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_507 br[506] vdd vss bl[506] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_507 br[506] vdd vss bl[506] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_507 br[506] vdd vss bl[506] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_507 br[506] vdd vss bl[506] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_507 br[506] vdd vss bl[506] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_507 br[506] vdd vss bl[506] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_507 br[506] vdd vss bl[506] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_507 br[506] vdd vss bl[506] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_507 br[506] vdd vss bl[506] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_507 br[506] vdd vss bl[506] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_507 br[506] vdd vss bl[506] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_507 br[506] vdd vss bl[506] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_507 br[506] vdd vss bl[506] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_507 br[506] vdd vss bl[506] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_508 br[507] vdd vss bl[507] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_508 br[507] vdd vss bl[507] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_508 br[507] vdd vss bl[507] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_508 br[507] vdd vss bl[507] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_508 br[507] vdd vss bl[507] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_508 br[507] vdd vss bl[507] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_508 br[507] vdd vss bl[507] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_508 br[507] vdd vss bl[507] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_508 br[507] vdd vss bl[507] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_508 br[507] vdd vss bl[507] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_508 br[507] vdd vss bl[507] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_508 br[507] vdd vss bl[507] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_508 br[507] vdd vss bl[507] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_508 br[507] vdd vss bl[507] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_508 br[507] vdd vss bl[507] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_508 br[507] vdd vss bl[507] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_508 br[507] vdd vss bl[507] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_508 br[507] vdd vss bl[507] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_508 br[507] vdd vss bl[507] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_509 br[508] vdd vss bl[508] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_509 br[508] vdd vss bl[508] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_509 br[508] vdd vss bl[508] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_509 br[508] vdd vss bl[508] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_509 br[508] vdd vss bl[508] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_509 br[508] vdd vss bl[508] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_509 br[508] vdd vss bl[508] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_509 br[508] vdd vss bl[508] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_509 br[508] vdd vss bl[508] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_509 br[508] vdd vss bl[508] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_509 br[508] vdd vss bl[508] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_509 br[508] vdd vss bl[508] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_509 br[508] vdd vss bl[508] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_509 br[508] vdd vss bl[508] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_509 br[508] vdd vss bl[508] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_509 br[508] vdd vss bl[508] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_509 br[508] vdd vss bl[508] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_509 br[508] vdd vss bl[508] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_509 br[508] vdd vss bl[508] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_510 br[509] vdd vss bl[509] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_510 br[509] vdd vss bl[509] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_510 br[509] vdd vss bl[509] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_510 br[509] vdd vss bl[509] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_510 br[509] vdd vss bl[509] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_510 br[509] vdd vss bl[509] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_510 br[509] vdd vss bl[509] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_510 br[509] vdd vss bl[509] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_510 br[509] vdd vss bl[509] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_510 br[509] vdd vss bl[509] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_510 br[509] vdd vss bl[509] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_510 br[509] vdd vss bl[509] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_510 br[509] vdd vss bl[509] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_510 br[509] vdd vss bl[509] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_510 br[509] vdd vss bl[509] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_510 br[509] vdd vss bl[509] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_510 br[509] vdd vss bl[509] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_510 br[509] vdd vss bl[509] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_510 br[509] vdd vss bl[509] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_511 br[510] vdd vss bl[510] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_511 br[510] vdd vss bl[510] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_511 br[510] vdd vss bl[510] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_511 br[510] vdd vss bl[510] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_511 br[510] vdd vss bl[510] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_511 br[510] vdd vss bl[510] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_511 br[510] vdd vss bl[510] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_511 br[510] vdd vss bl[510] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_511 br[510] vdd vss bl[510] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_511 br[510] vdd vss bl[510] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_511 br[510] vdd vss bl[510] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_511 br[510] vdd vss bl[510] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_511 br[510] vdd vss bl[510] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_511 br[510] vdd vss bl[510] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_511 br[510] vdd vss bl[510] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_511 br[510] vdd vss bl[510] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_511 br[510] vdd vss bl[510] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_511 br[510] vdd vss bl[510] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_511 br[510] vdd vss bl[510] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_512 br[511] vdd vss bl[511] vss vdd sram_sp_colend_wrapper
  Xcolend_bot_512 br[511] vdd vss bl[511] vss vdd sram_sp_colend_wrapper
  Xhstrap_0_512 br[511] vdd vss bl[511] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_512 br[511] vdd vss bl[511] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_512 br[511] vdd vss bl[511] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_512 br[511] vdd vss bl[511] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_512 br[511] vdd vss bl[511] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_512 br[511] vdd vss bl[511] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_512 br[511] vdd vss bl[511] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_512 br[511] vdd vss bl[511] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_512 br[511] vdd vss bl[511] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_512 br[511] vdd vss bl[511] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_512 br[511] vdd vss bl[511] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_512 br[511] vdd vss bl[511] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_512 br[511] vdd vss bl[511] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_512 br[511] vdd vss bl[511] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_512 br[511] vdd vss bl[511] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_512 br[511] vdd vss bl[511] vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_512 br[511] vdd vss bl[511] vss vdd sram_sp_hstrap_wrapper
  Xcolend_top_513 vdd vdd vss vdd vss vdd sram_sp_colend_wrapper
  Xcolend_bot_513 vdd vdd vss vdd vss vdd sram_sp_colend_wrapper
  Xhstrap_0_513 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_513 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_513 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_513 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_4_513 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_5_513 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_6_513 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_7_513 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_8_513 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_9_513 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_10_513 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_11_513 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_12_513 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_13_513 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_14_513 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_15_513 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhstrap_16_513 vdd vdd vss vdd vss vdd sram_sp_hstrap_wrapper
  Xhoriz_wlstrap_0_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_0 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_1 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_2 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_3 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_4 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_5 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_6 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_7 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_8 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_9 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_9 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_9 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_9 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_9 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_9 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_9 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_9 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_9 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_9 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_9 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_9 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_9 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_9 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_9 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_9 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_9 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_10 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_10 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_10 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_10 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_10 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_10 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_10 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_10 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_10 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_10 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_10 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_10 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_10 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_10 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_10 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_10 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_10 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_11 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_11 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_11 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_11 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_11 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_11 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_11 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_11 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_11 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_11 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_11 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_11 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_11 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_11 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_11 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_11 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_11 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_12 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_12 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_12 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_12 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_12 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_12 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_12 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_12 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_12 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_12 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_12 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_12 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_12 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_12 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_12 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_12 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_12 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_13 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_13 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_13 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_13 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_13 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_13 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_13 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_13 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_13 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_13 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_13 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_13 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_13 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_13 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_13 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_13 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_13 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_14 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_14 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_14 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_14 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_14 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_14 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_14 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_14 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_14 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_14 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_14 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_14 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_14 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_14 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_14 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_14 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_14 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_15 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_15 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_15 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_15 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_15 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_15 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_15 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_15 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_15 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_15 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_15 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_15 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_15 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_15 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_15 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_15 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_15 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_16 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_16 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_16 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_16 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_16 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_16 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_16 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_16 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_16 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_16 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_16 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_16 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_16 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_16 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_16 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_16 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_16 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_17 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_17 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_17 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_17 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_17 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_17 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_17 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_17 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_17 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_17 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_17 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_17 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_17 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_17 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_17 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_17 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_17 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_18 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_18 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_18 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_18 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_18 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_18 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_18 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_18 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_18 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_18 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_18 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_18 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_18 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_18 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_18 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_18 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_18 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_19 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_19 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_19 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_19 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_19 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_19 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_19 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_19 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_19 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_19 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_19 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_19 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_19 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_19 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_19 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_19 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_19 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_20 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_20 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_20 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_20 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_20 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_20 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_20 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_20 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_20 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_20 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_20 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_20 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_20 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_20 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_20 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_20 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_20 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_21 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_21 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_21 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_21 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_21 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_21 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_21 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_21 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_21 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_21 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_21 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_21 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_21 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_21 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_21 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_21 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_21 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_22 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_22 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_22 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_22 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_22 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_22 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_22 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_22 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_22 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_22 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_22 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_22 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_22 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_22 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_22 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_22 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_22 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_23 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_23 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_23 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_23 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_23 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_23 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_23 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_23 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_23 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_23 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_23 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_23 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_23 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_23 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_23 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_23 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_23 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_24 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_24 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_24 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_24 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_24 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_24 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_24 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_24 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_24 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_24 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_24 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_24 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_24 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_24 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_24 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_24 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_24 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_25 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_25 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_25 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_25 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_25 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_25 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_25 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_25 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_25 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_25 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_25 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_25 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_25 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_25 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_25 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_25 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_25 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_26 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_26 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_26 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_26 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_26 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_26 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_26 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_26 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_26 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_26 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_26 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_26 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_26 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_26 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_26 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_26 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_26 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_27 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_27 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_27 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_27 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_27 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_27 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_27 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_27 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_27 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_27 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_27 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_27 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_27 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_27 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_27 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_27 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_27 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_28 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_28 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_28 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_28 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_28 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_28 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_28 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_28 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_28 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_28 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_28 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_28 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_28 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_28 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_28 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_28 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_28 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_29 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_29 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_29 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_29 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_29 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_29 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_29 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_29 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_29 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_29 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_29 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_29 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_29 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_29 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_29 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_29 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_29 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_30 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_30 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_30 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_30 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_30 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_30 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_30 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_30 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_30 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_30 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_30 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_30 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_30 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_30 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_30 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_30 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_30 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_31 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_31 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_31 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_31 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_31 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_31 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_31 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_31 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_31 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_31 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_31 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_31 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_31 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_31 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_31 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_31 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_31 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_32 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_32 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_32 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_32 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_32 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_32 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_32 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_32 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_32 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_32 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_32 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_32 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_32 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_32 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_32 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_32 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_32 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_33 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_33 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_33 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_33 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_33 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_33 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_33 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_33 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_33 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_33 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_33 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_33 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_33 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_33 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_33 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_33 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_33 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_34 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_34 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_34 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_34 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_34 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_34 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_34 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_34 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_34 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_34 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_34 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_34 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_34 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_34 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_34 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_34 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_34 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_35 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_35 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_35 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_35 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_35 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_35 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_35 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_35 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_35 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_35 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_35 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_35 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_35 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_35 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_35 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_35 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_35 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_36 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_36 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_36 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_36 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_36 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_36 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_36 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_36 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_36 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_36 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_36 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_36 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_36 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_36 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_36 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_36 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_36 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_37 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_37 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_37 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_37 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_37 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_37 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_37 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_37 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_37 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_37 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_37 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_37 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_37 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_37 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_37 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_37 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_37 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_38 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_38 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_38 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_38 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_38 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_38 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_38 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_38 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_38 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_38 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_38 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_38 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_38 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_38 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_38 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_38 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_38 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_39 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_39 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_39 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_39 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_39 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_39 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_39 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_39 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_39 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_39 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_39 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_39 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_39 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_39 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_39 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_39 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_39 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_40 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_40 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_40 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_40 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_40 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_40 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_40 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_40 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_40 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_40 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_40 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_40 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_40 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_40 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_40 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_40 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_40 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_41 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_41 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_41 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_41 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_41 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_41 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_41 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_41 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_41 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_41 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_41 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_41 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_41 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_41 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_41 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_41 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_41 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_42 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_42 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_42 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_42 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_42 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_42 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_42 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_42 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_42 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_42 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_42 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_42 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_42 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_42 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_42 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_42 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_42 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_43 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_43 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_43 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_43 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_43 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_43 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_43 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_43 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_43 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_43 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_43 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_43 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_43 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_43 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_43 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_43 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_43 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_44 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_44 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_44 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_44 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_44 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_44 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_44 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_44 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_44 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_44 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_44 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_44 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_44 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_44 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_44 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_44 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_44 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_45 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_45 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_45 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_45 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_45 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_45 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_45 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_45 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_45 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_45 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_45 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_45 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_45 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_45 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_45 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_45 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_45 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_46 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_46 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_46 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_46 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_46 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_46 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_46 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_46 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_46 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_46 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_46 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_46 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_46 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_46 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_46 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_46 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_46 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_47 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_47 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_47 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_47 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_47 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_47 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_47 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_47 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_47 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_47 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_47 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_47 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_47 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_47 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_47 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_47 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_47 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_48 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_48 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_48 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_48 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_48 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_48 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_48 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_48 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_48 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_48 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_48 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_48 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_48 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_48 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_48 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_48 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_48 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_49 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_49 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_49 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_49 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_49 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_49 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_49 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_49 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_49 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_49 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_49 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_49 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_49 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_49 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_49 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_49 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_49 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_50 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_50 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_50 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_50 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_50 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_50 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_50 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_50 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_50 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_50 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_50 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_50 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_50 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_50 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_50 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_50 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_50 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_51 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_51 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_51 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_51 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_51 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_51 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_51 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_51 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_51 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_51 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_51 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_51 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_51 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_51 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_51 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_51 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_51 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_52 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_52 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_52 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_52 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_52 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_52 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_52 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_52 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_52 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_52 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_52 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_52 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_52 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_52 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_52 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_52 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_52 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_53 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_53 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_53 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_53 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_53 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_53 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_53 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_53 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_53 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_53 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_53 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_53 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_53 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_53 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_53 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_53 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_53 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_54 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_54 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_54 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_54 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_54 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_54 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_54 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_54 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_54 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_54 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_54 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_54 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_54 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_54 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_54 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_54 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_54 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_55 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_55 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_55 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_55 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_55 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_55 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_55 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_55 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_55 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_55 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_55 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_55 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_55 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_55 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_55 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_55 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_55 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_56 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_56 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_56 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_56 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_56 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_56 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_56 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_56 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_56 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_56 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_56 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_56 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_56 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_56 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_56 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_56 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_56 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_57 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_57 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_57 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_57 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_57 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_57 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_57 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_57 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_57 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_57 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_57 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_57 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_57 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_57 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_57 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_57 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_57 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_58 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_58 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_58 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_58 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_58 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_58 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_58 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_58 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_58 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_58 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_58 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_58 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_58 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_58 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_58 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_58 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_58 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_59 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_59 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_59 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_59 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_59 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_59 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_59 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_59 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_59 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_59 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_59 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_59 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_59 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_59 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_59 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_59 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_59 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_60 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_60 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_60 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_60 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_60 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_60 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_60 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_60 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_60 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_60 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_60 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_60 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_60 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_60 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_60 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_60 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_60 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_61 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_61 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_61 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_61 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_61 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_61 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_61 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_61 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_61 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_61 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_61 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_61 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_61 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_61 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_61 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_61 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_61 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_62 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_62 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_62 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_62 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_62 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_62 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_62 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_62 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_62 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_62 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_62 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_62 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_62 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_62 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_62 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_62 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_62 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_63 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_63 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_63 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_63 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_63 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_63 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_63 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_63 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_63 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_63 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_63 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_63 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_63 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_63 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_63 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_63 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_63 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_64 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_64 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_64 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_64 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_64 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_64 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_64 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_64 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_64 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_64 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_64 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_64 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_64 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_64 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_64 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_64 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_64 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_65 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_65 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_65 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_65 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_65 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_65 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_65 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_65 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_65 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_65 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_65 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_65 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_65 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_65 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_65 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_65 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_65 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_66 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_66 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_66 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_66 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_66 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_66 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_66 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_66 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_66 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_66 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_66 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_66 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_66 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_66 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_66 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_66 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_66 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_67 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_67 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_67 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_67 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_67 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_67 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_67 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_67 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_67 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_67 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_67 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_67 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_67 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_67 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_67 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_67 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_67 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_68 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_68 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_68 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_68 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_68 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_68 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_68 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_68 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_68 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_68 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_68 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_68 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_68 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_68 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_68 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_68 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_68 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_69 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_69 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_69 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_69 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_69 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_69 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_69 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_69 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_69 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_69 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_69 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_69 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_69 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_69 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_69 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_69 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_69 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_70 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_70 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_70 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_70 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_70 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_70 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_70 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_70 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_70 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_70 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_70 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_70 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_70 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_70 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_70 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_70 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_70 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_71 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_71 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_71 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_71 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_71 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_71 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_71 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_71 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_71 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_71 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_71 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_71 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_71 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_71 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_71 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_71 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_71 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_72 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_72 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_72 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_72 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_72 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_72 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_72 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_72 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_72 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_72 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_72 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_72 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_72 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_72 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_72 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_72 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_72 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_73 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_73 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_73 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_73 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_73 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_73 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_73 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_73 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_73 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_73 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_73 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_73 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_73 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_73 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_73 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_73 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_73 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_74 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_74 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_74 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_74 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_74 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_74 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_74 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_74 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_74 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_74 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_74 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_74 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_74 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_74 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_74 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_74 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_74 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_75 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_75 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_75 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_75 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_75 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_75 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_75 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_75 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_75 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_75 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_75 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_75 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_75 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_75 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_75 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_75 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_75 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_76 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_76 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_76 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_76 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_76 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_76 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_76 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_76 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_76 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_76 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_76 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_76 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_76 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_76 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_76 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_76 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_76 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_77 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_77 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_77 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_77 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_77 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_77 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_77 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_77 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_77 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_77 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_77 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_77 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_77 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_77 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_77 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_77 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_77 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_78 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_78 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_78 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_78 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_78 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_78 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_78 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_78 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_78 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_78 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_78 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_78 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_78 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_78 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_78 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_78 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_78 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_79 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_79 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_79 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_79 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_79 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_79 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_79 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_79 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_79 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_79 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_79 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_79 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_79 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_79 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_79 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_79 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_79 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_80 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_80 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_80 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_80 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_80 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_80 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_80 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_80 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_80 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_80 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_80 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_80 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_80 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_80 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_80 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_80 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_80 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_81 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_81 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_81 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_81 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_81 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_81 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_81 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_81 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_81 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_81 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_81 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_81 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_81 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_81 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_81 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_81 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_81 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_82 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_82 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_82 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_82 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_82 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_82 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_82 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_82 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_82 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_82 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_82 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_82 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_82 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_82 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_82 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_82 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_82 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_83 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_83 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_83 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_83 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_83 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_83 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_83 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_83 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_83 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_83 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_83 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_83 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_83 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_83 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_83 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_83 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_83 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_84 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_84 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_84 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_84 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_84 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_84 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_84 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_84 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_84 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_84 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_84 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_84 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_84 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_84 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_84 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_84 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_84 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_85 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_85 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_85 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_85 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_85 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_85 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_85 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_85 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_85 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_85 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_85 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_85 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_85 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_85 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_85 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_85 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_85 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_86 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_86 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_86 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_86 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_86 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_86 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_86 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_86 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_86 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_86 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_86 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_86 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_86 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_86 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_86 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_86 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_86 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_87 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_87 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_87 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_87 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_87 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_87 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_87 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_87 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_87 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_87 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_87 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_87 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_87 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_87 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_87 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_87 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_87 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_88 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_88 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_88 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_88 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_88 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_88 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_88 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_88 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_88 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_88 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_88 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_88 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_88 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_88 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_88 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_88 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_88 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_89 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_89 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_89 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_89 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_89 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_89 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_89 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_89 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_89 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_89 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_89 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_89 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_89 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_89 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_89 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_89 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_89 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_90 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_90 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_90 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_90 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_90 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_90 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_90 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_90 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_90 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_90 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_90 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_90 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_90 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_90 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_90 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_90 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_90 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_91 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_91 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_91 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_91 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_91 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_91 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_91 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_91 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_91 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_91 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_91 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_91 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_91 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_91 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_91 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_91 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_91 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_92 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_92 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_92 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_92 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_92 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_92 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_92 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_92 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_92 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_92 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_92 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_92 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_92 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_92 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_92 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_92 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_92 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_93 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_93 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_93 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_93 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_93 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_93 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_93 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_93 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_93 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_93 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_93 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_93 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_93 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_93 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_93 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_93 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_93 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_94 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_94 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_94 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_94 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_94 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_94 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_94 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_94 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_94 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_94 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_94 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_94 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_94 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_94 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_94 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_94 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_94 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_95 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_95 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_95 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_95 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_95 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_95 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_95 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_95 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_95 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_95 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_95 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_95 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_95 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_95 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_95 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_95 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_95 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_96 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_96 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_96 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_96 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_96 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_96 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_96 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_96 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_96 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_96 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_96 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_96 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_96 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_96 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_96 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_96 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_96 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_97 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_97 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_97 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_97 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_97 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_97 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_97 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_97 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_97 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_97 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_97 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_97 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_97 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_97 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_97 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_97 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_97 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_98 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_98 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_98 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_98 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_98 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_98 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_98 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_98 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_98 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_98 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_98 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_98 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_98 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_98 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_98 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_98 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_98 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_99 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_99 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_99 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_99 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_99 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_99 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_99 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_99 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_99 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_99 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_99 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_99 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_99 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_99 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_99 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_99 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_99 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_100 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_100 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_100 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_100 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_100 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_100 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_100 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_100 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_100 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_100 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_100 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_100 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_100 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_100 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_100 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_100 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_100 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_101 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_101 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_101 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_101 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_101 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_101 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_101 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_101 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_101 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_101 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_101 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_101 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_101 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_101 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_101 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_101 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_101 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_102 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_102 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_102 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_102 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_102 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_102 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_102 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_102 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_102 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_102 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_102 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_102 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_102 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_102 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_102 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_102 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_102 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_103 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_103 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_103 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_103 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_103 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_103 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_103 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_103 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_103 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_103 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_103 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_103 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_103 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_103 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_103 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_103 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_103 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_104 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_104 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_104 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_104 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_104 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_104 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_104 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_104 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_104 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_104 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_104 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_104 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_104 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_104 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_104 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_104 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_104 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_105 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_105 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_105 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_105 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_105 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_105 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_105 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_105 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_105 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_105 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_105 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_105 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_105 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_105 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_105 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_105 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_105 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_106 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_106 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_106 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_106 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_106 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_106 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_106 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_106 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_106 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_106 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_106 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_106 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_106 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_106 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_106 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_106 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_106 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_107 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_107 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_107 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_107 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_107 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_107 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_107 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_107 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_107 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_107 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_107 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_107 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_107 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_107 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_107 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_107 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_107 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_108 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_108 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_108 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_108 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_108 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_108 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_108 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_108 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_108 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_108 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_108 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_108 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_108 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_108 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_108 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_108 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_108 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_109 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_109 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_109 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_109 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_109 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_109 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_109 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_109 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_109 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_109 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_109 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_109 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_109 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_109 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_109 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_109 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_109 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_110 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_110 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_110 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_110 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_110 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_110 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_110 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_110 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_110 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_110 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_110 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_110 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_110 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_110 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_110 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_110 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_110 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_111 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_111 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_111 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_111 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_111 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_111 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_111 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_111 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_111 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_111 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_111 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_111 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_111 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_111 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_111 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_111 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_111 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_112 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_112 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_112 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_112 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_112 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_112 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_112 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_112 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_112 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_112 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_112 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_112 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_112 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_112 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_112 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_112 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_112 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_113 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_113 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_113 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_113 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_113 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_113 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_113 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_113 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_113 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_113 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_113 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_113 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_113 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_113 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_113 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_113 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_113 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_114 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_114 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_114 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_114 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_114 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_114 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_114 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_114 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_114 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_114 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_114 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_114 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_114 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_114 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_114 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_114 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_114 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_115 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_115 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_115 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_115 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_115 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_115 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_115 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_115 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_115 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_115 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_115 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_115 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_115 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_115 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_115 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_115 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_115 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_116 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_116 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_116 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_116 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_116 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_116 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_116 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_116 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_116 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_116 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_116 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_116 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_116 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_116 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_116 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_116 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_116 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_117 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_117 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_117 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_117 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_117 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_117 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_117 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_117 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_117 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_117 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_117 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_117 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_117 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_117 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_117 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_117 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_117 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_118 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_118 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_118 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_118 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_118 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_118 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_118 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_118 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_118 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_118 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_118 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_118 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_118 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_118 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_118 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_118 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_118 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_119 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_119 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_119 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_119 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_119 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_119 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_119 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_119 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_119 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_119 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_119 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_119 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_119 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_119 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_119 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_119 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_119 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_120 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_120 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_120 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_120 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_120 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_120 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_120 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_120 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_120 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_120 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_120 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_120 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_120 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_120 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_120 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_120 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_120 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_121 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_121 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_121 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_121 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_121 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_121 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_121 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_121 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_121 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_121 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_121 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_121 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_121 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_121 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_121 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_121 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_121 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_122 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_122 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_122 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_122 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_122 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_122 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_122 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_122 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_122 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_122 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_122 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_122 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_122 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_122 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_122 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_122 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_122 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_123 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_123 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_123 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_123 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_123 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_123 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_123 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_123 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_123 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_123 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_123 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_123 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_123 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_123 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_123 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_123 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_123 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_124 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_124 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_124 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_124 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_124 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_124 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_124 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_124 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_124 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_124 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_124 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_124 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_124 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_124 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_124 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_124 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_124 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_125 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_125 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_125 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_125 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_125 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_125 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_125 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_125 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_125 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_125 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_125 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_125 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_125 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_125 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_125 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_125 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_125 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_126 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_126 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_126 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_126 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_126 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_126 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_126 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_126 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_126 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_126 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_126 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_126 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_126 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_126 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_126 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_126 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_126 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_127 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_127 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_127 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_127 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_127 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_127 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_127 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_127 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_127 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_127 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_127 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_127 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_127 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_127 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_127 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_127 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_127 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_0_128 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_1_128 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_2_128 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_3_128 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_4_128 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_5_128 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_6_128 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_7_128 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_8_128 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_9_128 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_10_128 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_11_128 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_12_128 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_13_128 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_14_128 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_15_128 vss vss sram_sp_horiz_wlstrap_p2_wrapper
  Xhoriz_wlstrap_16_128 vss vss sram_sp_horiz_wlstrap_p2_wrapper

.ENDS sp_cell_array

.SUBCKT sram_sp_cell_replica BL BR VSS VDD VPB VNB WL

  X0 VDD WL BR VNB sky130_fd_pr__special_nfet_pass l=0.150 nf=1 w=0.140

  X1 Q VDD VSS VNB sky130_fd_pr__special_nfet_latch l=0.150 nf=1 w=0.210

  X2 BL WL Q VNB sky130_fd_pr__special_nfet_pass l=0.150 nf=1 w=0.140

  X3 Q WL Q VPB sky130_fd_pr__special_pfet_pass l=0.025 nf=1 w=0.140

  X4 VDD WL VDD VPB sky130_fd_pr__special_pfet_pass l=0.025 nf=1 w=0.140

  X5 VDD Q VDD VPB sky130_fd_pr__special_pfet_pass l=0.150 nf=1 w=0.140

  X6 Q VDD VDD VPB sky130_fd_pr__special_pfet_pass l=0.150 nf=1 w=0.140

  X7 VSS Q VDD VNB sky130_fd_pr__special_nfet_latch l=0.150 nf=1 w=0.210


.ENDS sram_sp_cell_replica

.SUBCKT sram_sp_cell_replica_wrapper BL BR VSS VDD VPB VNB WL

  X0 BL BR VSS VDD VPB VNB WL sram_sp_cell_replica

.ENDS sram_sp_cell_replica_wrapper

.SUBCKT sram_sp_rowtapend_replica VSS VNB

  X0 VSS VSS VSS VNB sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.420


.ENDS sram_sp_rowtapend_replica

.SUBCKT sram_sp_rowtapend_replica_wrapper VSS VNB

  X0 VSS VNB sram_sp_rowtapend_replica

.ENDS sram_sp_rowtapend_replica_wrapper

.SUBCKT replica_cell_array vdd vss rbl rbr rwl

  Xcell_0_0 rbl rbr vss vdd vdd vss rwl sram_sp_cell_replica_wrapper
  Xcell_0_1 rbl rbr vss vdd vdd vss rwl sram_sp_cell_replica_wrapper
  Xcell_1_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_1_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_2_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_2_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_3_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_3_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_4_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_4_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_5_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_5_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_6_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_6_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_7_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_7_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_8_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_8_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_9_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_9_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_10_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_10_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_11_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_11_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_12_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_12_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_13_0 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcell_13_1 rbl rbr vss vdd vdd vss vss sram_sp_cell_replica_wrapper
  Xcolend_0_0 rbr vdd vss rbl vss vdd sram_sp_colend_wrapper
  Xcolend_1_0 rbr vdd vss rbl vss vdd sram_sp_colend_wrapper
  Xcolend_0_1 rbr vdd vss rbl vss vdd sram_sp_colend_wrapper
  Xcolend_1_1 rbr vdd vss rbl vss vdd sram_sp_colend_wrapper
  Xrowtapend_0_0 vss vss sram_sp_rowtapend_replica_wrapper
  Xrowtapend_0_1 vss vss sram_sp_rowtapend_replica_wrapper
  Xhstrap_0_0 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_0_1 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xrowtapend_1_0 vss vss sram_sp_rowtapend_replica_wrapper
  Xrowtapend_1_1 vss vss sram_sp_rowtapend_replica_wrapper
  Xhstrap_1_0 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_1_1 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xrowtapend_2_0 vss vss sram_sp_rowtapend_replica_wrapper
  Xrowtapend_2_1 vss vss sram_sp_rowtapend_replica_wrapper
  Xhstrap_2_0 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_2_1 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xrowtapend_3_0 vss vss sram_sp_rowtapend_replica_wrapper
  Xrowtapend_3_1 vss vss sram_sp_rowtapend_replica_wrapper
  Xhstrap_3_0 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper
  Xhstrap_3_1 rbr vdd vss rbl vss vdd sram_sp_hstrap_wrapper

.ENDS replica_cell_array

.SUBCKT dff_array_16 vdd vss clk rb d[0] d[1] d[2] d[3] d[4] d[5] d[6] d[7] d[8] d[9] d[10] d[11] d[12] d[13] d[14] d[15] q[0] q[1] q[2] q[3] q[4] q[5] q[6] q[7] q[8] q[9] q[10] q[11] q[12] q[13] q[14] q[15] qn[0] qn[1] qn[2] qn[3] qn[4] qn[5] qn[6] qn[7] qn[8] qn[9] qn[10] qn[11] qn[12] qn[13] qn[14] qn[15]

  Xdff_0 clk d[0] rb vss vss vdd vdd q[0] qn[0] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_1 clk d[1] rb vss vss vdd vdd q[1] qn[1] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_2 clk d[2] rb vss vss vdd vdd q[2] qn[2] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_3 clk d[3] rb vss vss vdd vdd q[3] qn[3] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_4 clk d[4] rb vss vss vdd vdd q[4] qn[4] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_5 clk d[5] rb vss vss vdd vdd q[5] qn[5] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_6 clk d[6] rb vss vss vdd vdd q[6] qn[6] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_7 clk d[7] rb vss vss vdd vdd q[7] qn[7] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_8 clk d[8] rb vss vss vdd vdd q[8] qn[8] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_9 clk d[9] rb vss vss vdd vdd q[9] qn[9] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_10 clk d[10] rb vss vss vdd vdd q[10] qn[10] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_11 clk d[11] rb vss vss vdd vdd q[11] qn[11] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_12 clk d[12] rb vss vss vdd vdd q[12] qn[12] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_13 clk d[13] rb vss vss vdd vdd q[13] qn[13] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_14 clk d[14] rb vss vss vdd vdd q[14] qn[14] sky130_fd_sc_hs__dfrbp_2_wrapper
  Xdff_15 clk d[15] rb vss vss vdd vdd q[15] qn[15] sky130_fd_sc_hs__dfrbp_2_wrapper

.ENDS dff_array_16

.SUBCKT mos_w1300_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=1.300


.ENDS mos_w1300_l150_m1_nf1_id0

.SUBCKT folded_inv_2 vdd vss a y

  XMP0 y a vdd vdd mos_w3230_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w1300_l150_m1_nf1_id0
  XMP1 y a vdd vdd mos_w3230_l150_m1_nf1_id1
  XMN1 y a vss vss mos_w1300_l150_m1_nf1_id0

.ENDS folded_inv_2

.SUBCKT mos_w2890_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=2.890


.ENDS mos_w2890_l150_m1_nf1_id1

.SUBCKT mos_w1160_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=1.160


.ENDS mos_w1160_l150_m1_nf1_id0

.SUBCKT folded_inv_3 vdd vss a y

  XMP0 y a vdd vdd mos_w2890_l150_m1_nf1_id1
  XMN0 y a vss vss mos_w1160_l150_m1_nf1_id0
  XMP1 y a vdd vdd mos_w2890_l150_m1_nf1_id1
  XMN1 y a vss vss mos_w1160_l150_m1_nf1_id0

.ENDS folded_inv_3

.SUBCKT decoder_stage_7 vdd vss y y_b predecode_0_0 predecode_1_0

  Xgate_0_0_0 vdd vss predecode_0_0 predecode_1_0 x_0 nand2_1
  Xgate_1_0_0 vdd vss x_0 x_1 folded_inv_2
  Xgate_2_0_0 vdd vss x_1 y_b folded_inv_3
  Xgate_2_0_1 vdd vss x_1 y_b folded_inv_3
  Xgate_2_0_2 vdd vss x_1 y_b folded_inv_3
  Xgate_3_0_0 vdd vss y_b y folded_inv_3
  Xgate_3_0_1 vdd vss y_b y folded_inv_3
  Xgate_3_0_2 vdd vss y_b y folded_inv_3

.ENDS decoder_stage_7

.SUBCKT mos_w2600_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=2.600


.ENDS mos_w2600_l150_m1_nf1_id1

.SUBCKT mos_w1550_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.550


.ENDS mos_w1550_l150_m1_nf1_id1

.SUBCKT precharge_1 vdd bl br en_b

  Xbl_pull_up bl en_b vdd vdd mos_w2600_l150_m1_nf1_id1
  Xbr_pull_up br en_b vdd vdd mos_w2600_l150_m1_nf1_id1
  Xequalizer bl en_b br vdd mos_w1550_l150_m1_nf1_id1

.ENDS precharge_1

.SUBCKT mos_w3650_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=3.650


.ENDS mos_w3650_l150_m1_nf1_id1

.SUBCKT mos_w2400_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=2.400


.ENDS mos_w2400_l150_m1_nf1_id0

.SUBCKT tgate_mux sel_b sel bl br bl_out br_out vdd vss

  XMPBL bl_out sel_b bl vdd mos_w3650_l150_m1_nf1_id1
  XMPBR br_out sel_b br vdd mos_w3650_l150_m1_nf1_id1
  XMNBL bl_out sel bl vss mos_w2400_l150_m1_nf1_id0
  XMNBR br_out sel br vss mos_w2400_l150_m1_nf1_id0

.ENDS tgate_mux

.SUBCKT mos_w2600_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=2.600


.ENDS mos_w2600_l150_m1_nf1_id0

.SUBCKT tristate_inv din en en_b din_b vdd vss

  Xmn_en din_b en nint vss mos_w2600_l150_m1_nf1_id0
  Xmn_pd nint din vss vss mos_w2600_l150_m1_nf1_id0
  Xmp_en din_b en_b pint vdd mos_w2600_l150_m1_nf1_id1
  Xmp_pu pint din vdd vdd mos_w2600_l150_m1_nf1_id1

.ENDS tristate_inv

.SUBCKT write_driver en en_b data data_b bl br vdd vss

  Xbldriver data_b en en_b bl vdd vss tristate_inv
  Xbrdriver data en en_b br vdd vss tristate_inv

.ENDS write_driver

.SUBCKT sramgen_sp_sense_amp clk inn inp outn outp VDD VSS

  XSWOP outp clk VDD VDD sky130_fd_pr__pfet_01v8 l=0.150 nf=2 w=1.000

  XSWON outn clk VDD VDD sky130_fd_pr__pfet_01v8 l=0.150 nf=2 w=1.000

  XSWMP midp clk VDD VDD sky130_fd_pr__pfet_01v8 l=0.150 nf=2 w=1.000

  XSWMN midn clk VDD VDD sky130_fd_pr__pfet_01v8 l=0.150 nf=2 w=1.000

  XPFBP outp outn VDD VDD sky130_fd_pr__pfet_01v8 l=0.150 nf=2 w=2.000

  XPFBN outn outp VDD VDD sky130_fd_pr__pfet_01v8 l=0.150 nf=2 w=2.000

  XTAIL tail clk VSS VSS sky130_fd_pr__nfet_01v8 l=0.150 nf=4 w=1.680

  XNFBP outp outn midp VSS sky130_fd_pr__nfet_01v8 l=0.150 nf=2 w=1.680

  XNFBN outn outp midn VSS sky130_fd_pr__nfet_01v8 l=0.150 nf=2 w=1.680

  XINP midn inp tail VSS sky130_fd_pr__nfet_01v8 l=0.150 nf=2 w=1.680

  XINN midp inn tail VSS sky130_fd_pr__nfet_01v8 l=0.150 nf=2 w=1.680


.ENDS sramgen_sp_sense_amp

.SUBCKT sramgen_sp_sense_amp_wrapper clk inn inp outn outp VDD VSS

  X0 clk inn inp outn outp VDD VSS sramgen_sp_sense_amp

.ENDS sramgen_sp_sense_amp_wrapper

.SUBCKT column clk rstb vdd vss bl[0] bl[1] bl[2] bl[3] br[0] br[1] br[2] br[3] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we we_b din dout sense_en

  Xprecharge_0 vdd bl[0] br[0] pc_b precharge_1
  Xmux_0 sel_b[0] sel[0] bl[0] br[0] bl_out br_out vdd vss tgate_mux
  Xprecharge_1 vdd bl[1] br[1] pc_b precharge_1
  Xmux_1 sel_b[1] sel[1] bl[1] br[1] bl_out br_out vdd vss tgate_mux
  Xprecharge_2 vdd bl[2] br[2] pc_b precharge_1
  Xmux_2 sel_b[2] sel[2] bl[2] br[2] bl_out br_out vdd vss tgate_mux
  Xprecharge_3 vdd bl[3] br[3] pc_b precharge_1
  Xmux_3 sel_b[3] sel[3] bl[3] br[3] bl_out br_out vdd vss tgate_mux
  Xwrite_driver we we_b q q_b bl_out br_out vdd vss write_driver
  Xsense_amp sense_en br_out bl_out sa_outn sa_outp vdd vss sramgen_sp_sense_amp_wrapper
  Xlatch vdd vss sa_outp sa_outn dout diff_latch_outn diff_latch
  Xdff clk din rstb vss vss vdd vdd q q_b sky130_fd_sc_hs__dfrbp_2_wrapper

.ENDS column

.SUBCKT col_peripherals clk rstb vdd vss sense_en bl[0] bl[1] bl[2] bl[3] bl[4] bl[5] bl[6] bl[7] bl[8] bl[9] bl[10] bl[11] bl[12] bl[13] bl[14] bl[15] bl[16] bl[17] bl[18] bl[19] bl[20] bl[21] bl[22] bl[23] bl[24] bl[25] bl[26] bl[27] bl[28] bl[29] bl[30] bl[31] bl[32] bl[33] bl[34] bl[35] bl[36] bl[37] bl[38] bl[39] bl[40] bl[41] bl[42] bl[43] bl[44] bl[45] bl[46] bl[47] bl[48] bl[49] bl[50] bl[51] bl[52] bl[53] bl[54] bl[55] bl[56] bl[57] bl[58] bl[59] bl[60] bl[61] bl[62] bl[63] bl[64] bl[65] bl[66] bl[67] bl[68] bl[69] bl[70] bl[71] bl[72] bl[73] bl[74] bl[75] bl[76] bl[77] bl[78] bl[79] bl[80] bl[81] bl[82] bl[83] bl[84] bl[85] bl[86] bl[87] bl[88] bl[89] bl[90] bl[91] bl[92] bl[93] bl[94] bl[95] bl[96] bl[97] bl[98] bl[99] bl[100] bl[101] bl[102] bl[103] bl[104] bl[105] bl[106] bl[107] bl[108] bl[109] bl[110] bl[111] bl[112] bl[113] bl[114] bl[115] bl[116] bl[117] bl[118] bl[119] bl[120] bl[121] bl[122] bl[123] bl[124] bl[125] bl[126] bl[127] bl[128] bl[129] bl[130] bl[131] bl[132] bl[133] bl[134] bl[135] bl[136] bl[137] bl[138] bl[139] bl[140] bl[141] bl[142] bl[143] bl[144] bl[145] bl[146] bl[147] bl[148] bl[149] bl[150] bl[151] bl[152] bl[153] bl[154] bl[155] bl[156] bl[157] bl[158] bl[159] bl[160] bl[161] bl[162] bl[163] bl[164] bl[165] bl[166] bl[167] bl[168] bl[169] bl[170] bl[171] bl[172] bl[173] bl[174] bl[175] bl[176] bl[177] bl[178] bl[179] bl[180] bl[181] bl[182] bl[183] bl[184] bl[185] bl[186] bl[187] bl[188] bl[189] bl[190] bl[191] bl[192] bl[193] bl[194] bl[195] bl[196] bl[197] bl[198] bl[199] bl[200] bl[201] bl[202] bl[203] bl[204] bl[205] bl[206] bl[207] bl[208] bl[209] bl[210] bl[211] bl[212] bl[213] bl[214] bl[215] bl[216] bl[217] bl[218] bl[219] bl[220] bl[221] bl[222] bl[223] bl[224] bl[225] bl[226] bl[227] bl[228] bl[229] bl[230] bl[231] bl[232] bl[233] bl[234] bl[235] bl[236] bl[237] bl[238] bl[239] bl[240] bl[241] bl[242] bl[243] bl[244] bl[245] bl[246] bl[247] bl[248] bl[249] bl[250] bl[251] bl[252] bl[253] bl[254] bl[255] bl[256] bl[257] bl[258] bl[259] bl[260] bl[261] bl[262] bl[263] bl[264] bl[265] bl[266] bl[267] bl[268] bl[269] bl[270] bl[271] bl[272] bl[273] bl[274] bl[275] bl[276] bl[277] bl[278] bl[279] bl[280] bl[281] bl[282] bl[283] bl[284] bl[285] bl[286] bl[287] bl[288] bl[289] bl[290] bl[291] bl[292] bl[293] bl[294] bl[295] bl[296] bl[297] bl[298] bl[299] bl[300] bl[301] bl[302] bl[303] bl[304] bl[305] bl[306] bl[307] bl[308] bl[309] bl[310] bl[311] bl[312] bl[313] bl[314] bl[315] bl[316] bl[317] bl[318] bl[319] bl[320] bl[321] bl[322] bl[323] bl[324] bl[325] bl[326] bl[327] bl[328] bl[329] bl[330] bl[331] bl[332] bl[333] bl[334] bl[335] bl[336] bl[337] bl[338] bl[339] bl[340] bl[341] bl[342] bl[343] bl[344] bl[345] bl[346] bl[347] bl[348] bl[349] bl[350] bl[351] bl[352] bl[353] bl[354] bl[355] bl[356] bl[357] bl[358] bl[359] bl[360] bl[361] bl[362] bl[363] bl[364] bl[365] bl[366] bl[367] bl[368] bl[369] bl[370] bl[371] bl[372] bl[373] bl[374] bl[375] bl[376] bl[377] bl[378] bl[379] bl[380] bl[381] bl[382] bl[383] bl[384] bl[385] bl[386] bl[387] bl[388] bl[389] bl[390] bl[391] bl[392] bl[393] bl[394] bl[395] bl[396] bl[397] bl[398] bl[399] bl[400] bl[401] bl[402] bl[403] bl[404] bl[405] bl[406] bl[407] bl[408] bl[409] bl[410] bl[411] bl[412] bl[413] bl[414] bl[415] bl[416] bl[417] bl[418] bl[419] bl[420] bl[421] bl[422] bl[423] bl[424] bl[425] bl[426] bl[427] bl[428] bl[429] bl[430] bl[431] bl[432] bl[433] bl[434] bl[435] bl[436] bl[437] bl[438] bl[439] bl[440] bl[441] bl[442] bl[443] bl[444] bl[445] bl[446] bl[447] bl[448] bl[449] bl[450] bl[451] bl[452] bl[453] bl[454] bl[455] bl[456] bl[457] bl[458] bl[459] bl[460] bl[461] bl[462] bl[463] bl[464] bl[465] bl[466] bl[467] bl[468] bl[469] bl[470] bl[471] bl[472] bl[473] bl[474] bl[475] bl[476] bl[477] bl[478] bl[479] bl[480] bl[481] bl[482] bl[483] bl[484] bl[485] bl[486] bl[487] bl[488] bl[489] bl[490] bl[491] bl[492] bl[493] bl[494] bl[495] bl[496] bl[497] bl[498] bl[499] bl[500] bl[501] bl[502] bl[503] bl[504] bl[505] bl[506] bl[507] bl[508] bl[509] bl[510] bl[511] br[0] br[1] br[2] br[3] br[4] br[5] br[6] br[7] br[8] br[9] br[10] br[11] br[12] br[13] br[14] br[15] br[16] br[17] br[18] br[19] br[20] br[21] br[22] br[23] br[24] br[25] br[26] br[27] br[28] br[29] br[30] br[31] br[32] br[33] br[34] br[35] br[36] br[37] br[38] br[39] br[40] br[41] br[42] br[43] br[44] br[45] br[46] br[47] br[48] br[49] br[50] br[51] br[52] br[53] br[54] br[55] br[56] br[57] br[58] br[59] br[60] br[61] br[62] br[63] br[64] br[65] br[66] br[67] br[68] br[69] br[70] br[71] br[72] br[73] br[74] br[75] br[76] br[77] br[78] br[79] br[80] br[81] br[82] br[83] br[84] br[85] br[86] br[87] br[88] br[89] br[90] br[91] br[92] br[93] br[94] br[95] br[96] br[97] br[98] br[99] br[100] br[101] br[102] br[103] br[104] br[105] br[106] br[107] br[108] br[109] br[110] br[111] br[112] br[113] br[114] br[115] br[116] br[117] br[118] br[119] br[120] br[121] br[122] br[123] br[124] br[125] br[126] br[127] br[128] br[129] br[130] br[131] br[132] br[133] br[134] br[135] br[136] br[137] br[138] br[139] br[140] br[141] br[142] br[143] br[144] br[145] br[146] br[147] br[148] br[149] br[150] br[151] br[152] br[153] br[154] br[155] br[156] br[157] br[158] br[159] br[160] br[161] br[162] br[163] br[164] br[165] br[166] br[167] br[168] br[169] br[170] br[171] br[172] br[173] br[174] br[175] br[176] br[177] br[178] br[179] br[180] br[181] br[182] br[183] br[184] br[185] br[186] br[187] br[188] br[189] br[190] br[191] br[192] br[193] br[194] br[195] br[196] br[197] br[198] br[199] br[200] br[201] br[202] br[203] br[204] br[205] br[206] br[207] br[208] br[209] br[210] br[211] br[212] br[213] br[214] br[215] br[216] br[217] br[218] br[219] br[220] br[221] br[222] br[223] br[224] br[225] br[226] br[227] br[228] br[229] br[230] br[231] br[232] br[233] br[234] br[235] br[236] br[237] br[238] br[239] br[240] br[241] br[242] br[243] br[244] br[245] br[246] br[247] br[248] br[249] br[250] br[251] br[252] br[253] br[254] br[255] br[256] br[257] br[258] br[259] br[260] br[261] br[262] br[263] br[264] br[265] br[266] br[267] br[268] br[269] br[270] br[271] br[272] br[273] br[274] br[275] br[276] br[277] br[278] br[279] br[280] br[281] br[282] br[283] br[284] br[285] br[286] br[287] br[288] br[289] br[290] br[291] br[292] br[293] br[294] br[295] br[296] br[297] br[298] br[299] br[300] br[301] br[302] br[303] br[304] br[305] br[306] br[307] br[308] br[309] br[310] br[311] br[312] br[313] br[314] br[315] br[316] br[317] br[318] br[319] br[320] br[321] br[322] br[323] br[324] br[325] br[326] br[327] br[328] br[329] br[330] br[331] br[332] br[333] br[334] br[335] br[336] br[337] br[338] br[339] br[340] br[341] br[342] br[343] br[344] br[345] br[346] br[347] br[348] br[349] br[350] br[351] br[352] br[353] br[354] br[355] br[356] br[357] br[358] br[359] br[360] br[361] br[362] br[363] br[364] br[365] br[366] br[367] br[368] br[369] br[370] br[371] br[372] br[373] br[374] br[375] br[376] br[377] br[378] br[379] br[380] br[381] br[382] br[383] br[384] br[385] br[386] br[387] br[388] br[389] br[390] br[391] br[392] br[393] br[394] br[395] br[396] br[397] br[398] br[399] br[400] br[401] br[402] br[403] br[404] br[405] br[406] br[407] br[408] br[409] br[410] br[411] br[412] br[413] br[414] br[415] br[416] br[417] br[418] br[419] br[420] br[421] br[422] br[423] br[424] br[425] br[426] br[427] br[428] br[429] br[430] br[431] br[432] br[433] br[434] br[435] br[436] br[437] br[438] br[439] br[440] br[441] br[442] br[443] br[444] br[445] br[446] br[447] br[448] br[449] br[450] br[451] br[452] br[453] br[454] br[455] br[456] br[457] br[458] br[459] br[460] br[461] br[462] br[463] br[464] br[465] br[466] br[467] br[468] br[469] br[470] br[471] br[472] br[473] br[474] br[475] br[476] br[477] br[478] br[479] br[480] br[481] br[482] br[483] br[484] br[485] br[486] br[487] br[488] br[489] br[490] br[491] br[492] br[493] br[494] br[495] br[496] br[497] br[498] br[499] br[500] br[501] br[502] br[503] br[504] br[505] br[506] br[507] br[508] br[509] br[510] br[511] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we wmask[0] wmask[1] wmask[2] wmask[3] wmask[4] wmask[5] wmask[6] wmask[7] wmask[8] wmask[9] wmask[10] wmask[11] wmask[12] wmask[13] wmask[14] wmask[15] din[0] din[1] din[2] din[3] din[4] din[5] din[6] din[7] din[8] din[9] din[10] din[11] din[12] din[13] din[14] din[15] din[16] din[17] din[18] din[19] din[20] din[21] din[22] din[23] din[24] din[25] din[26] din[27] din[28] din[29] din[30] din[31] din[32] din[33] din[34] din[35] din[36] din[37] din[38] din[39] din[40] din[41] din[42] din[43] din[44] din[45] din[46] din[47] din[48] din[49] din[50] din[51] din[52] din[53] din[54] din[55] din[56] din[57] din[58] din[59] din[60] din[61] din[62] din[63] din[64] din[65] din[66] din[67] din[68] din[69] din[70] din[71] din[72] din[73] din[74] din[75] din[76] din[77] din[78] din[79] din[80] din[81] din[82] din[83] din[84] din[85] din[86] din[87] din[88] din[89] din[90] din[91] din[92] din[93] din[94] din[95] din[96] din[97] din[98] din[99] din[100] din[101] din[102] din[103] din[104] din[105] din[106] din[107] din[108] din[109] din[110] din[111] din[112] din[113] din[114] din[115] din[116] din[117] din[118] din[119] din[120] din[121] din[122] din[123] din[124] din[125] din[126] din[127] dout[0] dout[1] dout[2] dout[3] dout[4] dout[5] dout[6] dout[7] dout[8] dout[9] dout[10] dout[11] dout[12] dout[13] dout[14] dout[15] dout[16] dout[17] dout[18] dout[19] dout[20] dout[21] dout[22] dout[23] dout[24] dout[25] dout[26] dout[27] dout[28] dout[29] dout[30] dout[31] dout[32] dout[33] dout[34] dout[35] dout[36] dout[37] dout[38] dout[39] dout[40] dout[41] dout[42] dout[43] dout[44] dout[45] dout[46] dout[47] dout[48] dout[49] dout[50] dout[51] dout[52] dout[53] dout[54] dout[55] dout[56] dout[57] dout[58] dout[59] dout[60] dout[61] dout[62] dout[63] dout[64] dout[65] dout[66] dout[67] dout[68] dout[69] dout[70] dout[71] dout[72] dout[73] dout[74] dout[75] dout[76] dout[77] dout[78] dout[79] dout[80] dout[81] dout[82] dout[83] dout[84] dout[85] dout[86] dout[87] dout[88] dout[89] dout[90] dout[91] dout[92] dout[93] dout[94] dout[95] dout[96] dout[97] dout[98] dout[99] dout[100] dout[101] dout[102] dout[103] dout[104] dout[105] dout[106] dout[107] dout[108] dout[109] dout[110] dout[111] dout[112] dout[113] dout[114] dout[115] dout[116] dout[117] dout[118] dout[119] dout[120] dout[121] dout[122] dout[123] dout[124] dout[125] dout[126] dout[127]

  Xwmask_dffs vdd vss clk rstb wmask[0] wmask[1] wmask[2] wmask[3] wmask[4] wmask[5] wmask[6] wmask[7] wmask[8] wmask[9] wmask[10] wmask[11] wmask[12] wmask[13] wmask[14] wmask[15] wmask_in[0] wmask_in[1] wmask_in[2] wmask_in[3] wmask_in[4] wmask_in[5] wmask_in[6] wmask_in[7] wmask_in[8] wmask_in[9] wmask_in[10] wmask_in[11] wmask_in[12] wmask_in[13] wmask_in[14] wmask_in[15] wmask_in_b[0] wmask_in_b[1] wmask_in_b[2] wmask_in_b[3] wmask_in_b[4] wmask_in_b[5] wmask_in_b[6] wmask_in_b[7] wmask_in_b[8] wmask_in_b[9] wmask_in_b[10] wmask_in_b[11] wmask_in_b[12] wmask_in_b[13] wmask_in_b[14] wmask_in_b[15] dff_array_16
  Xwmask_and_0 vdd vss we_i[0] we_ib[0] we wmask_in[0] decoder_stage_7
  Xwmask_and_1 vdd vss we_i[1] we_ib[1] we wmask_in[1] decoder_stage_7
  Xwmask_and_2 vdd vss we_i[2] we_ib[2] we wmask_in[2] decoder_stage_7
  Xwmask_and_3 vdd vss we_i[3] we_ib[3] we wmask_in[3] decoder_stage_7
  Xwmask_and_4 vdd vss we_i[4] we_ib[4] we wmask_in[4] decoder_stage_7
  Xwmask_and_5 vdd vss we_i[5] we_ib[5] we wmask_in[5] decoder_stage_7
  Xwmask_and_6 vdd vss we_i[6] we_ib[6] we wmask_in[6] decoder_stage_7
  Xwmask_and_7 vdd vss we_i[7] we_ib[7] we wmask_in[7] decoder_stage_7
  Xwmask_and_8 vdd vss we_i[8] we_ib[8] we wmask_in[8] decoder_stage_7
  Xwmask_and_9 vdd vss we_i[9] we_ib[9] we wmask_in[9] decoder_stage_7
  Xwmask_and_10 vdd vss we_i[10] we_ib[10] we wmask_in[10] decoder_stage_7
  Xwmask_and_11 vdd vss we_i[11] we_ib[11] we wmask_in[11] decoder_stage_7
  Xwmask_and_12 vdd vss we_i[12] we_ib[12] we wmask_in[12] decoder_stage_7
  Xwmask_and_13 vdd vss we_i[13] we_ib[13] we wmask_in[13] decoder_stage_7
  Xwmask_and_14 vdd vss we_i[14] we_ib[14] we wmask_in[14] decoder_stage_7
  Xwmask_and_15 vdd vss we_i[15] we_ib[15] we wmask_in[15] decoder_stage_7
  Xcol_group_0 clk rstb vdd vss bl[0] bl[1] bl[2] bl[3] br[0] br[1] br[2] br[3] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[0] we_ib[0] din[0] dout[0] sense_en column
  Xcol_group_1 clk rstb vdd vss bl[4] bl[5] bl[6] bl[7] br[4] br[5] br[6] br[7] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[0] we_ib[0] din[1] dout[1] sense_en column
  Xcol_group_2 clk rstb vdd vss bl[8] bl[9] bl[10] bl[11] br[8] br[9] br[10] br[11] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[0] we_ib[0] din[2] dout[2] sense_en column
  Xcol_group_3 clk rstb vdd vss bl[12] bl[13] bl[14] bl[15] br[12] br[13] br[14] br[15] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[0] we_ib[0] din[3] dout[3] sense_en column
  Xcol_group_4 clk rstb vdd vss bl[16] bl[17] bl[18] bl[19] br[16] br[17] br[18] br[19] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[0] we_ib[0] din[4] dout[4] sense_en column
  Xcol_group_5 clk rstb vdd vss bl[20] bl[21] bl[22] bl[23] br[20] br[21] br[22] br[23] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[0] we_ib[0] din[5] dout[5] sense_en column
  Xcol_group_6 clk rstb vdd vss bl[24] bl[25] bl[26] bl[27] br[24] br[25] br[26] br[27] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[0] we_ib[0] din[6] dout[6] sense_en column
  Xcol_group_7 clk rstb vdd vss bl[28] bl[29] bl[30] bl[31] br[28] br[29] br[30] br[31] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[0] we_ib[0] din[7] dout[7] sense_en column
  Xcol_group_8 clk rstb vdd vss bl[32] bl[33] bl[34] bl[35] br[32] br[33] br[34] br[35] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[1] we_ib[1] din[8] dout[8] sense_en column
  Xcol_group_9 clk rstb vdd vss bl[36] bl[37] bl[38] bl[39] br[36] br[37] br[38] br[39] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[1] we_ib[1] din[9] dout[9] sense_en column
  Xcol_group_10 clk rstb vdd vss bl[40] bl[41] bl[42] bl[43] br[40] br[41] br[42] br[43] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[1] we_ib[1] din[10] dout[10] sense_en column
  Xcol_group_11 clk rstb vdd vss bl[44] bl[45] bl[46] bl[47] br[44] br[45] br[46] br[47] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[1] we_ib[1] din[11] dout[11] sense_en column
  Xcol_group_12 clk rstb vdd vss bl[48] bl[49] bl[50] bl[51] br[48] br[49] br[50] br[51] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[1] we_ib[1] din[12] dout[12] sense_en column
  Xcol_group_13 clk rstb vdd vss bl[52] bl[53] bl[54] bl[55] br[52] br[53] br[54] br[55] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[1] we_ib[1] din[13] dout[13] sense_en column
  Xcol_group_14 clk rstb vdd vss bl[56] bl[57] bl[58] bl[59] br[56] br[57] br[58] br[59] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[1] we_ib[1] din[14] dout[14] sense_en column
  Xcol_group_15 clk rstb vdd vss bl[60] bl[61] bl[62] bl[63] br[60] br[61] br[62] br[63] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[1] we_ib[1] din[15] dout[15] sense_en column
  Xcol_group_16 clk rstb vdd vss bl[64] bl[65] bl[66] bl[67] br[64] br[65] br[66] br[67] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[2] we_ib[2] din[16] dout[16] sense_en column
  Xcol_group_17 clk rstb vdd vss bl[68] bl[69] bl[70] bl[71] br[68] br[69] br[70] br[71] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[2] we_ib[2] din[17] dout[17] sense_en column
  Xcol_group_18 clk rstb vdd vss bl[72] bl[73] bl[74] bl[75] br[72] br[73] br[74] br[75] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[2] we_ib[2] din[18] dout[18] sense_en column
  Xcol_group_19 clk rstb vdd vss bl[76] bl[77] bl[78] bl[79] br[76] br[77] br[78] br[79] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[2] we_ib[2] din[19] dout[19] sense_en column
  Xcol_group_20 clk rstb vdd vss bl[80] bl[81] bl[82] bl[83] br[80] br[81] br[82] br[83] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[2] we_ib[2] din[20] dout[20] sense_en column
  Xcol_group_21 clk rstb vdd vss bl[84] bl[85] bl[86] bl[87] br[84] br[85] br[86] br[87] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[2] we_ib[2] din[21] dout[21] sense_en column
  Xcol_group_22 clk rstb vdd vss bl[88] bl[89] bl[90] bl[91] br[88] br[89] br[90] br[91] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[2] we_ib[2] din[22] dout[22] sense_en column
  Xcol_group_23 clk rstb vdd vss bl[92] bl[93] bl[94] bl[95] br[92] br[93] br[94] br[95] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[2] we_ib[2] din[23] dout[23] sense_en column
  Xcol_group_24 clk rstb vdd vss bl[96] bl[97] bl[98] bl[99] br[96] br[97] br[98] br[99] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[3] we_ib[3] din[24] dout[24] sense_en column
  Xcol_group_25 clk rstb vdd vss bl[100] bl[101] bl[102] bl[103] br[100] br[101] br[102] br[103] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[3] we_ib[3] din[25] dout[25] sense_en column
  Xcol_group_26 clk rstb vdd vss bl[104] bl[105] bl[106] bl[107] br[104] br[105] br[106] br[107] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[3] we_ib[3] din[26] dout[26] sense_en column
  Xcol_group_27 clk rstb vdd vss bl[108] bl[109] bl[110] bl[111] br[108] br[109] br[110] br[111] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[3] we_ib[3] din[27] dout[27] sense_en column
  Xcol_group_28 clk rstb vdd vss bl[112] bl[113] bl[114] bl[115] br[112] br[113] br[114] br[115] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[3] we_ib[3] din[28] dout[28] sense_en column
  Xcol_group_29 clk rstb vdd vss bl[116] bl[117] bl[118] bl[119] br[116] br[117] br[118] br[119] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[3] we_ib[3] din[29] dout[29] sense_en column
  Xcol_group_30 clk rstb vdd vss bl[120] bl[121] bl[122] bl[123] br[120] br[121] br[122] br[123] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[3] we_ib[3] din[30] dout[30] sense_en column
  Xcol_group_31 clk rstb vdd vss bl[124] bl[125] bl[126] bl[127] br[124] br[125] br[126] br[127] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[3] we_ib[3] din[31] dout[31] sense_en column
  Xcol_group_32 clk rstb vdd vss bl[128] bl[129] bl[130] bl[131] br[128] br[129] br[130] br[131] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[4] we_ib[4] din[32] dout[32] sense_en column
  Xcol_group_33 clk rstb vdd vss bl[132] bl[133] bl[134] bl[135] br[132] br[133] br[134] br[135] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[4] we_ib[4] din[33] dout[33] sense_en column
  Xcol_group_34 clk rstb vdd vss bl[136] bl[137] bl[138] bl[139] br[136] br[137] br[138] br[139] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[4] we_ib[4] din[34] dout[34] sense_en column
  Xcol_group_35 clk rstb vdd vss bl[140] bl[141] bl[142] bl[143] br[140] br[141] br[142] br[143] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[4] we_ib[4] din[35] dout[35] sense_en column
  Xcol_group_36 clk rstb vdd vss bl[144] bl[145] bl[146] bl[147] br[144] br[145] br[146] br[147] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[4] we_ib[4] din[36] dout[36] sense_en column
  Xcol_group_37 clk rstb vdd vss bl[148] bl[149] bl[150] bl[151] br[148] br[149] br[150] br[151] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[4] we_ib[4] din[37] dout[37] sense_en column
  Xcol_group_38 clk rstb vdd vss bl[152] bl[153] bl[154] bl[155] br[152] br[153] br[154] br[155] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[4] we_ib[4] din[38] dout[38] sense_en column
  Xcol_group_39 clk rstb vdd vss bl[156] bl[157] bl[158] bl[159] br[156] br[157] br[158] br[159] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[4] we_ib[4] din[39] dout[39] sense_en column
  Xcol_group_40 clk rstb vdd vss bl[160] bl[161] bl[162] bl[163] br[160] br[161] br[162] br[163] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[5] we_ib[5] din[40] dout[40] sense_en column
  Xcol_group_41 clk rstb vdd vss bl[164] bl[165] bl[166] bl[167] br[164] br[165] br[166] br[167] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[5] we_ib[5] din[41] dout[41] sense_en column
  Xcol_group_42 clk rstb vdd vss bl[168] bl[169] bl[170] bl[171] br[168] br[169] br[170] br[171] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[5] we_ib[5] din[42] dout[42] sense_en column
  Xcol_group_43 clk rstb vdd vss bl[172] bl[173] bl[174] bl[175] br[172] br[173] br[174] br[175] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[5] we_ib[5] din[43] dout[43] sense_en column
  Xcol_group_44 clk rstb vdd vss bl[176] bl[177] bl[178] bl[179] br[176] br[177] br[178] br[179] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[5] we_ib[5] din[44] dout[44] sense_en column
  Xcol_group_45 clk rstb vdd vss bl[180] bl[181] bl[182] bl[183] br[180] br[181] br[182] br[183] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[5] we_ib[5] din[45] dout[45] sense_en column
  Xcol_group_46 clk rstb vdd vss bl[184] bl[185] bl[186] bl[187] br[184] br[185] br[186] br[187] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[5] we_ib[5] din[46] dout[46] sense_en column
  Xcol_group_47 clk rstb vdd vss bl[188] bl[189] bl[190] bl[191] br[188] br[189] br[190] br[191] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[5] we_ib[5] din[47] dout[47] sense_en column
  Xcol_group_48 clk rstb vdd vss bl[192] bl[193] bl[194] bl[195] br[192] br[193] br[194] br[195] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[6] we_ib[6] din[48] dout[48] sense_en column
  Xcol_group_49 clk rstb vdd vss bl[196] bl[197] bl[198] bl[199] br[196] br[197] br[198] br[199] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[6] we_ib[6] din[49] dout[49] sense_en column
  Xcol_group_50 clk rstb vdd vss bl[200] bl[201] bl[202] bl[203] br[200] br[201] br[202] br[203] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[6] we_ib[6] din[50] dout[50] sense_en column
  Xcol_group_51 clk rstb vdd vss bl[204] bl[205] bl[206] bl[207] br[204] br[205] br[206] br[207] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[6] we_ib[6] din[51] dout[51] sense_en column
  Xcol_group_52 clk rstb vdd vss bl[208] bl[209] bl[210] bl[211] br[208] br[209] br[210] br[211] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[6] we_ib[6] din[52] dout[52] sense_en column
  Xcol_group_53 clk rstb vdd vss bl[212] bl[213] bl[214] bl[215] br[212] br[213] br[214] br[215] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[6] we_ib[6] din[53] dout[53] sense_en column
  Xcol_group_54 clk rstb vdd vss bl[216] bl[217] bl[218] bl[219] br[216] br[217] br[218] br[219] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[6] we_ib[6] din[54] dout[54] sense_en column
  Xcol_group_55 clk rstb vdd vss bl[220] bl[221] bl[222] bl[223] br[220] br[221] br[222] br[223] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[6] we_ib[6] din[55] dout[55] sense_en column
  Xcol_group_56 clk rstb vdd vss bl[224] bl[225] bl[226] bl[227] br[224] br[225] br[226] br[227] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[7] we_ib[7] din[56] dout[56] sense_en column
  Xcol_group_57 clk rstb vdd vss bl[228] bl[229] bl[230] bl[231] br[228] br[229] br[230] br[231] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[7] we_ib[7] din[57] dout[57] sense_en column
  Xcol_group_58 clk rstb vdd vss bl[232] bl[233] bl[234] bl[235] br[232] br[233] br[234] br[235] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[7] we_ib[7] din[58] dout[58] sense_en column
  Xcol_group_59 clk rstb vdd vss bl[236] bl[237] bl[238] bl[239] br[236] br[237] br[238] br[239] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[7] we_ib[7] din[59] dout[59] sense_en column
  Xcol_group_60 clk rstb vdd vss bl[240] bl[241] bl[242] bl[243] br[240] br[241] br[242] br[243] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[7] we_ib[7] din[60] dout[60] sense_en column
  Xcol_group_61 clk rstb vdd vss bl[244] bl[245] bl[246] bl[247] br[244] br[245] br[246] br[247] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[7] we_ib[7] din[61] dout[61] sense_en column
  Xcol_group_62 clk rstb vdd vss bl[248] bl[249] bl[250] bl[251] br[248] br[249] br[250] br[251] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[7] we_ib[7] din[62] dout[62] sense_en column
  Xcol_group_63 clk rstb vdd vss bl[252] bl[253] bl[254] bl[255] br[252] br[253] br[254] br[255] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[7] we_ib[7] din[63] dout[63] sense_en column
  Xcol_group_64 clk rstb vdd vss bl[256] bl[257] bl[258] bl[259] br[256] br[257] br[258] br[259] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[8] we_ib[8] din[64] dout[64] sense_en column
  Xcol_group_65 clk rstb vdd vss bl[260] bl[261] bl[262] bl[263] br[260] br[261] br[262] br[263] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[8] we_ib[8] din[65] dout[65] sense_en column
  Xcol_group_66 clk rstb vdd vss bl[264] bl[265] bl[266] bl[267] br[264] br[265] br[266] br[267] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[8] we_ib[8] din[66] dout[66] sense_en column
  Xcol_group_67 clk rstb vdd vss bl[268] bl[269] bl[270] bl[271] br[268] br[269] br[270] br[271] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[8] we_ib[8] din[67] dout[67] sense_en column
  Xcol_group_68 clk rstb vdd vss bl[272] bl[273] bl[274] bl[275] br[272] br[273] br[274] br[275] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[8] we_ib[8] din[68] dout[68] sense_en column
  Xcol_group_69 clk rstb vdd vss bl[276] bl[277] bl[278] bl[279] br[276] br[277] br[278] br[279] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[8] we_ib[8] din[69] dout[69] sense_en column
  Xcol_group_70 clk rstb vdd vss bl[280] bl[281] bl[282] bl[283] br[280] br[281] br[282] br[283] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[8] we_ib[8] din[70] dout[70] sense_en column
  Xcol_group_71 clk rstb vdd vss bl[284] bl[285] bl[286] bl[287] br[284] br[285] br[286] br[287] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[8] we_ib[8] din[71] dout[71] sense_en column
  Xcol_group_72 clk rstb vdd vss bl[288] bl[289] bl[290] bl[291] br[288] br[289] br[290] br[291] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[9] we_ib[9] din[72] dout[72] sense_en column
  Xcol_group_73 clk rstb vdd vss bl[292] bl[293] bl[294] bl[295] br[292] br[293] br[294] br[295] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[9] we_ib[9] din[73] dout[73] sense_en column
  Xcol_group_74 clk rstb vdd vss bl[296] bl[297] bl[298] bl[299] br[296] br[297] br[298] br[299] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[9] we_ib[9] din[74] dout[74] sense_en column
  Xcol_group_75 clk rstb vdd vss bl[300] bl[301] bl[302] bl[303] br[300] br[301] br[302] br[303] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[9] we_ib[9] din[75] dout[75] sense_en column
  Xcol_group_76 clk rstb vdd vss bl[304] bl[305] bl[306] bl[307] br[304] br[305] br[306] br[307] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[9] we_ib[9] din[76] dout[76] sense_en column
  Xcol_group_77 clk rstb vdd vss bl[308] bl[309] bl[310] bl[311] br[308] br[309] br[310] br[311] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[9] we_ib[9] din[77] dout[77] sense_en column
  Xcol_group_78 clk rstb vdd vss bl[312] bl[313] bl[314] bl[315] br[312] br[313] br[314] br[315] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[9] we_ib[9] din[78] dout[78] sense_en column
  Xcol_group_79 clk rstb vdd vss bl[316] bl[317] bl[318] bl[319] br[316] br[317] br[318] br[319] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[9] we_ib[9] din[79] dout[79] sense_en column
  Xcol_group_80 clk rstb vdd vss bl[320] bl[321] bl[322] bl[323] br[320] br[321] br[322] br[323] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[10] we_ib[10] din[80] dout[80] sense_en column
  Xcol_group_81 clk rstb vdd vss bl[324] bl[325] bl[326] bl[327] br[324] br[325] br[326] br[327] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[10] we_ib[10] din[81] dout[81] sense_en column
  Xcol_group_82 clk rstb vdd vss bl[328] bl[329] bl[330] bl[331] br[328] br[329] br[330] br[331] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[10] we_ib[10] din[82] dout[82] sense_en column
  Xcol_group_83 clk rstb vdd vss bl[332] bl[333] bl[334] bl[335] br[332] br[333] br[334] br[335] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[10] we_ib[10] din[83] dout[83] sense_en column
  Xcol_group_84 clk rstb vdd vss bl[336] bl[337] bl[338] bl[339] br[336] br[337] br[338] br[339] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[10] we_ib[10] din[84] dout[84] sense_en column
  Xcol_group_85 clk rstb vdd vss bl[340] bl[341] bl[342] bl[343] br[340] br[341] br[342] br[343] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[10] we_ib[10] din[85] dout[85] sense_en column
  Xcol_group_86 clk rstb vdd vss bl[344] bl[345] bl[346] bl[347] br[344] br[345] br[346] br[347] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[10] we_ib[10] din[86] dout[86] sense_en column
  Xcol_group_87 clk rstb vdd vss bl[348] bl[349] bl[350] bl[351] br[348] br[349] br[350] br[351] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[10] we_ib[10] din[87] dout[87] sense_en column
  Xcol_group_88 clk rstb vdd vss bl[352] bl[353] bl[354] bl[355] br[352] br[353] br[354] br[355] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[11] we_ib[11] din[88] dout[88] sense_en column
  Xcol_group_89 clk rstb vdd vss bl[356] bl[357] bl[358] bl[359] br[356] br[357] br[358] br[359] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[11] we_ib[11] din[89] dout[89] sense_en column
  Xcol_group_90 clk rstb vdd vss bl[360] bl[361] bl[362] bl[363] br[360] br[361] br[362] br[363] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[11] we_ib[11] din[90] dout[90] sense_en column
  Xcol_group_91 clk rstb vdd vss bl[364] bl[365] bl[366] bl[367] br[364] br[365] br[366] br[367] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[11] we_ib[11] din[91] dout[91] sense_en column
  Xcol_group_92 clk rstb vdd vss bl[368] bl[369] bl[370] bl[371] br[368] br[369] br[370] br[371] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[11] we_ib[11] din[92] dout[92] sense_en column
  Xcol_group_93 clk rstb vdd vss bl[372] bl[373] bl[374] bl[375] br[372] br[373] br[374] br[375] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[11] we_ib[11] din[93] dout[93] sense_en column
  Xcol_group_94 clk rstb vdd vss bl[376] bl[377] bl[378] bl[379] br[376] br[377] br[378] br[379] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[11] we_ib[11] din[94] dout[94] sense_en column
  Xcol_group_95 clk rstb vdd vss bl[380] bl[381] bl[382] bl[383] br[380] br[381] br[382] br[383] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[11] we_ib[11] din[95] dout[95] sense_en column
  Xcol_group_96 clk rstb vdd vss bl[384] bl[385] bl[386] bl[387] br[384] br[385] br[386] br[387] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[12] we_ib[12] din[96] dout[96] sense_en column
  Xcol_group_97 clk rstb vdd vss bl[388] bl[389] bl[390] bl[391] br[388] br[389] br[390] br[391] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[12] we_ib[12] din[97] dout[97] sense_en column
  Xcol_group_98 clk rstb vdd vss bl[392] bl[393] bl[394] bl[395] br[392] br[393] br[394] br[395] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[12] we_ib[12] din[98] dout[98] sense_en column
  Xcol_group_99 clk rstb vdd vss bl[396] bl[397] bl[398] bl[399] br[396] br[397] br[398] br[399] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[12] we_ib[12] din[99] dout[99] sense_en column
  Xcol_group_100 clk rstb vdd vss bl[400] bl[401] bl[402] bl[403] br[400] br[401] br[402] br[403] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[12] we_ib[12] din[100] dout[100] sense_en column
  Xcol_group_101 clk rstb vdd vss bl[404] bl[405] bl[406] bl[407] br[404] br[405] br[406] br[407] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[12] we_ib[12] din[101] dout[101] sense_en column
  Xcol_group_102 clk rstb vdd vss bl[408] bl[409] bl[410] bl[411] br[408] br[409] br[410] br[411] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[12] we_ib[12] din[102] dout[102] sense_en column
  Xcol_group_103 clk rstb vdd vss bl[412] bl[413] bl[414] bl[415] br[412] br[413] br[414] br[415] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[12] we_ib[12] din[103] dout[103] sense_en column
  Xcol_group_104 clk rstb vdd vss bl[416] bl[417] bl[418] bl[419] br[416] br[417] br[418] br[419] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[13] we_ib[13] din[104] dout[104] sense_en column
  Xcol_group_105 clk rstb vdd vss bl[420] bl[421] bl[422] bl[423] br[420] br[421] br[422] br[423] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[13] we_ib[13] din[105] dout[105] sense_en column
  Xcol_group_106 clk rstb vdd vss bl[424] bl[425] bl[426] bl[427] br[424] br[425] br[426] br[427] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[13] we_ib[13] din[106] dout[106] sense_en column
  Xcol_group_107 clk rstb vdd vss bl[428] bl[429] bl[430] bl[431] br[428] br[429] br[430] br[431] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[13] we_ib[13] din[107] dout[107] sense_en column
  Xcol_group_108 clk rstb vdd vss bl[432] bl[433] bl[434] bl[435] br[432] br[433] br[434] br[435] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[13] we_ib[13] din[108] dout[108] sense_en column
  Xcol_group_109 clk rstb vdd vss bl[436] bl[437] bl[438] bl[439] br[436] br[437] br[438] br[439] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[13] we_ib[13] din[109] dout[109] sense_en column
  Xcol_group_110 clk rstb vdd vss bl[440] bl[441] bl[442] bl[443] br[440] br[441] br[442] br[443] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[13] we_ib[13] din[110] dout[110] sense_en column
  Xcol_group_111 clk rstb vdd vss bl[444] bl[445] bl[446] bl[447] br[444] br[445] br[446] br[447] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[13] we_ib[13] din[111] dout[111] sense_en column
  Xcol_group_112 clk rstb vdd vss bl[448] bl[449] bl[450] bl[451] br[448] br[449] br[450] br[451] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[14] we_ib[14] din[112] dout[112] sense_en column
  Xcol_group_113 clk rstb vdd vss bl[452] bl[453] bl[454] bl[455] br[452] br[453] br[454] br[455] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[14] we_ib[14] din[113] dout[113] sense_en column
  Xcol_group_114 clk rstb vdd vss bl[456] bl[457] bl[458] bl[459] br[456] br[457] br[458] br[459] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[14] we_ib[14] din[114] dout[114] sense_en column
  Xcol_group_115 clk rstb vdd vss bl[460] bl[461] bl[462] bl[463] br[460] br[461] br[462] br[463] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[14] we_ib[14] din[115] dout[115] sense_en column
  Xcol_group_116 clk rstb vdd vss bl[464] bl[465] bl[466] bl[467] br[464] br[465] br[466] br[467] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[14] we_ib[14] din[116] dout[116] sense_en column
  Xcol_group_117 clk rstb vdd vss bl[468] bl[469] bl[470] bl[471] br[468] br[469] br[470] br[471] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[14] we_ib[14] din[117] dout[117] sense_en column
  Xcol_group_118 clk rstb vdd vss bl[472] bl[473] bl[474] bl[475] br[472] br[473] br[474] br[475] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[14] we_ib[14] din[118] dout[118] sense_en column
  Xcol_group_119 clk rstb vdd vss bl[476] bl[477] bl[478] bl[479] br[476] br[477] br[478] br[479] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[14] we_ib[14] din[119] dout[119] sense_en column
  Xcol_group_120 clk rstb vdd vss bl[480] bl[481] bl[482] bl[483] br[480] br[481] br[482] br[483] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[15] we_ib[15] din[120] dout[120] sense_en column
  Xcol_group_121 clk rstb vdd vss bl[484] bl[485] bl[486] bl[487] br[484] br[485] br[486] br[487] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[15] we_ib[15] din[121] dout[121] sense_en column
  Xcol_group_122 clk rstb vdd vss bl[488] bl[489] bl[490] bl[491] br[488] br[489] br[490] br[491] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[15] we_ib[15] din[122] dout[122] sense_en column
  Xcol_group_123 clk rstb vdd vss bl[492] bl[493] bl[494] bl[495] br[492] br[493] br[494] br[495] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[15] we_ib[15] din[123] dout[123] sense_en column
  Xcol_group_124 clk rstb vdd vss bl[496] bl[497] bl[498] bl[499] br[496] br[497] br[498] br[499] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[15] we_ib[15] din[124] dout[124] sense_en column
  Xcol_group_125 clk rstb vdd vss bl[500] bl[501] bl[502] bl[503] br[500] br[501] br[502] br[503] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[15] we_ib[15] din[125] dout[125] sense_en column
  Xcol_group_126 clk rstb vdd vss bl[504] bl[505] bl[506] bl[507] br[504] br[505] br[506] br[507] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[15] we_ib[15] din[126] dout[126] sense_en column
  Xcol_group_127 clk rstb vdd vss bl[508] bl[509] bl[510] bl[511] br[508] br[509] br[510] br[511] pc_b sel[0] sel[1] sel[2] sel[3] sel_b[0] sel_b[1] sel_b[2] sel_b[3] we_i[15] we_ib[15] din[127] dout[127] sense_en column

.ENDS col_peripherals

.SUBCKT mos_w800_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=0.800


.ENDS mos_w800_l150_m1_nf1_id0

.SUBCKT mos_w1200_l150_m1_nf1_id0 d g s b

  X0 d g s b sky130_fd_pr__nfet_01v8 l=0.150 nf=1 w=1.200


.ENDS mos_w1200_l150_m1_nf1_id0

.SUBCKT mos_w1700_l150_m1_nf1_id1 d g s b

  X0 d g s b sky130_fd_pr__pfet_01v8 l=0.150 nf=1 w=1.700


.ENDS mos_w1700_l150_m1_nf1_id1

.SUBCKT column_mos vdd vss bl

  Xgate_nmos vss bl vss vss mos_w800_l150_m1_nf1_id0
  Xdrain_nmos bl vss vss vss mos_w1200_l150_m1_nf1_id0
  Xdrain_pmos bl vdd vdd vdd mos_w1700_l150_m1_nf1_id1

.ENDS column_mos

.SUBCKT column_mos_1 vdd vss bl

  Xdrain_nmos bl vss vss vss mos_w1200_l150_m1_nf1_id0
  Xdrain_pmos bl vdd vdd vdd mos_w1700_l150_m1_nf1_id1

.ENDS column_mos_1

.SUBCKT replica_column_mos vdd vss bl

  Xunit0 vdd vss bl column_mos
  Xunit1 vdd vss bl column_mos_1
  Xunit2 vdd vss bl column_mos_1

.ENDS replica_column_mos

.SUBCKT sram22_inner vdd vss clk we ce rstb addr[0] addr[1] addr[2] addr[3] addr[4] addr[5] addr[6] addr[7] wmask[0] wmask[1] wmask[2] wmask[3] wmask[4] wmask[5] wmask[6] wmask[7] wmask[8] wmask[9] wmask[10] wmask[11] wmask[12] wmask[13] wmask[14] wmask[15] din[0] din[1] din[2] din[3] din[4] din[5] din[6] din[7] din[8] din[9] din[10] din[11] din[12] din[13] din[14] din[15] din[16] din[17] din[18] din[19] din[20] din[21] din[22] din[23] din[24] din[25] din[26] din[27] din[28] din[29] din[30] din[31] din[32] din[33] din[34] din[35] din[36] din[37] din[38] din[39] din[40] din[41] din[42] din[43] din[44] din[45] din[46] din[47] din[48] din[49] din[50] din[51] din[52] din[53] din[54] din[55] din[56] din[57] din[58] din[59] din[60] din[61] din[62] din[63] din[64] din[65] din[66] din[67] din[68] din[69] din[70] din[71] din[72] din[73] din[74] din[75] din[76] din[77] din[78] din[79] din[80] din[81] din[82] din[83] din[84] din[85] din[86] din[87] din[88] din[89] din[90] din[91] din[92] din[93] din[94] din[95] din[96] din[97] din[98] din[99] din[100] din[101] din[102] din[103] din[104] din[105] din[106] din[107] din[108] din[109] din[110] din[111] din[112] din[113] din[114] din[115] din[116] din[117] din[118] din[119] din[120] din[121] din[122] din[123] din[124] din[125] din[126] din[127] dout[0] dout[1] dout[2] dout[3] dout[4] dout[5] dout[6] dout[7] dout[8] dout[9] dout[10] dout[11] dout[12] dout[13] dout[14] dout[15] dout[16] dout[17] dout[18] dout[19] dout[20] dout[21] dout[22] dout[23] dout[24] dout[25] dout[26] dout[27] dout[28] dout[29] dout[30] dout[31] dout[32] dout[33] dout[34] dout[35] dout[36] dout[37] dout[38] dout[39] dout[40] dout[41] dout[42] dout[43] dout[44] dout[45] dout[46] dout[47] dout[48] dout[49] dout[50] dout[51] dout[52] dout[53] dout[54] dout[55] dout[56] dout[57] dout[58] dout[59] dout[60] dout[61] dout[62] dout[63] dout[64] dout[65] dout[66] dout[67] dout[68] dout[69] dout[70] dout[71] dout[72] dout[73] dout[74] dout[75] dout[76] dout[77] dout[78] dout[79] dout[80] dout[81] dout[82] dout[83] dout[84] dout[85] dout[86] dout[87] dout[88] dout[89] dout[90] dout[91] dout[92] dout[93] dout[94] dout[95] dout[96] dout[97] dout[98] dout[99] dout[100] dout[101] dout[102] dout[103] dout[104] dout[105] dout[106] dout[107] dout[108] dout[109] dout[110] dout[111] dout[112] dout[113] dout[114] dout[115] dout[116] dout[117] dout[118] dout[119] dout[120] dout[121] dout[122] dout[123] dout[124] dout[125] dout[126] dout[127]

  Xaddr_gate vdd vss addr_gated[0] addr_gated[1] addr_gated[2] addr_gated[3] addr_gated[4] addr_gated[5] addr_b_gated[0] addr_b_gated[1] addr_b_gated[2] addr_b_gated[3] addr_b_gated[4] addr_b_gated[5] addr_gate_y_b_noconn[0] addr_gate_y_b_noconn[1] addr_gate_y_b_noconn[2] addr_gate_y_b_noconn[3] addr_gate_y_b_noconn[4] addr_gate_y_b_noconn[5] addr_gate_y_b_noconn[6] addr_gate_y_b_noconn[7] addr_gate_y_b_noconn[8] addr_gate_y_b_noconn[9] addr_gate_y_b_noconn[10] addr_gate_y_b_noconn[11] wl_en addr_in[2] addr_in[3] addr_in[4] addr_in[5] addr_in[6] addr_in[7] addr_in_b[2] addr_in_b[3] addr_in_b[4] addr_in_b[5] addr_in_b[6] addr_in_b[7] decoder_stage
  Xdecoder vdd vss wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl_b[0] wl_b[1] wl_b[2] wl_b[3] wl_b[4] wl_b[5] wl_b[6] wl_b[7] wl_b[8] wl_b[9] wl_b[10] wl_b[11] wl_b[12] wl_b[13] wl_b[14] wl_b[15] wl_b[16] wl_b[17] wl_b[18] wl_b[19] wl_b[20] wl_b[21] wl_b[22] wl_b[23] wl_b[24] wl_b[25] wl_b[26] wl_b[27] wl_b[28] wl_b[29] wl_b[30] wl_b[31] wl_b[32] wl_b[33] wl_b[34] wl_b[35] wl_b[36] wl_b[37] wl_b[38] wl_b[39] wl_b[40] wl_b[41] wl_b[42] wl_b[43] wl_b[44] wl_b[45] wl_b[46] wl_b[47] wl_b[48] wl_b[49] wl_b[50] wl_b[51] wl_b[52] wl_b[53] wl_b[54] wl_b[55] wl_b[56] wl_b[57] wl_b[58] wl_b[59] wl_b[60] wl_b[61] wl_b[62] wl_b[63] addr_b_gated[0] addr_gated[0] addr_b_gated[1] addr_gated[1] addr_b_gated[2] addr_gated[2] addr_b_gated[3] addr_gated[3] addr_b_gated[4] addr_gated[4] addr_b_gated[5] addr_gated[5] decoder
  Xcolumn_decoder vdd vss col_sel[0] col_sel[1] col_sel[2] col_sel[3] col_sel_b[0] col_sel_b[1] col_sel_b[2] col_sel_b[3] addr_in_b[0] addr_in[0] addr_in_b[1] addr_in[1] decoder_1
  Xcontrol_logic clk ce_in we_in rstb rbl sense_en0 pc_b0 rwl wl_en0 write_driver_en0 vdd vss control_logic_replica_v2
  Xpc_b_buffer vdd vss pc_b pc pc_b0 decoder_stage_1
  Xwlen_buffer vdd vss wl_en wl_en_b wl_en0 decoder_stage_2
  Xwrite_driver_en_buffer vdd vss write_driver_en write_driver_en_b write_driver_en0 decoder_stage_3
  Xsense_en_buffer vdd vss sense_en sense_en_b sense_en0 decoder_stage_4
  Xaddr_we_ce_dffs vdd vss clk rstb addr[0] addr[1] addr[2] addr[3] addr[4] addr[5] addr[6] addr[7] we ce addr_in[0] addr_in[1] addr_in[2] addr_in[3] addr_in[4] addr_in[5] addr_in[6] addr_in[7] we_in ce_in addr_in_b[0] addr_in_b[1] addr_in_b[2] addr_in_b[3] addr_in_b[4] addr_in_b[5] addr_in_b[6] addr_in_b[7] we_in_b ce_in_b dff_array_10
  Xbitcell_array vdd vss vdd vdd bl[0] bl[1] bl[2] bl[3] bl[4] bl[5] bl[6] bl[7] bl[8] bl[9] bl[10] bl[11] bl[12] bl[13] bl[14] bl[15] bl[16] bl[17] bl[18] bl[19] bl[20] bl[21] bl[22] bl[23] bl[24] bl[25] bl[26] bl[27] bl[28] bl[29] bl[30] bl[31] bl[32] bl[33] bl[34] bl[35] bl[36] bl[37] bl[38] bl[39] bl[40] bl[41] bl[42] bl[43] bl[44] bl[45] bl[46] bl[47] bl[48] bl[49] bl[50] bl[51] bl[52] bl[53] bl[54] bl[55] bl[56] bl[57] bl[58] bl[59] bl[60] bl[61] bl[62] bl[63] bl[64] bl[65] bl[66] bl[67] bl[68] bl[69] bl[70] bl[71] bl[72] bl[73] bl[74] bl[75] bl[76] bl[77] bl[78] bl[79] bl[80] bl[81] bl[82] bl[83] bl[84] bl[85] bl[86] bl[87] bl[88] bl[89] bl[90] bl[91] bl[92] bl[93] bl[94] bl[95] bl[96] bl[97] bl[98] bl[99] bl[100] bl[101] bl[102] bl[103] bl[104] bl[105] bl[106] bl[107] bl[108] bl[109] bl[110] bl[111] bl[112] bl[113] bl[114] bl[115] bl[116] bl[117] bl[118] bl[119] bl[120] bl[121] bl[122] bl[123] bl[124] bl[125] bl[126] bl[127] bl[128] bl[129] bl[130] bl[131] bl[132] bl[133] bl[134] bl[135] bl[136] bl[137] bl[138] bl[139] bl[140] bl[141] bl[142] bl[143] bl[144] bl[145] bl[146] bl[147] bl[148] bl[149] bl[150] bl[151] bl[152] bl[153] bl[154] bl[155] bl[156] bl[157] bl[158] bl[159] bl[160] bl[161] bl[162] bl[163] bl[164] bl[165] bl[166] bl[167] bl[168] bl[169] bl[170] bl[171] bl[172] bl[173] bl[174] bl[175] bl[176] bl[177] bl[178] bl[179] bl[180] bl[181] bl[182] bl[183] bl[184] bl[185] bl[186] bl[187] bl[188] bl[189] bl[190] bl[191] bl[192] bl[193] bl[194] bl[195] bl[196] bl[197] bl[198] bl[199] bl[200] bl[201] bl[202] bl[203] bl[204] bl[205] bl[206] bl[207] bl[208] bl[209] bl[210] bl[211] bl[212] bl[213] bl[214] bl[215] bl[216] bl[217] bl[218] bl[219] bl[220] bl[221] bl[222] bl[223] bl[224] bl[225] bl[226] bl[227] bl[228] bl[229] bl[230] bl[231] bl[232] bl[233] bl[234] bl[235] bl[236] bl[237] bl[238] bl[239] bl[240] bl[241] bl[242] bl[243] bl[244] bl[245] bl[246] bl[247] bl[248] bl[249] bl[250] bl[251] bl[252] bl[253] bl[254] bl[255] bl[256] bl[257] bl[258] bl[259] bl[260] bl[261] bl[262] bl[263] bl[264] bl[265] bl[266] bl[267] bl[268] bl[269] bl[270] bl[271] bl[272] bl[273] bl[274] bl[275] bl[276] bl[277] bl[278] bl[279] bl[280] bl[281] bl[282] bl[283] bl[284] bl[285] bl[286] bl[287] bl[288] bl[289] bl[290] bl[291] bl[292] bl[293] bl[294] bl[295] bl[296] bl[297] bl[298] bl[299] bl[300] bl[301] bl[302] bl[303] bl[304] bl[305] bl[306] bl[307] bl[308] bl[309] bl[310] bl[311] bl[312] bl[313] bl[314] bl[315] bl[316] bl[317] bl[318] bl[319] bl[320] bl[321] bl[322] bl[323] bl[324] bl[325] bl[326] bl[327] bl[328] bl[329] bl[330] bl[331] bl[332] bl[333] bl[334] bl[335] bl[336] bl[337] bl[338] bl[339] bl[340] bl[341] bl[342] bl[343] bl[344] bl[345] bl[346] bl[347] bl[348] bl[349] bl[350] bl[351] bl[352] bl[353] bl[354] bl[355] bl[356] bl[357] bl[358] bl[359] bl[360] bl[361] bl[362] bl[363] bl[364] bl[365] bl[366] bl[367] bl[368] bl[369] bl[370] bl[371] bl[372] bl[373] bl[374] bl[375] bl[376] bl[377] bl[378] bl[379] bl[380] bl[381] bl[382] bl[383] bl[384] bl[385] bl[386] bl[387] bl[388] bl[389] bl[390] bl[391] bl[392] bl[393] bl[394] bl[395] bl[396] bl[397] bl[398] bl[399] bl[400] bl[401] bl[402] bl[403] bl[404] bl[405] bl[406] bl[407] bl[408] bl[409] bl[410] bl[411] bl[412] bl[413] bl[414] bl[415] bl[416] bl[417] bl[418] bl[419] bl[420] bl[421] bl[422] bl[423] bl[424] bl[425] bl[426] bl[427] bl[428] bl[429] bl[430] bl[431] bl[432] bl[433] bl[434] bl[435] bl[436] bl[437] bl[438] bl[439] bl[440] bl[441] bl[442] bl[443] bl[444] bl[445] bl[446] bl[447] bl[448] bl[449] bl[450] bl[451] bl[452] bl[453] bl[454] bl[455] bl[456] bl[457] bl[458] bl[459] bl[460] bl[461] bl[462] bl[463] bl[464] bl[465] bl[466] bl[467] bl[468] bl[469] bl[470] bl[471] bl[472] bl[473] bl[474] bl[475] bl[476] bl[477] bl[478] bl[479] bl[480] bl[481] bl[482] bl[483] bl[484] bl[485] bl[486] bl[487] bl[488] bl[489] bl[490] bl[491] bl[492] bl[493] bl[494] bl[495] bl[496] bl[497] bl[498] bl[499] bl[500] bl[501] bl[502] bl[503] bl[504] bl[505] bl[506] bl[507] bl[508] bl[509] bl[510] bl[511] br[0] br[1] br[2] br[3] br[4] br[5] br[6] br[7] br[8] br[9] br[10] br[11] br[12] br[13] br[14] br[15] br[16] br[17] br[18] br[19] br[20] br[21] br[22] br[23] br[24] br[25] br[26] br[27] br[28] br[29] br[30] br[31] br[32] br[33] br[34] br[35] br[36] br[37] br[38] br[39] br[40] br[41] br[42] br[43] br[44] br[45] br[46] br[47] br[48] br[49] br[50] br[51] br[52] br[53] br[54] br[55] br[56] br[57] br[58] br[59] br[60] br[61] br[62] br[63] br[64] br[65] br[66] br[67] br[68] br[69] br[70] br[71] br[72] br[73] br[74] br[75] br[76] br[77] br[78] br[79] br[80] br[81] br[82] br[83] br[84] br[85] br[86] br[87] br[88] br[89] br[90] br[91] br[92] br[93] br[94] br[95] br[96] br[97] br[98] br[99] br[100] br[101] br[102] br[103] br[104] br[105] br[106] br[107] br[108] br[109] br[110] br[111] br[112] br[113] br[114] br[115] br[116] br[117] br[118] br[119] br[120] br[121] br[122] br[123] br[124] br[125] br[126] br[127] br[128] br[129] br[130] br[131] br[132] br[133] br[134] br[135] br[136] br[137] br[138] br[139] br[140] br[141] br[142] br[143] br[144] br[145] br[146] br[147] br[148] br[149] br[150] br[151] br[152] br[153] br[154] br[155] br[156] br[157] br[158] br[159] br[160] br[161] br[162] br[163] br[164] br[165] br[166] br[167] br[168] br[169] br[170] br[171] br[172] br[173] br[174] br[175] br[176] br[177] br[178] br[179] br[180] br[181] br[182] br[183] br[184] br[185] br[186] br[187] br[188] br[189] br[190] br[191] br[192] br[193] br[194] br[195] br[196] br[197] br[198] br[199] br[200] br[201] br[202] br[203] br[204] br[205] br[206] br[207] br[208] br[209] br[210] br[211] br[212] br[213] br[214] br[215] br[216] br[217] br[218] br[219] br[220] br[221] br[222] br[223] br[224] br[225] br[226] br[227] br[228] br[229] br[230] br[231] br[232] br[233] br[234] br[235] br[236] br[237] br[238] br[239] br[240] br[241] br[242] br[243] br[244] br[245] br[246] br[247] br[248] br[249] br[250] br[251] br[252] br[253] br[254] br[255] br[256] br[257] br[258] br[259] br[260] br[261] br[262] br[263] br[264] br[265] br[266] br[267] br[268] br[269] br[270] br[271] br[272] br[273] br[274] br[275] br[276] br[277] br[278] br[279] br[280] br[281] br[282] br[283] br[284] br[285] br[286] br[287] br[288] br[289] br[290] br[291] br[292] br[293] br[294] br[295] br[296] br[297] br[298] br[299] br[300] br[301] br[302] br[303] br[304] br[305] br[306] br[307] br[308] br[309] br[310] br[311] br[312] br[313] br[314] br[315] br[316] br[317] br[318] br[319] br[320] br[321] br[322] br[323] br[324] br[325] br[326] br[327] br[328] br[329] br[330] br[331] br[332] br[333] br[334] br[335] br[336] br[337] br[338] br[339] br[340] br[341] br[342] br[343] br[344] br[345] br[346] br[347] br[348] br[349] br[350] br[351] br[352] br[353] br[354] br[355] br[356] br[357] br[358] br[359] br[360] br[361] br[362] br[363] br[364] br[365] br[366] br[367] br[368] br[369] br[370] br[371] br[372] br[373] br[374] br[375] br[376] br[377] br[378] br[379] br[380] br[381] br[382] br[383] br[384] br[385] br[386] br[387] br[388] br[389] br[390] br[391] br[392] br[393] br[394] br[395] br[396] br[397] br[398] br[399] br[400] br[401] br[402] br[403] br[404] br[405] br[406] br[407] br[408] br[409] br[410] br[411] br[412] br[413] br[414] br[415] br[416] br[417] br[418] br[419] br[420] br[421] br[422] br[423] br[424] br[425] br[426] br[427] br[428] br[429] br[430] br[431] br[432] br[433] br[434] br[435] br[436] br[437] br[438] br[439] br[440] br[441] br[442] br[443] br[444] br[445] br[446] br[447] br[448] br[449] br[450] br[451] br[452] br[453] br[454] br[455] br[456] br[457] br[458] br[459] br[460] br[461] br[462] br[463] br[464] br[465] br[466] br[467] br[468] br[469] br[470] br[471] br[472] br[473] br[474] br[475] br[476] br[477] br[478] br[479] br[480] br[481] br[482] br[483] br[484] br[485] br[486] br[487] br[488] br[489] br[490] br[491] br[492] br[493] br[494] br[495] br[496] br[497] br[498] br[499] br[500] br[501] br[502] br[503] br[504] br[505] br[506] br[507] br[508] br[509] br[510] br[511] wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] sp_cell_array
  Xreplica_bitcell_array vdd vss rbl rbr rwl replica_cell_array
  Xcol_circuitry clk rstb vdd vss sense_en bl[0] bl[1] bl[2] bl[3] bl[4] bl[5] bl[6] bl[7] bl[8] bl[9] bl[10] bl[11] bl[12] bl[13] bl[14] bl[15] bl[16] bl[17] bl[18] bl[19] bl[20] bl[21] bl[22] bl[23] bl[24] bl[25] bl[26] bl[27] bl[28] bl[29] bl[30] bl[31] bl[32] bl[33] bl[34] bl[35] bl[36] bl[37] bl[38] bl[39] bl[40] bl[41] bl[42] bl[43] bl[44] bl[45] bl[46] bl[47] bl[48] bl[49] bl[50] bl[51] bl[52] bl[53] bl[54] bl[55] bl[56] bl[57] bl[58] bl[59] bl[60] bl[61] bl[62] bl[63] bl[64] bl[65] bl[66] bl[67] bl[68] bl[69] bl[70] bl[71] bl[72] bl[73] bl[74] bl[75] bl[76] bl[77] bl[78] bl[79] bl[80] bl[81] bl[82] bl[83] bl[84] bl[85] bl[86] bl[87] bl[88] bl[89] bl[90] bl[91] bl[92] bl[93] bl[94] bl[95] bl[96] bl[97] bl[98] bl[99] bl[100] bl[101] bl[102] bl[103] bl[104] bl[105] bl[106] bl[107] bl[108] bl[109] bl[110] bl[111] bl[112] bl[113] bl[114] bl[115] bl[116] bl[117] bl[118] bl[119] bl[120] bl[121] bl[122] bl[123] bl[124] bl[125] bl[126] bl[127] bl[128] bl[129] bl[130] bl[131] bl[132] bl[133] bl[134] bl[135] bl[136] bl[137] bl[138] bl[139] bl[140] bl[141] bl[142] bl[143] bl[144] bl[145] bl[146] bl[147] bl[148] bl[149] bl[150] bl[151] bl[152] bl[153] bl[154] bl[155] bl[156] bl[157] bl[158] bl[159] bl[160] bl[161] bl[162] bl[163] bl[164] bl[165] bl[166] bl[167] bl[168] bl[169] bl[170] bl[171] bl[172] bl[173] bl[174] bl[175] bl[176] bl[177] bl[178] bl[179] bl[180] bl[181] bl[182] bl[183] bl[184] bl[185] bl[186] bl[187] bl[188] bl[189] bl[190] bl[191] bl[192] bl[193] bl[194] bl[195] bl[196] bl[197] bl[198] bl[199] bl[200] bl[201] bl[202] bl[203] bl[204] bl[205] bl[206] bl[207] bl[208] bl[209] bl[210] bl[211] bl[212] bl[213] bl[214] bl[215] bl[216] bl[217] bl[218] bl[219] bl[220] bl[221] bl[222] bl[223] bl[224] bl[225] bl[226] bl[227] bl[228] bl[229] bl[230] bl[231] bl[232] bl[233] bl[234] bl[235] bl[236] bl[237] bl[238] bl[239] bl[240] bl[241] bl[242] bl[243] bl[244] bl[245] bl[246] bl[247] bl[248] bl[249] bl[250] bl[251] bl[252] bl[253] bl[254] bl[255] bl[256] bl[257] bl[258] bl[259] bl[260] bl[261] bl[262] bl[263] bl[264] bl[265] bl[266] bl[267] bl[268] bl[269] bl[270] bl[271] bl[272] bl[273] bl[274] bl[275] bl[276] bl[277] bl[278] bl[279] bl[280] bl[281] bl[282] bl[283] bl[284] bl[285] bl[286] bl[287] bl[288] bl[289] bl[290] bl[291] bl[292] bl[293] bl[294] bl[295] bl[296] bl[297] bl[298] bl[299] bl[300] bl[301] bl[302] bl[303] bl[304] bl[305] bl[306] bl[307] bl[308] bl[309] bl[310] bl[311] bl[312] bl[313] bl[314] bl[315] bl[316] bl[317] bl[318] bl[319] bl[320] bl[321] bl[322] bl[323] bl[324] bl[325] bl[326] bl[327] bl[328] bl[329] bl[330] bl[331] bl[332] bl[333] bl[334] bl[335] bl[336] bl[337] bl[338] bl[339] bl[340] bl[341] bl[342] bl[343] bl[344] bl[345] bl[346] bl[347] bl[348] bl[349] bl[350] bl[351] bl[352] bl[353] bl[354] bl[355] bl[356] bl[357] bl[358] bl[359] bl[360] bl[361] bl[362] bl[363] bl[364] bl[365] bl[366] bl[367] bl[368] bl[369] bl[370] bl[371] bl[372] bl[373] bl[374] bl[375] bl[376] bl[377] bl[378] bl[379] bl[380] bl[381] bl[382] bl[383] bl[384] bl[385] bl[386] bl[387] bl[388] bl[389] bl[390] bl[391] bl[392] bl[393] bl[394] bl[395] bl[396] bl[397] bl[398] bl[399] bl[400] bl[401] bl[402] bl[403] bl[404] bl[405] bl[406] bl[407] bl[408] bl[409] bl[410] bl[411] bl[412] bl[413] bl[414] bl[415] bl[416] bl[417] bl[418] bl[419] bl[420] bl[421] bl[422] bl[423] bl[424] bl[425] bl[426] bl[427] bl[428] bl[429] bl[430] bl[431] bl[432] bl[433] bl[434] bl[435] bl[436] bl[437] bl[438] bl[439] bl[440] bl[441] bl[442] bl[443] bl[444] bl[445] bl[446] bl[447] bl[448] bl[449] bl[450] bl[451] bl[452] bl[453] bl[454] bl[455] bl[456] bl[457] bl[458] bl[459] bl[460] bl[461] bl[462] bl[463] bl[464] bl[465] bl[466] bl[467] bl[468] bl[469] bl[470] bl[471] bl[472] bl[473] bl[474] bl[475] bl[476] bl[477] bl[478] bl[479] bl[480] bl[481] bl[482] bl[483] bl[484] bl[485] bl[486] bl[487] bl[488] bl[489] bl[490] bl[491] bl[492] bl[493] bl[494] bl[495] bl[496] bl[497] bl[498] bl[499] bl[500] bl[501] bl[502] bl[503] bl[504] bl[505] bl[506] bl[507] bl[508] bl[509] bl[510] bl[511] br[0] br[1] br[2] br[3] br[4] br[5] br[6] br[7] br[8] br[9] br[10] br[11] br[12] br[13] br[14] br[15] br[16] br[17] br[18] br[19] br[20] br[21] br[22] br[23] br[24] br[25] br[26] br[27] br[28] br[29] br[30] br[31] br[32] br[33] br[34] br[35] br[36] br[37] br[38] br[39] br[40] br[41] br[42] br[43] br[44] br[45] br[46] br[47] br[48] br[49] br[50] br[51] br[52] br[53] br[54] br[55] br[56] br[57] br[58] br[59] br[60] br[61] br[62] br[63] br[64] br[65] br[66] br[67] br[68] br[69] br[70] br[71] br[72] br[73] br[74] br[75] br[76] br[77] br[78] br[79] br[80] br[81] br[82] br[83] br[84] br[85] br[86] br[87] br[88] br[89] br[90] br[91] br[92] br[93] br[94] br[95] br[96] br[97] br[98] br[99] br[100] br[101] br[102] br[103] br[104] br[105] br[106] br[107] br[108] br[109] br[110] br[111] br[112] br[113] br[114] br[115] br[116] br[117] br[118] br[119] br[120] br[121] br[122] br[123] br[124] br[125] br[126] br[127] br[128] br[129] br[130] br[131] br[132] br[133] br[134] br[135] br[136] br[137] br[138] br[139] br[140] br[141] br[142] br[143] br[144] br[145] br[146] br[147] br[148] br[149] br[150] br[151] br[152] br[153] br[154] br[155] br[156] br[157] br[158] br[159] br[160] br[161] br[162] br[163] br[164] br[165] br[166] br[167] br[168] br[169] br[170] br[171] br[172] br[173] br[174] br[175] br[176] br[177] br[178] br[179] br[180] br[181] br[182] br[183] br[184] br[185] br[186] br[187] br[188] br[189] br[190] br[191] br[192] br[193] br[194] br[195] br[196] br[197] br[198] br[199] br[200] br[201] br[202] br[203] br[204] br[205] br[206] br[207] br[208] br[209] br[210] br[211] br[212] br[213] br[214] br[215] br[216] br[217] br[218] br[219] br[220] br[221] br[222] br[223] br[224] br[225] br[226] br[227] br[228] br[229] br[230] br[231] br[232] br[233] br[234] br[235] br[236] br[237] br[238] br[239] br[240] br[241] br[242] br[243] br[244] br[245] br[246] br[247] br[248] br[249] br[250] br[251] br[252] br[253] br[254] br[255] br[256] br[257] br[258] br[259] br[260] br[261] br[262] br[263] br[264] br[265] br[266] br[267] br[268] br[269] br[270] br[271] br[272] br[273] br[274] br[275] br[276] br[277] br[278] br[279] br[280] br[281] br[282] br[283] br[284] br[285] br[286] br[287] br[288] br[289] br[290] br[291] br[292] br[293] br[294] br[295] br[296] br[297] br[298] br[299] br[300] br[301] br[302] br[303] br[304] br[305] br[306] br[307] br[308] br[309] br[310] br[311] br[312] br[313] br[314] br[315] br[316] br[317] br[318] br[319] br[320] br[321] br[322] br[323] br[324] br[325] br[326] br[327] br[328] br[329] br[330] br[331] br[332] br[333] br[334] br[335] br[336] br[337] br[338] br[339] br[340] br[341] br[342] br[343] br[344] br[345] br[346] br[347] br[348] br[349] br[350] br[351] br[352] br[353] br[354] br[355] br[356] br[357] br[358] br[359] br[360] br[361] br[362] br[363] br[364] br[365] br[366] br[367] br[368] br[369] br[370] br[371] br[372] br[373] br[374] br[375] br[376] br[377] br[378] br[379] br[380] br[381] br[382] br[383] br[384] br[385] br[386] br[387] br[388] br[389] br[390] br[391] br[392] br[393] br[394] br[395] br[396] br[397] br[398] br[399] br[400] br[401] br[402] br[403] br[404] br[405] br[406] br[407] br[408] br[409] br[410] br[411] br[412] br[413] br[414] br[415] br[416] br[417] br[418] br[419] br[420] br[421] br[422] br[423] br[424] br[425] br[426] br[427] br[428] br[429] br[430] br[431] br[432] br[433] br[434] br[435] br[436] br[437] br[438] br[439] br[440] br[441] br[442] br[443] br[444] br[445] br[446] br[447] br[448] br[449] br[450] br[451] br[452] br[453] br[454] br[455] br[456] br[457] br[458] br[459] br[460] br[461] br[462] br[463] br[464] br[465] br[466] br[467] br[468] br[469] br[470] br[471] br[472] br[473] br[474] br[475] br[476] br[477] br[478] br[479] br[480] br[481] br[482] br[483] br[484] br[485] br[486] br[487] br[488] br[489] br[490] br[491] br[492] br[493] br[494] br[495] br[496] br[497] br[498] br[499] br[500] br[501] br[502] br[503] br[504] br[505] br[506] br[507] br[508] br[509] br[510] br[511] pc_b col_sel[0] col_sel[1] col_sel[2] col_sel[3] col_sel_b[0] col_sel_b[1] col_sel_b[2] col_sel_b[3] write_driver_en wmask[0] wmask[1] wmask[2] wmask[3] wmask[4] wmask[5] wmask[6] wmask[7] wmask[8] wmask[9] wmask[10] wmask[11] wmask[12] wmask[13] wmask[14] wmask[15] din[0] din[1] din[2] din[3] din[4] din[5] din[6] din[7] din[8] din[9] din[10] din[11] din[12] din[13] din[14] din[15] din[16] din[17] din[18] din[19] din[20] din[21] din[22] din[23] din[24] din[25] din[26] din[27] din[28] din[29] din[30] din[31] din[32] din[33] din[34] din[35] din[36] din[37] din[38] din[39] din[40] din[41] din[42] din[43] din[44] din[45] din[46] din[47] din[48] din[49] din[50] din[51] din[52] din[53] din[54] din[55] din[56] din[57] din[58] din[59] din[60] din[61] din[62] din[63] din[64] din[65] din[66] din[67] din[68] din[69] din[70] din[71] din[72] din[73] din[74] din[75] din[76] din[77] din[78] din[79] din[80] din[81] din[82] din[83] din[84] din[85] din[86] din[87] din[88] din[89] din[90] din[91] din[92] din[93] din[94] din[95] din[96] din[97] din[98] din[99] din[100] din[101] din[102] din[103] din[104] din[105] din[106] din[107] din[108] din[109] din[110] din[111] din[112] din[113] din[114] din[115] din[116] din[117] din[118] din[119] din[120] din[121] din[122] din[123] din[124] din[125] din[126] din[127] dout[0] dout[1] dout[2] dout[3] dout[4] dout[5] dout[6] dout[7] dout[8] dout[9] dout[10] dout[11] dout[12] dout[13] dout[14] dout[15] dout[16] dout[17] dout[18] dout[19] dout[20] dout[21] dout[22] dout[23] dout[24] dout[25] dout[26] dout[27] dout[28] dout[29] dout[30] dout[31] dout[32] dout[33] dout[34] dout[35] dout[36] dout[37] dout[38] dout[39] dout[40] dout[41] dout[42] dout[43] dout[44] dout[45] dout[46] dout[47] dout[48] dout[49] dout[50] dout[51] dout[52] dout[53] dout[54] dout[55] dout[56] dout[57] dout[58] dout[59] dout[60] dout[61] dout[62] dout[63] dout[64] dout[65] dout[66] dout[67] dout[68] dout[69] dout[70] dout[71] dout[72] dout[73] dout[74] dout[75] dout[76] dout[77] dout[78] dout[79] dout[80] dout[81] dout[82] dout[83] dout[84] dout[85] dout[86] dout[87] dout[88] dout[89] dout[90] dout[91] dout[92] dout[93] dout[94] dout[95] dout[96] dout[97] dout[98] dout[99] dout[100] dout[101] dout[102] dout[103] dout[104] dout[105] dout[106] dout[107] dout[108] dout[109] dout[110] dout[111] dout[112] dout[113] dout[114] dout[115] dout[116] dout[117] dout[118] dout[119] dout[120] dout[121] dout[122] dout[123] dout[124] dout[125] dout[126] dout[127] col_peripherals
  Xreplica_precharge_0 vdd rbl rbr pc_b0 precharge
  Xreplica_precharge_1 vdd rbl rbr pc_b0 precharge
  Xreplica_mos vdd vss rbl replica_column_mos

.ENDS sram22_inner

.SUBCKT sram22_256x128m4w8 vdd vss clk we ce rstb addr[0] addr[1] addr[2] addr[3] addr[4] addr[5] addr[6] addr[7] wmask[0] wmask[1] wmask[2] wmask[3] wmask[4] wmask[5] wmask[6] wmask[7] wmask[8] wmask[9] wmask[10] wmask[11] wmask[12] wmask[13] wmask[14] wmask[15] din[0] din[1] din[2] din[3] din[4] din[5] din[6] din[7] din[8] din[9] din[10] din[11] din[12] din[13] din[14] din[15] din[16] din[17] din[18] din[19] din[20] din[21] din[22] din[23] din[24] din[25] din[26] din[27] din[28] din[29] din[30] din[31] din[32] din[33] din[34] din[35] din[36] din[37] din[38] din[39] din[40] din[41] din[42] din[43] din[44] din[45] din[46] din[47] din[48] din[49] din[50] din[51] din[52] din[53] din[54] din[55] din[56] din[57] din[58] din[59] din[60] din[61] din[62] din[63] din[64] din[65] din[66] din[67] din[68] din[69] din[70] din[71] din[72] din[73] din[74] din[75] din[76] din[77] din[78] din[79] din[80] din[81] din[82] din[83] din[84] din[85] din[86] din[87] din[88] din[89] din[90] din[91] din[92] din[93] din[94] din[95] din[96] din[97] din[98] din[99] din[100] din[101] din[102] din[103] din[104] din[105] din[106] din[107] din[108] din[109] din[110] din[111] din[112] din[113] din[114] din[115] din[116] din[117] din[118] din[119] din[120] din[121] din[122] din[123] din[124] din[125] din[126] din[127] dout[0] dout[1] dout[2] dout[3] dout[4] dout[5] dout[6] dout[7] dout[8] dout[9] dout[10] dout[11] dout[12] dout[13] dout[14] dout[15] dout[16] dout[17] dout[18] dout[19] dout[20] dout[21] dout[22] dout[23] dout[24] dout[25] dout[26] dout[27] dout[28] dout[29] dout[30] dout[31] dout[32] dout[33] dout[34] dout[35] dout[36] dout[37] dout[38] dout[39] dout[40] dout[41] dout[42] dout[43] dout[44] dout[45] dout[46] dout[47] dout[48] dout[49] dout[50] dout[51] dout[52] dout[53] dout[54] dout[55] dout[56] dout[57] dout[58] dout[59] dout[60] dout[61] dout[62] dout[63] dout[64] dout[65] dout[66] dout[67] dout[68] dout[69] dout[70] dout[71] dout[72] dout[73] dout[74] dout[75] dout[76] dout[77] dout[78] dout[79] dout[80] dout[81] dout[82] dout[83] dout[84] dout[85] dout[86] dout[87] dout[88] dout[89] dout[90] dout[91] dout[92] dout[93] dout[94] dout[95] dout[96] dout[97] dout[98] dout[99] dout[100] dout[101] dout[102] dout[103] dout[104] dout[105] dout[106] dout[107] dout[108] dout[109] dout[110] dout[111] dout[112] dout[113] dout[114] dout[115] dout[116] dout[117] dout[118] dout[119] dout[120] dout[121] dout[122] dout[123] dout[124] dout[125] dout[126] dout[127]

  X0 vdd vss clk we ce rstb addr[0] addr[1] addr[2] addr[3] addr[4] addr[5] addr[6] addr[7] wmask[0] wmask[1] wmask[2] wmask[3] wmask[4] wmask[5] wmask[6] wmask[7] wmask[8] wmask[9] wmask[10] wmask[11] wmask[12] wmask[13] wmask[14] wmask[15] din[0] din[1] din[2] din[3] din[4] din[5] din[6] din[7] din[8] din[9] din[10] din[11] din[12] din[13] din[14] din[15] din[16] din[17] din[18] din[19] din[20] din[21] din[22] din[23] din[24] din[25] din[26] din[27] din[28] din[29] din[30] din[31] din[32] din[33] din[34] din[35] din[36] din[37] din[38] din[39] din[40] din[41] din[42] din[43] din[44] din[45] din[46] din[47] din[48] din[49] din[50] din[51] din[52] din[53] din[54] din[55] din[56] din[57] din[58] din[59] din[60] din[61] din[62] din[63] din[64] din[65] din[66] din[67] din[68] din[69] din[70] din[71] din[72] din[73] din[74] din[75] din[76] din[77] din[78] din[79] din[80] din[81] din[82] din[83] din[84] din[85] din[86] din[87] din[88] din[89] din[90] din[91] din[92] din[93] din[94] din[95] din[96] din[97] din[98] din[99] din[100] din[101] din[102] din[103] din[104] din[105] din[106] din[107] din[108] din[109] din[110] din[111] din[112] din[113] din[114] din[115] din[116] din[117] din[118] din[119] din[120] din[121] din[122] din[123] din[124] din[125] din[126] din[127] dout[0] dout[1] dout[2] dout[3] dout[4] dout[5] dout[6] dout[7] dout[8] dout[9] dout[10] dout[11] dout[12] dout[13] dout[14] dout[15] dout[16] dout[17] dout[18] dout[19] dout[20] dout[21] dout[22] dout[23] dout[24] dout[25] dout[26] dout[27] dout[28] dout[29] dout[30] dout[31] dout[32] dout[33] dout[34] dout[35] dout[36] dout[37] dout[38] dout[39] dout[40] dout[41] dout[42] dout[43] dout[44] dout[45] dout[46] dout[47] dout[48] dout[49] dout[50] dout[51] dout[52] dout[53] dout[54] dout[55] dout[56] dout[57] dout[58] dout[59] dout[60] dout[61] dout[62] dout[63] dout[64] dout[65] dout[66] dout[67] dout[68] dout[69] dout[70] dout[71] dout[72] dout[73] dout[74] dout[75] dout[76] dout[77] dout[78] dout[79] dout[80] dout[81] dout[82] dout[83] dout[84] dout[85] dout[86] dout[87] dout[88] dout[89] dout[90] dout[91] dout[92] dout[93] dout[94] dout[95] dout[96] dout[97] dout[98] dout[99] dout[100] dout[101] dout[102] dout[103] dout[104] dout[105] dout[106] dout[107] dout[108] dout[109] dout[110] dout[111] dout[112] dout[113] dout[114] dout[115] dout[116] dout[117] dout[118] dout[119] dout[120] dout[121] dout[122] dout[123] dout[124] dout[125] dout[126] dout[127] sram22_inner

.ENDS sram22_256x128m4w8

