* circuit.Package sramgen_sramgen_sram_64x32m4w32_replica_v1
* Written by SpiceNetlister
* 

.SUBCKT hierarchical_decoder_nand_2 
+ gnd vdd a b y 

xn1 
+ x a gnd gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='3.2' l='0.15' 

xn2 
+ y b x gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='3.2' l='0.15' 

xp1 
+ y a vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.4' l='0.15' 

xp2 
+ y b vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.4' l='0.15' 

.ENDS

.SUBCKT hierarchical_decoder_inv_3 
+ gnd vdd din din_b 

xn 
+ din_b din gnd gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='1.6' l='0.15' 

xp 
+ din_b din vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.4' l='0.15' 

.ENDS

.SUBCKT hierarchical_decoder 
+ vdd gnd addr[3] addr[2] addr[1] addr[0] addr_b[3] addr_b[2] addr_b[1] addr_b[0] decode[15] decode[14] decode[13] decode[12] decode[11] decode[10] decode[9] decode[8] decode[7] decode[6] decode[5] decode[4] decode[3] decode[2] decode[1] decode[0] decode_b[15] decode_b[14] decode_b[13] decode_b[12] decode_b[11] decode_b[10] decode_b[9] decode_b[8] decode_b[7] decode_b[6] decode_b[5] decode_b[4] decode_b[3] decode_b[2] decode_b[1] decode_b[0] 

xnand_5 
+ gnd vdd addr_b[3] addr_b[2] net_4 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_6 
+ gnd vdd net_4 predecode_1[0] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_8 
+ gnd vdd addr_b[3] addr[2] net_7 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_9 
+ gnd vdd net_7 predecode_1[1] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_11 
+ gnd vdd addr[3] addr_b[2] net_10 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_12 
+ gnd vdd net_10 predecode_1[2] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_14 
+ gnd vdd addr[3] addr[2] net_13 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_15 
+ gnd vdd net_13 predecode_1[3] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_18 
+ gnd vdd addr_b[1] addr_b[0] net_17 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_19 
+ gnd vdd net_17 predecode_16[0] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_21 
+ gnd vdd addr_b[1] addr[0] net_20 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_22 
+ gnd vdd net_20 predecode_16[1] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_24 
+ gnd vdd addr[1] addr_b[0] net_23 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_25 
+ gnd vdd net_23 predecode_16[2] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_27 
+ gnd vdd addr[1] addr[0] net_26 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_28 
+ gnd vdd net_26 predecode_16[3] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_29 
+ gnd vdd predecode_1[0] predecode_16[0] decode_b[0] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_30 
+ gnd vdd decode_b[0] decode[0] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_31 
+ gnd vdd predecode_1[0] predecode_16[1] decode_b[1] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_32 
+ gnd vdd decode_b[1] decode[1] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_33 
+ gnd vdd predecode_1[0] predecode_16[2] decode_b[2] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_34 
+ gnd vdd decode_b[2] decode[2] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_35 
+ gnd vdd predecode_1[0] predecode_16[3] decode_b[3] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_36 
+ gnd vdd decode_b[3] decode[3] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_37 
+ gnd vdd predecode_1[1] predecode_16[0] decode_b[4] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_38 
+ gnd vdd decode_b[4] decode[4] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_39 
+ gnd vdd predecode_1[1] predecode_16[1] decode_b[5] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_40 
+ gnd vdd decode_b[5] decode[5] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_41 
+ gnd vdd predecode_1[1] predecode_16[2] decode_b[6] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_42 
+ gnd vdd decode_b[6] decode[6] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_43 
+ gnd vdd predecode_1[1] predecode_16[3] decode_b[7] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_44 
+ gnd vdd decode_b[7] decode[7] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_45 
+ gnd vdd predecode_1[2] predecode_16[0] decode_b[8] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_46 
+ gnd vdd decode_b[8] decode[8] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_47 
+ gnd vdd predecode_1[2] predecode_16[1] decode_b[9] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_48 
+ gnd vdd decode_b[9] decode[9] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_49 
+ gnd vdd predecode_1[2] predecode_16[2] decode_b[10] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_50 
+ gnd vdd decode_b[10] decode[10] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_51 
+ gnd vdd predecode_1[2] predecode_16[3] decode_b[11] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_52 
+ gnd vdd decode_b[11] decode[11] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_53 
+ gnd vdd predecode_1[3] predecode_16[0] decode_b[12] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_54 
+ gnd vdd decode_b[12] decode[12] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_55 
+ gnd vdd predecode_1[3] predecode_16[1] decode_b[13] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_56 
+ gnd vdd decode_b[13] decode[13] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_57 
+ gnd vdd predecode_1[3] predecode_16[2] decode_b[14] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_58 
+ gnd vdd decode_b[14] decode[14] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_59 
+ gnd vdd predecode_1[3] predecode_16[3] decode_b[15] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_60 
+ gnd vdd decode_b[15] decode[15] 
+ hierarchical_decoder_inv_3 
* No parameters

.ENDS

.SUBCKT column_decoder_nand_1 
+ gnd vdd a b y 

xn1 
+ x a gnd gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='3.2' l='0.15' 

xn2 
+ y b x gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='3.2' l='0.15' 

xp1 
+ y a vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.4' l='0.15' 

xp2 
+ y b vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.4' l='0.15' 

.ENDS

.SUBCKT column_decoder_inv_2 
+ gnd vdd din din_b 

xn 
+ din_b din gnd gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='1.6' l='0.15' 

xp 
+ din_b din vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.4' l='0.15' 

.ENDS

.SUBCKT column_decoder 
+ vdd gnd addr[1] addr[0] addr_b[1] addr_b[0] decode[3] decode[2] decode[1] decode[0] decode_b[3] decode_b[2] decode_b[1] decode_b[0] 

xnand_3 
+ gnd vdd addr_b[1] addr_b[0] decode_b[0] 
+ column_decoder_nand_1 
* No parameters

xinv_4 
+ gnd vdd decode_b[0] decode[0] 
+ column_decoder_inv_2 
* No parameters

xnand_5 
+ gnd vdd addr_b[1] addr[0] decode_b[1] 
+ column_decoder_nand_1 
* No parameters

xinv_6 
+ gnd vdd decode_b[1] decode[1] 
+ column_decoder_inv_2 
* No parameters

xnand_7 
+ gnd vdd addr[1] addr_b[0] decode_b[2] 
+ column_decoder_nand_1 
* No parameters

xinv_8 
+ gnd vdd decode_b[2] decode[2] 
+ column_decoder_inv_2 
* No parameters

xnand_9 
+ gnd vdd addr[1] addr[0] decode_b[3] 
+ column_decoder_nand_1 
* No parameters

xinv_10 
+ gnd vdd decode_b[3] decode[3] 
+ column_decoder_inv_2 
* No parameters

.ENDS

.SUBCKT wordline_driver_and2_nand 
+ gnd vdd a b y 

xn1 
+ x a gnd gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='3.2' l='0.15' 

xn2 
+ y b x gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='3.2' l='0.15' 

xp1 
+ y a vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.4' l='0.15' 

xp2 
+ y b vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.4' l='0.15' 

.ENDS

.SUBCKT wordline_driver_and2_inv 
+ gnd vdd din din_b 

xn 
+ din_b din gnd gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='1.6' l='0.15' 

xp 
+ din_b din vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.4' l='0.15' 

.ENDS

.SUBCKT wordline_driver_and2 
+ a b y vdd vss 

xnand 
+ vss vdd a b tmp 
+ wordline_driver_and2_nand 
* No parameters

xinv 
+ vss vdd tmp y 
+ wordline_driver_and2_inv 
* No parameters

.ENDS

.SUBCKT wordline_driver 
+ vdd vss din wl_en wl 

xand2 
+ din wl_en wl vdd vss 
+ wordline_driver_and2 
* No parameters

.ENDS

.SUBCKT wordline_driver_array 
+ vdd vss din[15] din[14] din[13] din[12] din[11] din[10] din[9] din[8] din[7] din[6] din[5] din[4] din[3] din[2] din[1] din[0] wl_en wl[15] wl[14] wl[13] wl[12] wl[11] wl[10] wl[9] wl[8] wl[7] wl[6] wl[5] wl[4] wl[3] wl[2] wl[1] wl[0] 

xwl_driver_0 
+ vdd vss din[0] wl_en wl[0] 
+ wordline_driver 
* No parameters

xwl_driver_1 
+ vdd vss din[1] wl_en wl[1] 
+ wordline_driver 
* No parameters

xwl_driver_2 
+ vdd vss din[2] wl_en wl[2] 
+ wordline_driver 
* No parameters

xwl_driver_3 
+ vdd vss din[3] wl_en wl[3] 
+ wordline_driver 
* No parameters

xwl_driver_4 
+ vdd vss din[4] wl_en wl[4] 
+ wordline_driver 
* No parameters

xwl_driver_5 
+ vdd vss din[5] wl_en wl[5] 
+ wordline_driver 
* No parameters

xwl_driver_6 
+ vdd vss din[6] wl_en wl[6] 
+ wordline_driver 
* No parameters

xwl_driver_7 
+ vdd vss din[7] wl_en wl[7] 
+ wordline_driver 
* No parameters

xwl_driver_8 
+ vdd vss din[8] wl_en wl[8] 
+ wordline_driver 
* No parameters

xwl_driver_9 
+ vdd vss din[9] wl_en wl[9] 
+ wordline_driver 
* No parameters

xwl_driver_10 
+ vdd vss din[10] wl_en wl[10] 
+ wordline_driver 
* No parameters

xwl_driver_11 
+ vdd vss din[11] wl_en wl[11] 
+ wordline_driver 
* No parameters

xwl_driver_12 
+ vdd vss din[12] wl_en wl[12] 
+ wordline_driver 
* No parameters

xwl_driver_13 
+ vdd vss din[13] wl_en wl[13] 
+ wordline_driver 
* No parameters

xwl_driver_14 
+ vdd vss din[14] wl_en wl[14] 
+ wordline_driver 
* No parameters

xwl_driver_15 
+ vdd vss din[15] wl_en wl[15] 
+ wordline_driver 
* No parameters

.ENDS

.SUBCKT bitcell_array 
+ vdd vss bl[127] bl[126] bl[125] bl[124] bl[123] bl[122] bl[121] bl[120] bl[119] bl[118] bl[117] bl[116] bl[115] bl[114] bl[113] bl[112] bl[111] bl[110] bl[109] bl[108] bl[107] bl[106] bl[105] bl[104] bl[103] bl[102] bl[101] bl[100] bl[99] bl[98] bl[97] bl[96] bl[95] bl[94] bl[93] bl[92] bl[91] bl[90] bl[89] bl[88] bl[87] bl[86] bl[85] bl[84] bl[83] bl[82] bl[81] bl[80] bl[79] bl[78] bl[77] bl[76] bl[75] bl[74] bl[73] bl[72] bl[71] bl[70] bl[69] bl[68] bl[67] bl[66] bl[65] bl[64] bl[63] bl[62] bl[61] bl[60] bl[59] bl[58] bl[57] bl[56] bl[55] bl[54] bl[53] bl[52] bl[51] bl[50] bl[49] bl[48] bl[47] bl[46] bl[45] bl[44] bl[43] bl[42] bl[41] bl[40] bl[39] bl[38] bl[37] bl[36] bl[35] bl[34] bl[33] bl[32] bl[31] bl[30] bl[29] bl[28] bl[27] bl[26] bl[25] bl[24] bl[23] bl[22] bl[21] bl[20] bl[19] bl[18] bl[17] bl[16] bl[15] bl[14] bl[13] bl[12] bl[11] bl[10] bl[9] bl[8] bl[7] bl[6] bl[5] bl[4] bl[3] bl[2] bl[1] bl[0] br[127] br[126] br[125] br[124] br[123] br[122] br[121] br[120] br[119] br[118] br[117] br[116] br[115] br[114] br[113] br[112] br[111] br[110] br[109] br[108] br[107] br[106] br[105] br[104] br[103] br[102] br[101] br[100] br[99] br[98] br[97] br[96] br[95] br[94] br[93] br[92] br[91] br[90] br[89] br[88] br[87] br[86] br[85] br[84] br[83] br[82] br[81] br[80] br[79] br[78] br[77] br[76] br[75] br[74] br[73] br[72] br[71] br[70] br[69] br[68] br[67] br[66] br[65] br[64] br[63] br[62] br[61] br[60] br[59] br[58] br[57] br[56] br[55] br[54] br[53] br[52] br[51] br[50] br[49] br[48] br[47] br[46] br[45] br[44] br[43] br[42] br[41] br[40] br[39] br[38] br[37] br[36] br[35] br[34] br[33] br[32] br[31] br[30] br[29] br[28] br[27] br[26] br[25] br[24] br[23] br[22] br[21] br[20] br[19] br[18] br[17] br[16] br[15] br[14] br[13] br[12] br[11] br[10] br[9] br[8] br[7] br[6] br[5] br[4] br[3] br[2] br[1] br[0] wl[15] wl[14] wl[13] wl[12] wl[11] wl[10] wl[9] wl[8] wl[7] wl[6] wl[5] wl[4] wl[3] wl[2] wl[1] wl[0] vnb vpb rbl rbr 

xbitcell_0_0 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_1 
+ rbl rbr vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_2 
+ bl[0] br[0] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_3 
+ bl[1] br[1] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_4 
+ bl[2] br[2] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_5 
+ bl[3] br[3] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_6 
+ bl[4] br[4] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_7 
+ bl[5] br[5] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_8 
+ bl[6] br[6] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_9 
+ bl[7] br[7] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_10 
+ bl[8] br[8] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_11 
+ bl[9] br[9] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_12 
+ bl[10] br[10] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_13 
+ bl[11] br[11] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_14 
+ bl[12] br[12] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_15 
+ bl[13] br[13] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_16 
+ bl[14] br[14] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_17 
+ bl[15] br[15] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_18 
+ bl[16] br[16] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_19 
+ bl[17] br[17] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_20 
+ bl[18] br[18] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_21 
+ bl[19] br[19] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_22 
+ bl[20] br[20] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_23 
+ bl[21] br[21] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_24 
+ bl[22] br[22] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_25 
+ bl[23] br[23] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_26 
+ bl[24] br[24] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_27 
+ bl[25] br[25] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_28 
+ bl[26] br[26] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_29 
+ bl[27] br[27] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_30 
+ bl[28] br[28] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_31 
+ bl[29] br[29] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_32 
+ bl[30] br[30] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_33 
+ bl[31] br[31] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_34 
+ bl[32] br[32] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_35 
+ bl[33] br[33] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_36 
+ bl[34] br[34] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_37 
+ bl[35] br[35] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_38 
+ bl[36] br[36] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_39 
+ bl[37] br[37] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_40 
+ bl[38] br[38] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_41 
+ bl[39] br[39] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_42 
+ bl[40] br[40] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_43 
+ bl[41] br[41] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_44 
+ bl[42] br[42] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_45 
+ bl[43] br[43] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_46 
+ bl[44] br[44] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_47 
+ bl[45] br[45] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_48 
+ bl[46] br[46] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_49 
+ bl[47] br[47] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_50 
+ bl[48] br[48] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_51 
+ bl[49] br[49] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_52 
+ bl[50] br[50] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_53 
+ bl[51] br[51] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_54 
+ bl[52] br[52] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_55 
+ bl[53] br[53] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_56 
+ bl[54] br[54] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_57 
+ bl[55] br[55] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_58 
+ bl[56] br[56] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_59 
+ bl[57] br[57] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_60 
+ bl[58] br[58] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_61 
+ bl[59] br[59] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_62 
+ bl[60] br[60] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_63 
+ bl[61] br[61] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_64 
+ bl[62] br[62] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_65 
+ bl[63] br[63] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_66 
+ bl[64] br[64] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_67 
+ bl[65] br[65] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_68 
+ bl[66] br[66] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_69 
+ bl[67] br[67] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_70 
+ bl[68] br[68] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_71 
+ bl[69] br[69] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_72 
+ bl[70] br[70] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_73 
+ bl[71] br[71] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_74 
+ bl[72] br[72] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_75 
+ bl[73] br[73] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_76 
+ bl[74] br[74] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_77 
+ bl[75] br[75] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_78 
+ bl[76] br[76] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_79 
+ bl[77] br[77] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_80 
+ bl[78] br[78] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_81 
+ bl[79] br[79] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_82 
+ bl[80] br[80] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_83 
+ bl[81] br[81] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_84 
+ bl[82] br[82] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_85 
+ bl[83] br[83] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_86 
+ bl[84] br[84] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_87 
+ bl[85] br[85] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_88 
+ bl[86] br[86] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_89 
+ bl[87] br[87] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_90 
+ bl[88] br[88] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_91 
+ bl[89] br[89] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_92 
+ bl[90] br[90] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_93 
+ bl[91] br[91] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_94 
+ bl[92] br[92] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_95 
+ bl[93] br[93] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_96 
+ bl[94] br[94] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_97 
+ bl[95] br[95] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_98 
+ bl[96] br[96] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_99 
+ bl[97] br[97] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_100 
+ bl[98] br[98] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_101 
+ bl[99] br[99] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_102 
+ bl[100] br[100] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_103 
+ bl[101] br[101] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_104 
+ bl[102] br[102] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_105 
+ bl[103] br[103] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_106 
+ bl[104] br[104] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_107 
+ bl[105] br[105] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_108 
+ bl[106] br[106] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_109 
+ bl[107] br[107] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_110 
+ bl[108] br[108] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_111 
+ bl[109] br[109] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_112 
+ bl[110] br[110] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_113 
+ bl[111] br[111] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_114 
+ bl[112] br[112] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_115 
+ bl[113] br[113] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_116 
+ bl[114] br[114] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_117 
+ bl[115] br[115] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_118 
+ bl[116] br[116] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_119 
+ bl[117] br[117] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_120 
+ bl[118] br[118] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_121 
+ bl[119] br[119] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_122 
+ bl[120] br[120] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_123 
+ bl[121] br[121] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_124 
+ bl[122] br[122] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_125 
+ bl[123] br[123] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_126 
+ bl[124] br[124] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_127 
+ bl[125] br[125] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_128 
+ bl[126] br[126] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_129 
+ bl[127] br[127] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_130 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_131 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_0 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_1 
+ rbl rbr vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_2 
+ bl[0] br[0] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_3 
+ bl[1] br[1] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_4 
+ bl[2] br[2] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_5 
+ bl[3] br[3] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_6 
+ bl[4] br[4] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_7 
+ bl[5] br[5] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_8 
+ bl[6] br[6] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_9 
+ bl[7] br[7] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_10 
+ bl[8] br[8] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_11 
+ bl[9] br[9] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_12 
+ bl[10] br[10] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_13 
+ bl[11] br[11] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_14 
+ bl[12] br[12] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_15 
+ bl[13] br[13] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_16 
+ bl[14] br[14] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_17 
+ bl[15] br[15] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_18 
+ bl[16] br[16] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_19 
+ bl[17] br[17] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_20 
+ bl[18] br[18] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_21 
+ bl[19] br[19] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_22 
+ bl[20] br[20] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_23 
+ bl[21] br[21] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_24 
+ bl[22] br[22] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_25 
+ bl[23] br[23] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_26 
+ bl[24] br[24] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_27 
+ bl[25] br[25] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_28 
+ bl[26] br[26] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_29 
+ bl[27] br[27] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_30 
+ bl[28] br[28] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_31 
+ bl[29] br[29] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_32 
+ bl[30] br[30] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_33 
+ bl[31] br[31] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_34 
+ bl[32] br[32] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_35 
+ bl[33] br[33] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_36 
+ bl[34] br[34] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_37 
+ bl[35] br[35] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_38 
+ bl[36] br[36] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_39 
+ bl[37] br[37] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_40 
+ bl[38] br[38] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_41 
+ bl[39] br[39] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_42 
+ bl[40] br[40] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_43 
+ bl[41] br[41] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_44 
+ bl[42] br[42] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_45 
+ bl[43] br[43] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_46 
+ bl[44] br[44] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_47 
+ bl[45] br[45] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_48 
+ bl[46] br[46] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_49 
+ bl[47] br[47] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_50 
+ bl[48] br[48] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_51 
+ bl[49] br[49] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_52 
+ bl[50] br[50] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_53 
+ bl[51] br[51] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_54 
+ bl[52] br[52] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_55 
+ bl[53] br[53] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_56 
+ bl[54] br[54] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_57 
+ bl[55] br[55] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_58 
+ bl[56] br[56] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_59 
+ bl[57] br[57] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_60 
+ bl[58] br[58] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_61 
+ bl[59] br[59] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_62 
+ bl[60] br[60] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_63 
+ bl[61] br[61] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_64 
+ bl[62] br[62] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_65 
+ bl[63] br[63] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_66 
+ bl[64] br[64] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_67 
+ bl[65] br[65] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_68 
+ bl[66] br[66] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_69 
+ bl[67] br[67] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_70 
+ bl[68] br[68] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_71 
+ bl[69] br[69] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_72 
+ bl[70] br[70] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_73 
+ bl[71] br[71] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_74 
+ bl[72] br[72] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_75 
+ bl[73] br[73] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_76 
+ bl[74] br[74] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_77 
+ bl[75] br[75] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_78 
+ bl[76] br[76] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_79 
+ bl[77] br[77] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_80 
+ bl[78] br[78] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_81 
+ bl[79] br[79] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_82 
+ bl[80] br[80] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_83 
+ bl[81] br[81] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_84 
+ bl[82] br[82] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_85 
+ bl[83] br[83] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_86 
+ bl[84] br[84] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_87 
+ bl[85] br[85] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_88 
+ bl[86] br[86] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_89 
+ bl[87] br[87] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_90 
+ bl[88] br[88] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_91 
+ bl[89] br[89] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_92 
+ bl[90] br[90] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_93 
+ bl[91] br[91] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_94 
+ bl[92] br[92] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_95 
+ bl[93] br[93] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_96 
+ bl[94] br[94] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_97 
+ bl[95] br[95] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_98 
+ bl[96] br[96] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_99 
+ bl[97] br[97] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_100 
+ bl[98] br[98] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_101 
+ bl[99] br[99] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_102 
+ bl[100] br[100] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_103 
+ bl[101] br[101] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_104 
+ bl[102] br[102] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_105 
+ bl[103] br[103] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_106 
+ bl[104] br[104] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_107 
+ bl[105] br[105] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_108 
+ bl[106] br[106] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_109 
+ bl[107] br[107] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_110 
+ bl[108] br[108] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_111 
+ bl[109] br[109] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_112 
+ bl[110] br[110] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_113 
+ bl[111] br[111] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_114 
+ bl[112] br[112] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_115 
+ bl[113] br[113] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_116 
+ bl[114] br[114] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_117 
+ bl[115] br[115] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_118 
+ bl[116] br[116] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_119 
+ bl[117] br[117] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_120 
+ bl[118] br[118] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_121 
+ bl[119] br[119] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_122 
+ bl[120] br[120] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_123 
+ bl[121] br[121] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_124 
+ bl[122] br[122] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_125 
+ bl[123] br[123] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_126 
+ bl[124] br[124] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_127 
+ bl[125] br[125] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_128 
+ bl[126] br[126] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_129 
+ bl[127] br[127] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_130 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_131 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_0 
+ vdd vdd vss vdd vpb vnb wl[0] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_2_1 
+ rbl rbr vss vdd vpb vnb wl[0] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_2_2 
+ bl[0] br[0] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_3 
+ bl[1] br[1] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_4 
+ bl[2] br[2] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_5 
+ bl[3] br[3] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_6 
+ bl[4] br[4] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_7 
+ bl[5] br[5] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_8 
+ bl[6] br[6] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_9 
+ bl[7] br[7] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_10 
+ bl[8] br[8] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_11 
+ bl[9] br[9] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_12 
+ bl[10] br[10] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_13 
+ bl[11] br[11] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_14 
+ bl[12] br[12] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_15 
+ bl[13] br[13] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_16 
+ bl[14] br[14] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_17 
+ bl[15] br[15] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_18 
+ bl[16] br[16] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_19 
+ bl[17] br[17] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_20 
+ bl[18] br[18] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_21 
+ bl[19] br[19] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_22 
+ bl[20] br[20] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_23 
+ bl[21] br[21] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_24 
+ bl[22] br[22] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_25 
+ bl[23] br[23] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_26 
+ bl[24] br[24] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_27 
+ bl[25] br[25] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_28 
+ bl[26] br[26] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_29 
+ bl[27] br[27] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_30 
+ bl[28] br[28] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_31 
+ bl[29] br[29] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_32 
+ bl[30] br[30] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_33 
+ bl[31] br[31] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_34 
+ bl[32] br[32] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_35 
+ bl[33] br[33] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_36 
+ bl[34] br[34] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_37 
+ bl[35] br[35] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_38 
+ bl[36] br[36] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_39 
+ bl[37] br[37] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_40 
+ bl[38] br[38] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_41 
+ bl[39] br[39] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_42 
+ bl[40] br[40] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_43 
+ bl[41] br[41] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_44 
+ bl[42] br[42] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_45 
+ bl[43] br[43] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_46 
+ bl[44] br[44] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_47 
+ bl[45] br[45] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_48 
+ bl[46] br[46] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_49 
+ bl[47] br[47] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_50 
+ bl[48] br[48] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_51 
+ bl[49] br[49] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_52 
+ bl[50] br[50] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_53 
+ bl[51] br[51] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_54 
+ bl[52] br[52] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_55 
+ bl[53] br[53] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_56 
+ bl[54] br[54] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_57 
+ bl[55] br[55] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_58 
+ bl[56] br[56] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_59 
+ bl[57] br[57] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_60 
+ bl[58] br[58] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_61 
+ bl[59] br[59] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_62 
+ bl[60] br[60] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_63 
+ bl[61] br[61] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_64 
+ bl[62] br[62] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_65 
+ bl[63] br[63] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_66 
+ bl[64] br[64] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_67 
+ bl[65] br[65] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_68 
+ bl[66] br[66] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_69 
+ bl[67] br[67] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_70 
+ bl[68] br[68] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_71 
+ bl[69] br[69] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_72 
+ bl[70] br[70] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_73 
+ bl[71] br[71] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_74 
+ bl[72] br[72] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_75 
+ bl[73] br[73] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_76 
+ bl[74] br[74] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_77 
+ bl[75] br[75] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_78 
+ bl[76] br[76] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_79 
+ bl[77] br[77] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_80 
+ bl[78] br[78] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_81 
+ bl[79] br[79] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_82 
+ bl[80] br[80] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_83 
+ bl[81] br[81] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_84 
+ bl[82] br[82] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_85 
+ bl[83] br[83] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_86 
+ bl[84] br[84] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_87 
+ bl[85] br[85] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_88 
+ bl[86] br[86] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_89 
+ bl[87] br[87] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_90 
+ bl[88] br[88] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_91 
+ bl[89] br[89] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_92 
+ bl[90] br[90] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_93 
+ bl[91] br[91] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_94 
+ bl[92] br[92] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_95 
+ bl[93] br[93] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_96 
+ bl[94] br[94] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_97 
+ bl[95] br[95] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_98 
+ bl[96] br[96] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_99 
+ bl[97] br[97] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_100 
+ bl[98] br[98] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_101 
+ bl[99] br[99] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_102 
+ bl[100] br[100] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_103 
+ bl[101] br[101] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_104 
+ bl[102] br[102] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_105 
+ bl[103] br[103] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_106 
+ bl[104] br[104] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_107 
+ bl[105] br[105] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_108 
+ bl[106] br[106] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_109 
+ bl[107] br[107] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_110 
+ bl[108] br[108] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_111 
+ bl[109] br[109] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_112 
+ bl[110] br[110] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_113 
+ bl[111] br[111] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_114 
+ bl[112] br[112] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_115 
+ bl[113] br[113] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_116 
+ bl[114] br[114] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_117 
+ bl[115] br[115] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_118 
+ bl[116] br[116] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_119 
+ bl[117] br[117] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_120 
+ bl[118] br[118] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_121 
+ bl[119] br[119] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_122 
+ bl[120] br[120] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_123 
+ bl[121] br[121] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_124 
+ bl[122] br[122] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_125 
+ bl[123] br[123] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_126 
+ bl[124] br[124] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_127 
+ bl[125] br[125] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_128 
+ bl[126] br[126] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_129 
+ bl[127] br[127] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_130 
+ vdd vdd vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_131 
+ vdd vdd vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_0 
+ vdd vdd vss vdd vpb vnb wl[1] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_3_1 
+ rbl rbr vss vdd vpb vnb wl[1] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_3_2 
+ bl[0] br[0] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_3 
+ bl[1] br[1] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_4 
+ bl[2] br[2] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_5 
+ bl[3] br[3] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_6 
+ bl[4] br[4] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_7 
+ bl[5] br[5] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_8 
+ bl[6] br[6] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_9 
+ bl[7] br[7] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_10 
+ bl[8] br[8] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_11 
+ bl[9] br[9] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_12 
+ bl[10] br[10] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_13 
+ bl[11] br[11] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_14 
+ bl[12] br[12] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_15 
+ bl[13] br[13] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_16 
+ bl[14] br[14] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_17 
+ bl[15] br[15] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_18 
+ bl[16] br[16] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_19 
+ bl[17] br[17] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_20 
+ bl[18] br[18] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_21 
+ bl[19] br[19] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_22 
+ bl[20] br[20] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_23 
+ bl[21] br[21] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_24 
+ bl[22] br[22] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_25 
+ bl[23] br[23] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_26 
+ bl[24] br[24] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_27 
+ bl[25] br[25] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_28 
+ bl[26] br[26] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_29 
+ bl[27] br[27] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_30 
+ bl[28] br[28] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_31 
+ bl[29] br[29] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_32 
+ bl[30] br[30] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_33 
+ bl[31] br[31] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_34 
+ bl[32] br[32] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_35 
+ bl[33] br[33] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_36 
+ bl[34] br[34] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_37 
+ bl[35] br[35] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_38 
+ bl[36] br[36] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_39 
+ bl[37] br[37] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_40 
+ bl[38] br[38] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_41 
+ bl[39] br[39] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_42 
+ bl[40] br[40] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_43 
+ bl[41] br[41] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_44 
+ bl[42] br[42] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_45 
+ bl[43] br[43] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_46 
+ bl[44] br[44] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_47 
+ bl[45] br[45] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_48 
+ bl[46] br[46] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_49 
+ bl[47] br[47] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_50 
+ bl[48] br[48] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_51 
+ bl[49] br[49] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_52 
+ bl[50] br[50] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_53 
+ bl[51] br[51] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_54 
+ bl[52] br[52] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_55 
+ bl[53] br[53] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_56 
+ bl[54] br[54] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_57 
+ bl[55] br[55] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_58 
+ bl[56] br[56] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_59 
+ bl[57] br[57] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_60 
+ bl[58] br[58] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_61 
+ bl[59] br[59] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_62 
+ bl[60] br[60] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_63 
+ bl[61] br[61] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_64 
+ bl[62] br[62] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_65 
+ bl[63] br[63] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_66 
+ bl[64] br[64] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_67 
+ bl[65] br[65] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_68 
+ bl[66] br[66] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_69 
+ bl[67] br[67] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_70 
+ bl[68] br[68] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_71 
+ bl[69] br[69] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_72 
+ bl[70] br[70] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_73 
+ bl[71] br[71] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_74 
+ bl[72] br[72] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_75 
+ bl[73] br[73] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_76 
+ bl[74] br[74] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_77 
+ bl[75] br[75] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_78 
+ bl[76] br[76] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_79 
+ bl[77] br[77] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_80 
+ bl[78] br[78] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_81 
+ bl[79] br[79] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_82 
+ bl[80] br[80] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_83 
+ bl[81] br[81] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_84 
+ bl[82] br[82] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_85 
+ bl[83] br[83] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_86 
+ bl[84] br[84] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_87 
+ bl[85] br[85] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_88 
+ bl[86] br[86] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_89 
+ bl[87] br[87] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_90 
+ bl[88] br[88] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_91 
+ bl[89] br[89] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_92 
+ bl[90] br[90] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_93 
+ bl[91] br[91] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_94 
+ bl[92] br[92] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_95 
+ bl[93] br[93] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_96 
+ bl[94] br[94] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_97 
+ bl[95] br[95] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_98 
+ bl[96] br[96] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_99 
+ bl[97] br[97] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_100 
+ bl[98] br[98] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_101 
+ bl[99] br[99] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_102 
+ bl[100] br[100] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_103 
+ bl[101] br[101] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_104 
+ bl[102] br[102] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_105 
+ bl[103] br[103] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_106 
+ bl[104] br[104] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_107 
+ bl[105] br[105] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_108 
+ bl[106] br[106] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_109 
+ bl[107] br[107] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_110 
+ bl[108] br[108] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_111 
+ bl[109] br[109] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_112 
+ bl[110] br[110] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_113 
+ bl[111] br[111] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_114 
+ bl[112] br[112] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_115 
+ bl[113] br[113] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_116 
+ bl[114] br[114] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_117 
+ bl[115] br[115] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_118 
+ bl[116] br[116] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_119 
+ bl[117] br[117] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_120 
+ bl[118] br[118] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_121 
+ bl[119] br[119] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_122 
+ bl[120] br[120] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_123 
+ bl[121] br[121] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_124 
+ bl[122] br[122] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_125 
+ bl[123] br[123] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_126 
+ bl[124] br[124] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_127 
+ bl[125] br[125] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_128 
+ bl[126] br[126] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_129 
+ bl[127] br[127] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_130 
+ vdd vdd vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_131 
+ vdd vdd vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_0 
+ vdd vdd vss vdd vpb vnb wl[2] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_4_1 
+ rbl rbr vss vdd vpb vnb wl[2] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_4_2 
+ bl[0] br[0] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_3 
+ bl[1] br[1] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_4 
+ bl[2] br[2] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_5 
+ bl[3] br[3] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_6 
+ bl[4] br[4] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_7 
+ bl[5] br[5] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_8 
+ bl[6] br[6] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_9 
+ bl[7] br[7] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_10 
+ bl[8] br[8] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_11 
+ bl[9] br[9] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_12 
+ bl[10] br[10] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_13 
+ bl[11] br[11] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_14 
+ bl[12] br[12] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_15 
+ bl[13] br[13] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_16 
+ bl[14] br[14] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_17 
+ bl[15] br[15] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_18 
+ bl[16] br[16] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_19 
+ bl[17] br[17] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_20 
+ bl[18] br[18] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_21 
+ bl[19] br[19] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_22 
+ bl[20] br[20] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_23 
+ bl[21] br[21] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_24 
+ bl[22] br[22] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_25 
+ bl[23] br[23] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_26 
+ bl[24] br[24] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_27 
+ bl[25] br[25] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_28 
+ bl[26] br[26] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_29 
+ bl[27] br[27] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_30 
+ bl[28] br[28] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_31 
+ bl[29] br[29] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_32 
+ bl[30] br[30] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_33 
+ bl[31] br[31] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_34 
+ bl[32] br[32] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_35 
+ bl[33] br[33] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_36 
+ bl[34] br[34] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_37 
+ bl[35] br[35] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_38 
+ bl[36] br[36] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_39 
+ bl[37] br[37] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_40 
+ bl[38] br[38] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_41 
+ bl[39] br[39] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_42 
+ bl[40] br[40] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_43 
+ bl[41] br[41] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_44 
+ bl[42] br[42] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_45 
+ bl[43] br[43] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_46 
+ bl[44] br[44] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_47 
+ bl[45] br[45] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_48 
+ bl[46] br[46] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_49 
+ bl[47] br[47] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_50 
+ bl[48] br[48] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_51 
+ bl[49] br[49] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_52 
+ bl[50] br[50] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_53 
+ bl[51] br[51] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_54 
+ bl[52] br[52] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_55 
+ bl[53] br[53] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_56 
+ bl[54] br[54] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_57 
+ bl[55] br[55] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_58 
+ bl[56] br[56] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_59 
+ bl[57] br[57] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_60 
+ bl[58] br[58] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_61 
+ bl[59] br[59] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_62 
+ bl[60] br[60] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_63 
+ bl[61] br[61] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_64 
+ bl[62] br[62] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_65 
+ bl[63] br[63] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_66 
+ bl[64] br[64] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_67 
+ bl[65] br[65] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_68 
+ bl[66] br[66] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_69 
+ bl[67] br[67] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_70 
+ bl[68] br[68] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_71 
+ bl[69] br[69] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_72 
+ bl[70] br[70] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_73 
+ bl[71] br[71] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_74 
+ bl[72] br[72] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_75 
+ bl[73] br[73] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_76 
+ bl[74] br[74] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_77 
+ bl[75] br[75] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_78 
+ bl[76] br[76] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_79 
+ bl[77] br[77] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_80 
+ bl[78] br[78] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_81 
+ bl[79] br[79] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_82 
+ bl[80] br[80] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_83 
+ bl[81] br[81] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_84 
+ bl[82] br[82] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_85 
+ bl[83] br[83] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_86 
+ bl[84] br[84] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_87 
+ bl[85] br[85] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_88 
+ bl[86] br[86] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_89 
+ bl[87] br[87] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_90 
+ bl[88] br[88] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_91 
+ bl[89] br[89] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_92 
+ bl[90] br[90] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_93 
+ bl[91] br[91] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_94 
+ bl[92] br[92] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_95 
+ bl[93] br[93] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_96 
+ bl[94] br[94] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_97 
+ bl[95] br[95] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_98 
+ bl[96] br[96] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_99 
+ bl[97] br[97] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_100 
+ bl[98] br[98] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_101 
+ bl[99] br[99] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_102 
+ bl[100] br[100] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_103 
+ bl[101] br[101] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_104 
+ bl[102] br[102] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_105 
+ bl[103] br[103] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_106 
+ bl[104] br[104] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_107 
+ bl[105] br[105] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_108 
+ bl[106] br[106] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_109 
+ bl[107] br[107] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_110 
+ bl[108] br[108] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_111 
+ bl[109] br[109] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_112 
+ bl[110] br[110] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_113 
+ bl[111] br[111] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_114 
+ bl[112] br[112] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_115 
+ bl[113] br[113] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_116 
+ bl[114] br[114] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_117 
+ bl[115] br[115] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_118 
+ bl[116] br[116] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_119 
+ bl[117] br[117] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_120 
+ bl[118] br[118] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_121 
+ bl[119] br[119] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_122 
+ bl[120] br[120] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_123 
+ bl[121] br[121] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_124 
+ bl[122] br[122] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_125 
+ bl[123] br[123] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_126 
+ bl[124] br[124] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_127 
+ bl[125] br[125] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_128 
+ bl[126] br[126] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_129 
+ bl[127] br[127] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_130 
+ vdd vdd vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_131 
+ vdd vdd vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_0 
+ vdd vdd vss vdd vpb vnb wl[3] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_5_1 
+ rbl rbr vss vdd vpb vnb wl[3] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_5_2 
+ bl[0] br[0] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_3 
+ bl[1] br[1] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_4 
+ bl[2] br[2] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_5 
+ bl[3] br[3] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_6 
+ bl[4] br[4] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_7 
+ bl[5] br[5] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_8 
+ bl[6] br[6] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_9 
+ bl[7] br[7] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_10 
+ bl[8] br[8] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_11 
+ bl[9] br[9] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_12 
+ bl[10] br[10] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_13 
+ bl[11] br[11] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_14 
+ bl[12] br[12] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_15 
+ bl[13] br[13] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_16 
+ bl[14] br[14] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_17 
+ bl[15] br[15] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_18 
+ bl[16] br[16] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_19 
+ bl[17] br[17] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_20 
+ bl[18] br[18] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_21 
+ bl[19] br[19] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_22 
+ bl[20] br[20] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_23 
+ bl[21] br[21] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_24 
+ bl[22] br[22] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_25 
+ bl[23] br[23] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_26 
+ bl[24] br[24] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_27 
+ bl[25] br[25] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_28 
+ bl[26] br[26] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_29 
+ bl[27] br[27] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_30 
+ bl[28] br[28] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_31 
+ bl[29] br[29] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_32 
+ bl[30] br[30] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_33 
+ bl[31] br[31] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_34 
+ bl[32] br[32] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_35 
+ bl[33] br[33] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_36 
+ bl[34] br[34] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_37 
+ bl[35] br[35] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_38 
+ bl[36] br[36] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_39 
+ bl[37] br[37] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_40 
+ bl[38] br[38] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_41 
+ bl[39] br[39] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_42 
+ bl[40] br[40] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_43 
+ bl[41] br[41] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_44 
+ bl[42] br[42] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_45 
+ bl[43] br[43] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_46 
+ bl[44] br[44] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_47 
+ bl[45] br[45] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_48 
+ bl[46] br[46] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_49 
+ bl[47] br[47] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_50 
+ bl[48] br[48] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_51 
+ bl[49] br[49] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_52 
+ bl[50] br[50] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_53 
+ bl[51] br[51] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_54 
+ bl[52] br[52] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_55 
+ bl[53] br[53] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_56 
+ bl[54] br[54] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_57 
+ bl[55] br[55] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_58 
+ bl[56] br[56] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_59 
+ bl[57] br[57] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_60 
+ bl[58] br[58] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_61 
+ bl[59] br[59] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_62 
+ bl[60] br[60] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_63 
+ bl[61] br[61] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_64 
+ bl[62] br[62] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_65 
+ bl[63] br[63] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_66 
+ bl[64] br[64] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_67 
+ bl[65] br[65] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_68 
+ bl[66] br[66] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_69 
+ bl[67] br[67] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_70 
+ bl[68] br[68] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_71 
+ bl[69] br[69] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_72 
+ bl[70] br[70] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_73 
+ bl[71] br[71] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_74 
+ bl[72] br[72] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_75 
+ bl[73] br[73] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_76 
+ bl[74] br[74] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_77 
+ bl[75] br[75] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_78 
+ bl[76] br[76] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_79 
+ bl[77] br[77] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_80 
+ bl[78] br[78] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_81 
+ bl[79] br[79] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_82 
+ bl[80] br[80] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_83 
+ bl[81] br[81] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_84 
+ bl[82] br[82] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_85 
+ bl[83] br[83] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_86 
+ bl[84] br[84] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_87 
+ bl[85] br[85] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_88 
+ bl[86] br[86] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_89 
+ bl[87] br[87] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_90 
+ bl[88] br[88] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_91 
+ bl[89] br[89] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_92 
+ bl[90] br[90] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_93 
+ bl[91] br[91] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_94 
+ bl[92] br[92] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_95 
+ bl[93] br[93] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_96 
+ bl[94] br[94] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_97 
+ bl[95] br[95] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_98 
+ bl[96] br[96] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_99 
+ bl[97] br[97] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_100 
+ bl[98] br[98] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_101 
+ bl[99] br[99] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_102 
+ bl[100] br[100] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_103 
+ bl[101] br[101] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_104 
+ bl[102] br[102] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_105 
+ bl[103] br[103] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_106 
+ bl[104] br[104] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_107 
+ bl[105] br[105] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_108 
+ bl[106] br[106] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_109 
+ bl[107] br[107] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_110 
+ bl[108] br[108] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_111 
+ bl[109] br[109] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_112 
+ bl[110] br[110] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_113 
+ bl[111] br[111] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_114 
+ bl[112] br[112] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_115 
+ bl[113] br[113] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_116 
+ bl[114] br[114] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_117 
+ bl[115] br[115] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_118 
+ bl[116] br[116] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_119 
+ bl[117] br[117] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_120 
+ bl[118] br[118] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_121 
+ bl[119] br[119] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_122 
+ bl[120] br[120] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_123 
+ bl[121] br[121] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_124 
+ bl[122] br[122] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_125 
+ bl[123] br[123] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_126 
+ bl[124] br[124] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_127 
+ bl[125] br[125] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_128 
+ bl[126] br[126] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_129 
+ bl[127] br[127] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_130 
+ vdd vdd vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_131 
+ vdd vdd vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_0 
+ vdd vdd vss vdd vpb vnb wl[4] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_6_1 
+ rbl rbr vss vdd vpb vnb wl[4] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_6_2 
+ bl[0] br[0] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_3 
+ bl[1] br[1] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_4 
+ bl[2] br[2] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_5 
+ bl[3] br[3] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_6 
+ bl[4] br[4] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_7 
+ bl[5] br[5] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_8 
+ bl[6] br[6] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_9 
+ bl[7] br[7] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_10 
+ bl[8] br[8] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_11 
+ bl[9] br[9] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_12 
+ bl[10] br[10] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_13 
+ bl[11] br[11] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_14 
+ bl[12] br[12] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_15 
+ bl[13] br[13] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_16 
+ bl[14] br[14] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_17 
+ bl[15] br[15] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_18 
+ bl[16] br[16] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_19 
+ bl[17] br[17] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_20 
+ bl[18] br[18] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_21 
+ bl[19] br[19] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_22 
+ bl[20] br[20] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_23 
+ bl[21] br[21] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_24 
+ bl[22] br[22] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_25 
+ bl[23] br[23] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_26 
+ bl[24] br[24] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_27 
+ bl[25] br[25] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_28 
+ bl[26] br[26] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_29 
+ bl[27] br[27] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_30 
+ bl[28] br[28] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_31 
+ bl[29] br[29] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_32 
+ bl[30] br[30] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_33 
+ bl[31] br[31] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_34 
+ bl[32] br[32] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_35 
+ bl[33] br[33] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_36 
+ bl[34] br[34] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_37 
+ bl[35] br[35] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_38 
+ bl[36] br[36] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_39 
+ bl[37] br[37] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_40 
+ bl[38] br[38] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_41 
+ bl[39] br[39] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_42 
+ bl[40] br[40] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_43 
+ bl[41] br[41] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_44 
+ bl[42] br[42] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_45 
+ bl[43] br[43] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_46 
+ bl[44] br[44] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_47 
+ bl[45] br[45] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_48 
+ bl[46] br[46] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_49 
+ bl[47] br[47] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_50 
+ bl[48] br[48] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_51 
+ bl[49] br[49] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_52 
+ bl[50] br[50] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_53 
+ bl[51] br[51] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_54 
+ bl[52] br[52] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_55 
+ bl[53] br[53] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_56 
+ bl[54] br[54] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_57 
+ bl[55] br[55] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_58 
+ bl[56] br[56] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_59 
+ bl[57] br[57] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_60 
+ bl[58] br[58] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_61 
+ bl[59] br[59] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_62 
+ bl[60] br[60] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_63 
+ bl[61] br[61] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_64 
+ bl[62] br[62] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_65 
+ bl[63] br[63] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_66 
+ bl[64] br[64] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_67 
+ bl[65] br[65] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_68 
+ bl[66] br[66] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_69 
+ bl[67] br[67] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_70 
+ bl[68] br[68] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_71 
+ bl[69] br[69] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_72 
+ bl[70] br[70] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_73 
+ bl[71] br[71] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_74 
+ bl[72] br[72] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_75 
+ bl[73] br[73] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_76 
+ bl[74] br[74] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_77 
+ bl[75] br[75] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_78 
+ bl[76] br[76] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_79 
+ bl[77] br[77] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_80 
+ bl[78] br[78] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_81 
+ bl[79] br[79] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_82 
+ bl[80] br[80] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_83 
+ bl[81] br[81] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_84 
+ bl[82] br[82] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_85 
+ bl[83] br[83] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_86 
+ bl[84] br[84] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_87 
+ bl[85] br[85] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_88 
+ bl[86] br[86] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_89 
+ bl[87] br[87] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_90 
+ bl[88] br[88] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_91 
+ bl[89] br[89] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_92 
+ bl[90] br[90] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_93 
+ bl[91] br[91] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_94 
+ bl[92] br[92] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_95 
+ bl[93] br[93] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_96 
+ bl[94] br[94] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_97 
+ bl[95] br[95] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_98 
+ bl[96] br[96] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_99 
+ bl[97] br[97] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_100 
+ bl[98] br[98] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_101 
+ bl[99] br[99] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_102 
+ bl[100] br[100] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_103 
+ bl[101] br[101] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_104 
+ bl[102] br[102] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_105 
+ bl[103] br[103] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_106 
+ bl[104] br[104] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_107 
+ bl[105] br[105] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_108 
+ bl[106] br[106] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_109 
+ bl[107] br[107] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_110 
+ bl[108] br[108] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_111 
+ bl[109] br[109] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_112 
+ bl[110] br[110] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_113 
+ bl[111] br[111] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_114 
+ bl[112] br[112] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_115 
+ bl[113] br[113] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_116 
+ bl[114] br[114] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_117 
+ bl[115] br[115] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_118 
+ bl[116] br[116] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_119 
+ bl[117] br[117] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_120 
+ bl[118] br[118] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_121 
+ bl[119] br[119] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_122 
+ bl[120] br[120] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_123 
+ bl[121] br[121] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_124 
+ bl[122] br[122] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_125 
+ bl[123] br[123] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_126 
+ bl[124] br[124] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_127 
+ bl[125] br[125] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_128 
+ bl[126] br[126] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_129 
+ bl[127] br[127] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_130 
+ vdd vdd vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_131 
+ vdd vdd vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_0 
+ vdd vdd vss vdd vpb vnb wl[5] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_7_1 
+ rbl rbr vss vdd vpb vnb wl[5] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_7_2 
+ bl[0] br[0] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_3 
+ bl[1] br[1] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_4 
+ bl[2] br[2] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_5 
+ bl[3] br[3] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_6 
+ bl[4] br[4] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_7 
+ bl[5] br[5] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_8 
+ bl[6] br[6] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_9 
+ bl[7] br[7] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_10 
+ bl[8] br[8] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_11 
+ bl[9] br[9] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_12 
+ bl[10] br[10] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_13 
+ bl[11] br[11] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_14 
+ bl[12] br[12] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_15 
+ bl[13] br[13] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_16 
+ bl[14] br[14] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_17 
+ bl[15] br[15] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_18 
+ bl[16] br[16] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_19 
+ bl[17] br[17] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_20 
+ bl[18] br[18] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_21 
+ bl[19] br[19] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_22 
+ bl[20] br[20] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_23 
+ bl[21] br[21] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_24 
+ bl[22] br[22] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_25 
+ bl[23] br[23] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_26 
+ bl[24] br[24] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_27 
+ bl[25] br[25] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_28 
+ bl[26] br[26] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_29 
+ bl[27] br[27] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_30 
+ bl[28] br[28] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_31 
+ bl[29] br[29] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_32 
+ bl[30] br[30] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_33 
+ bl[31] br[31] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_34 
+ bl[32] br[32] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_35 
+ bl[33] br[33] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_36 
+ bl[34] br[34] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_37 
+ bl[35] br[35] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_38 
+ bl[36] br[36] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_39 
+ bl[37] br[37] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_40 
+ bl[38] br[38] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_41 
+ bl[39] br[39] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_42 
+ bl[40] br[40] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_43 
+ bl[41] br[41] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_44 
+ bl[42] br[42] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_45 
+ bl[43] br[43] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_46 
+ bl[44] br[44] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_47 
+ bl[45] br[45] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_48 
+ bl[46] br[46] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_49 
+ bl[47] br[47] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_50 
+ bl[48] br[48] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_51 
+ bl[49] br[49] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_52 
+ bl[50] br[50] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_53 
+ bl[51] br[51] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_54 
+ bl[52] br[52] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_55 
+ bl[53] br[53] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_56 
+ bl[54] br[54] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_57 
+ bl[55] br[55] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_58 
+ bl[56] br[56] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_59 
+ bl[57] br[57] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_60 
+ bl[58] br[58] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_61 
+ bl[59] br[59] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_62 
+ bl[60] br[60] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_63 
+ bl[61] br[61] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_64 
+ bl[62] br[62] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_65 
+ bl[63] br[63] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_66 
+ bl[64] br[64] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_67 
+ bl[65] br[65] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_68 
+ bl[66] br[66] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_69 
+ bl[67] br[67] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_70 
+ bl[68] br[68] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_71 
+ bl[69] br[69] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_72 
+ bl[70] br[70] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_73 
+ bl[71] br[71] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_74 
+ bl[72] br[72] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_75 
+ bl[73] br[73] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_76 
+ bl[74] br[74] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_77 
+ bl[75] br[75] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_78 
+ bl[76] br[76] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_79 
+ bl[77] br[77] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_80 
+ bl[78] br[78] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_81 
+ bl[79] br[79] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_82 
+ bl[80] br[80] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_83 
+ bl[81] br[81] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_84 
+ bl[82] br[82] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_85 
+ bl[83] br[83] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_86 
+ bl[84] br[84] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_87 
+ bl[85] br[85] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_88 
+ bl[86] br[86] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_89 
+ bl[87] br[87] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_90 
+ bl[88] br[88] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_91 
+ bl[89] br[89] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_92 
+ bl[90] br[90] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_93 
+ bl[91] br[91] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_94 
+ bl[92] br[92] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_95 
+ bl[93] br[93] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_96 
+ bl[94] br[94] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_97 
+ bl[95] br[95] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_98 
+ bl[96] br[96] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_99 
+ bl[97] br[97] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_100 
+ bl[98] br[98] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_101 
+ bl[99] br[99] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_102 
+ bl[100] br[100] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_103 
+ bl[101] br[101] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_104 
+ bl[102] br[102] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_105 
+ bl[103] br[103] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_106 
+ bl[104] br[104] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_107 
+ bl[105] br[105] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_108 
+ bl[106] br[106] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_109 
+ bl[107] br[107] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_110 
+ bl[108] br[108] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_111 
+ bl[109] br[109] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_112 
+ bl[110] br[110] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_113 
+ bl[111] br[111] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_114 
+ bl[112] br[112] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_115 
+ bl[113] br[113] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_116 
+ bl[114] br[114] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_117 
+ bl[115] br[115] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_118 
+ bl[116] br[116] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_119 
+ bl[117] br[117] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_120 
+ bl[118] br[118] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_121 
+ bl[119] br[119] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_122 
+ bl[120] br[120] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_123 
+ bl[121] br[121] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_124 
+ bl[122] br[122] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_125 
+ bl[123] br[123] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_126 
+ bl[124] br[124] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_127 
+ bl[125] br[125] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_128 
+ bl[126] br[126] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_129 
+ bl[127] br[127] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_130 
+ vdd vdd vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_131 
+ vdd vdd vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_0 
+ vdd vdd vss vdd vpb vnb wl[6] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_8_1 
+ rbl rbr vss vdd vpb vnb wl[6] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_8_2 
+ bl[0] br[0] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_3 
+ bl[1] br[1] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_4 
+ bl[2] br[2] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_5 
+ bl[3] br[3] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_6 
+ bl[4] br[4] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_7 
+ bl[5] br[5] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_8 
+ bl[6] br[6] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_9 
+ bl[7] br[7] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_10 
+ bl[8] br[8] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_11 
+ bl[9] br[9] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_12 
+ bl[10] br[10] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_13 
+ bl[11] br[11] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_14 
+ bl[12] br[12] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_15 
+ bl[13] br[13] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_16 
+ bl[14] br[14] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_17 
+ bl[15] br[15] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_18 
+ bl[16] br[16] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_19 
+ bl[17] br[17] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_20 
+ bl[18] br[18] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_21 
+ bl[19] br[19] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_22 
+ bl[20] br[20] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_23 
+ bl[21] br[21] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_24 
+ bl[22] br[22] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_25 
+ bl[23] br[23] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_26 
+ bl[24] br[24] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_27 
+ bl[25] br[25] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_28 
+ bl[26] br[26] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_29 
+ bl[27] br[27] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_30 
+ bl[28] br[28] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_31 
+ bl[29] br[29] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_32 
+ bl[30] br[30] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_33 
+ bl[31] br[31] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_34 
+ bl[32] br[32] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_35 
+ bl[33] br[33] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_36 
+ bl[34] br[34] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_37 
+ bl[35] br[35] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_38 
+ bl[36] br[36] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_39 
+ bl[37] br[37] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_40 
+ bl[38] br[38] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_41 
+ bl[39] br[39] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_42 
+ bl[40] br[40] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_43 
+ bl[41] br[41] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_44 
+ bl[42] br[42] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_45 
+ bl[43] br[43] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_46 
+ bl[44] br[44] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_47 
+ bl[45] br[45] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_48 
+ bl[46] br[46] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_49 
+ bl[47] br[47] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_50 
+ bl[48] br[48] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_51 
+ bl[49] br[49] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_52 
+ bl[50] br[50] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_53 
+ bl[51] br[51] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_54 
+ bl[52] br[52] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_55 
+ bl[53] br[53] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_56 
+ bl[54] br[54] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_57 
+ bl[55] br[55] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_58 
+ bl[56] br[56] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_59 
+ bl[57] br[57] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_60 
+ bl[58] br[58] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_61 
+ bl[59] br[59] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_62 
+ bl[60] br[60] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_63 
+ bl[61] br[61] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_64 
+ bl[62] br[62] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_65 
+ bl[63] br[63] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_66 
+ bl[64] br[64] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_67 
+ bl[65] br[65] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_68 
+ bl[66] br[66] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_69 
+ bl[67] br[67] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_70 
+ bl[68] br[68] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_71 
+ bl[69] br[69] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_72 
+ bl[70] br[70] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_73 
+ bl[71] br[71] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_74 
+ bl[72] br[72] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_75 
+ bl[73] br[73] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_76 
+ bl[74] br[74] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_77 
+ bl[75] br[75] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_78 
+ bl[76] br[76] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_79 
+ bl[77] br[77] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_80 
+ bl[78] br[78] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_81 
+ bl[79] br[79] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_82 
+ bl[80] br[80] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_83 
+ bl[81] br[81] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_84 
+ bl[82] br[82] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_85 
+ bl[83] br[83] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_86 
+ bl[84] br[84] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_87 
+ bl[85] br[85] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_88 
+ bl[86] br[86] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_89 
+ bl[87] br[87] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_90 
+ bl[88] br[88] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_91 
+ bl[89] br[89] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_92 
+ bl[90] br[90] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_93 
+ bl[91] br[91] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_94 
+ bl[92] br[92] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_95 
+ bl[93] br[93] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_96 
+ bl[94] br[94] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_97 
+ bl[95] br[95] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_98 
+ bl[96] br[96] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_99 
+ bl[97] br[97] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_100 
+ bl[98] br[98] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_101 
+ bl[99] br[99] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_102 
+ bl[100] br[100] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_103 
+ bl[101] br[101] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_104 
+ bl[102] br[102] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_105 
+ bl[103] br[103] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_106 
+ bl[104] br[104] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_107 
+ bl[105] br[105] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_108 
+ bl[106] br[106] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_109 
+ bl[107] br[107] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_110 
+ bl[108] br[108] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_111 
+ bl[109] br[109] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_112 
+ bl[110] br[110] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_113 
+ bl[111] br[111] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_114 
+ bl[112] br[112] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_115 
+ bl[113] br[113] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_116 
+ bl[114] br[114] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_117 
+ bl[115] br[115] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_118 
+ bl[116] br[116] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_119 
+ bl[117] br[117] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_120 
+ bl[118] br[118] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_121 
+ bl[119] br[119] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_122 
+ bl[120] br[120] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_123 
+ bl[121] br[121] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_124 
+ bl[122] br[122] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_125 
+ bl[123] br[123] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_126 
+ bl[124] br[124] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_127 
+ bl[125] br[125] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_128 
+ bl[126] br[126] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_129 
+ bl[127] br[127] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_130 
+ vdd vdd vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_131 
+ vdd vdd vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_0 
+ vdd vdd vss vdd vpb vnb wl[7] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_9_1 
+ rbl rbr vss vdd vpb vnb wl[7] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_9_2 
+ bl[0] br[0] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_3 
+ bl[1] br[1] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_4 
+ bl[2] br[2] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_5 
+ bl[3] br[3] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_6 
+ bl[4] br[4] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_7 
+ bl[5] br[5] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_8 
+ bl[6] br[6] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_9 
+ bl[7] br[7] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_10 
+ bl[8] br[8] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_11 
+ bl[9] br[9] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_12 
+ bl[10] br[10] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_13 
+ bl[11] br[11] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_14 
+ bl[12] br[12] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_15 
+ bl[13] br[13] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_16 
+ bl[14] br[14] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_17 
+ bl[15] br[15] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_18 
+ bl[16] br[16] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_19 
+ bl[17] br[17] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_20 
+ bl[18] br[18] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_21 
+ bl[19] br[19] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_22 
+ bl[20] br[20] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_23 
+ bl[21] br[21] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_24 
+ bl[22] br[22] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_25 
+ bl[23] br[23] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_26 
+ bl[24] br[24] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_27 
+ bl[25] br[25] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_28 
+ bl[26] br[26] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_29 
+ bl[27] br[27] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_30 
+ bl[28] br[28] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_31 
+ bl[29] br[29] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_32 
+ bl[30] br[30] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_33 
+ bl[31] br[31] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_34 
+ bl[32] br[32] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_35 
+ bl[33] br[33] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_36 
+ bl[34] br[34] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_37 
+ bl[35] br[35] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_38 
+ bl[36] br[36] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_39 
+ bl[37] br[37] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_40 
+ bl[38] br[38] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_41 
+ bl[39] br[39] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_42 
+ bl[40] br[40] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_43 
+ bl[41] br[41] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_44 
+ bl[42] br[42] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_45 
+ bl[43] br[43] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_46 
+ bl[44] br[44] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_47 
+ bl[45] br[45] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_48 
+ bl[46] br[46] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_49 
+ bl[47] br[47] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_50 
+ bl[48] br[48] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_51 
+ bl[49] br[49] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_52 
+ bl[50] br[50] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_53 
+ bl[51] br[51] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_54 
+ bl[52] br[52] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_55 
+ bl[53] br[53] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_56 
+ bl[54] br[54] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_57 
+ bl[55] br[55] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_58 
+ bl[56] br[56] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_59 
+ bl[57] br[57] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_60 
+ bl[58] br[58] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_61 
+ bl[59] br[59] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_62 
+ bl[60] br[60] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_63 
+ bl[61] br[61] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_64 
+ bl[62] br[62] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_65 
+ bl[63] br[63] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_66 
+ bl[64] br[64] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_67 
+ bl[65] br[65] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_68 
+ bl[66] br[66] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_69 
+ bl[67] br[67] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_70 
+ bl[68] br[68] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_71 
+ bl[69] br[69] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_72 
+ bl[70] br[70] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_73 
+ bl[71] br[71] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_74 
+ bl[72] br[72] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_75 
+ bl[73] br[73] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_76 
+ bl[74] br[74] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_77 
+ bl[75] br[75] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_78 
+ bl[76] br[76] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_79 
+ bl[77] br[77] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_80 
+ bl[78] br[78] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_81 
+ bl[79] br[79] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_82 
+ bl[80] br[80] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_83 
+ bl[81] br[81] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_84 
+ bl[82] br[82] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_85 
+ bl[83] br[83] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_86 
+ bl[84] br[84] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_87 
+ bl[85] br[85] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_88 
+ bl[86] br[86] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_89 
+ bl[87] br[87] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_90 
+ bl[88] br[88] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_91 
+ bl[89] br[89] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_92 
+ bl[90] br[90] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_93 
+ bl[91] br[91] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_94 
+ bl[92] br[92] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_95 
+ bl[93] br[93] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_96 
+ bl[94] br[94] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_97 
+ bl[95] br[95] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_98 
+ bl[96] br[96] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_99 
+ bl[97] br[97] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_100 
+ bl[98] br[98] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_101 
+ bl[99] br[99] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_102 
+ bl[100] br[100] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_103 
+ bl[101] br[101] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_104 
+ bl[102] br[102] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_105 
+ bl[103] br[103] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_106 
+ bl[104] br[104] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_107 
+ bl[105] br[105] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_108 
+ bl[106] br[106] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_109 
+ bl[107] br[107] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_110 
+ bl[108] br[108] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_111 
+ bl[109] br[109] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_112 
+ bl[110] br[110] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_113 
+ bl[111] br[111] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_114 
+ bl[112] br[112] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_115 
+ bl[113] br[113] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_116 
+ bl[114] br[114] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_117 
+ bl[115] br[115] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_118 
+ bl[116] br[116] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_119 
+ bl[117] br[117] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_120 
+ bl[118] br[118] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_121 
+ bl[119] br[119] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_122 
+ bl[120] br[120] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_123 
+ bl[121] br[121] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_124 
+ bl[122] br[122] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_125 
+ bl[123] br[123] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_126 
+ bl[124] br[124] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_127 
+ bl[125] br[125] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_128 
+ bl[126] br[126] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_129 
+ bl[127] br[127] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_130 
+ vdd vdd vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_131 
+ vdd vdd vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_0 
+ vdd vdd vss vdd vpb vnb wl[8] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_10_1 
+ rbl rbr vss vdd vpb vnb wl[8] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_10_2 
+ bl[0] br[0] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_3 
+ bl[1] br[1] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_4 
+ bl[2] br[2] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_5 
+ bl[3] br[3] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_6 
+ bl[4] br[4] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_7 
+ bl[5] br[5] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_8 
+ bl[6] br[6] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_9 
+ bl[7] br[7] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_10 
+ bl[8] br[8] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_11 
+ bl[9] br[9] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_12 
+ bl[10] br[10] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_13 
+ bl[11] br[11] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_14 
+ bl[12] br[12] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_15 
+ bl[13] br[13] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_16 
+ bl[14] br[14] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_17 
+ bl[15] br[15] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_18 
+ bl[16] br[16] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_19 
+ bl[17] br[17] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_20 
+ bl[18] br[18] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_21 
+ bl[19] br[19] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_22 
+ bl[20] br[20] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_23 
+ bl[21] br[21] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_24 
+ bl[22] br[22] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_25 
+ bl[23] br[23] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_26 
+ bl[24] br[24] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_27 
+ bl[25] br[25] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_28 
+ bl[26] br[26] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_29 
+ bl[27] br[27] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_30 
+ bl[28] br[28] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_31 
+ bl[29] br[29] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_32 
+ bl[30] br[30] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_33 
+ bl[31] br[31] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_34 
+ bl[32] br[32] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_35 
+ bl[33] br[33] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_36 
+ bl[34] br[34] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_37 
+ bl[35] br[35] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_38 
+ bl[36] br[36] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_39 
+ bl[37] br[37] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_40 
+ bl[38] br[38] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_41 
+ bl[39] br[39] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_42 
+ bl[40] br[40] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_43 
+ bl[41] br[41] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_44 
+ bl[42] br[42] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_45 
+ bl[43] br[43] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_46 
+ bl[44] br[44] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_47 
+ bl[45] br[45] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_48 
+ bl[46] br[46] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_49 
+ bl[47] br[47] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_50 
+ bl[48] br[48] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_51 
+ bl[49] br[49] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_52 
+ bl[50] br[50] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_53 
+ bl[51] br[51] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_54 
+ bl[52] br[52] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_55 
+ bl[53] br[53] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_56 
+ bl[54] br[54] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_57 
+ bl[55] br[55] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_58 
+ bl[56] br[56] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_59 
+ bl[57] br[57] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_60 
+ bl[58] br[58] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_61 
+ bl[59] br[59] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_62 
+ bl[60] br[60] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_63 
+ bl[61] br[61] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_64 
+ bl[62] br[62] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_65 
+ bl[63] br[63] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_66 
+ bl[64] br[64] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_67 
+ bl[65] br[65] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_68 
+ bl[66] br[66] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_69 
+ bl[67] br[67] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_70 
+ bl[68] br[68] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_71 
+ bl[69] br[69] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_72 
+ bl[70] br[70] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_73 
+ bl[71] br[71] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_74 
+ bl[72] br[72] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_75 
+ bl[73] br[73] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_76 
+ bl[74] br[74] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_77 
+ bl[75] br[75] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_78 
+ bl[76] br[76] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_79 
+ bl[77] br[77] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_80 
+ bl[78] br[78] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_81 
+ bl[79] br[79] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_82 
+ bl[80] br[80] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_83 
+ bl[81] br[81] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_84 
+ bl[82] br[82] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_85 
+ bl[83] br[83] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_86 
+ bl[84] br[84] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_87 
+ bl[85] br[85] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_88 
+ bl[86] br[86] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_89 
+ bl[87] br[87] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_90 
+ bl[88] br[88] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_91 
+ bl[89] br[89] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_92 
+ bl[90] br[90] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_93 
+ bl[91] br[91] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_94 
+ bl[92] br[92] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_95 
+ bl[93] br[93] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_96 
+ bl[94] br[94] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_97 
+ bl[95] br[95] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_98 
+ bl[96] br[96] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_99 
+ bl[97] br[97] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_100 
+ bl[98] br[98] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_101 
+ bl[99] br[99] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_102 
+ bl[100] br[100] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_103 
+ bl[101] br[101] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_104 
+ bl[102] br[102] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_105 
+ bl[103] br[103] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_106 
+ bl[104] br[104] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_107 
+ bl[105] br[105] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_108 
+ bl[106] br[106] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_109 
+ bl[107] br[107] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_110 
+ bl[108] br[108] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_111 
+ bl[109] br[109] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_112 
+ bl[110] br[110] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_113 
+ bl[111] br[111] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_114 
+ bl[112] br[112] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_115 
+ bl[113] br[113] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_116 
+ bl[114] br[114] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_117 
+ bl[115] br[115] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_118 
+ bl[116] br[116] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_119 
+ bl[117] br[117] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_120 
+ bl[118] br[118] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_121 
+ bl[119] br[119] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_122 
+ bl[120] br[120] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_123 
+ bl[121] br[121] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_124 
+ bl[122] br[122] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_125 
+ bl[123] br[123] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_126 
+ bl[124] br[124] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_127 
+ bl[125] br[125] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_128 
+ bl[126] br[126] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_129 
+ bl[127] br[127] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_130 
+ vdd vdd vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_131 
+ vdd vdd vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_0 
+ vdd vdd vss vdd vpb vnb wl[9] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_11_1 
+ rbl rbr vss vdd vpb vnb wl[9] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_11_2 
+ bl[0] br[0] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_3 
+ bl[1] br[1] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_4 
+ bl[2] br[2] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_5 
+ bl[3] br[3] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_6 
+ bl[4] br[4] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_7 
+ bl[5] br[5] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_8 
+ bl[6] br[6] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_9 
+ bl[7] br[7] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_10 
+ bl[8] br[8] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_11 
+ bl[9] br[9] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_12 
+ bl[10] br[10] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_13 
+ bl[11] br[11] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_14 
+ bl[12] br[12] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_15 
+ bl[13] br[13] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_16 
+ bl[14] br[14] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_17 
+ bl[15] br[15] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_18 
+ bl[16] br[16] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_19 
+ bl[17] br[17] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_20 
+ bl[18] br[18] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_21 
+ bl[19] br[19] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_22 
+ bl[20] br[20] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_23 
+ bl[21] br[21] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_24 
+ bl[22] br[22] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_25 
+ bl[23] br[23] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_26 
+ bl[24] br[24] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_27 
+ bl[25] br[25] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_28 
+ bl[26] br[26] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_29 
+ bl[27] br[27] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_30 
+ bl[28] br[28] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_31 
+ bl[29] br[29] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_32 
+ bl[30] br[30] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_33 
+ bl[31] br[31] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_34 
+ bl[32] br[32] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_35 
+ bl[33] br[33] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_36 
+ bl[34] br[34] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_37 
+ bl[35] br[35] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_38 
+ bl[36] br[36] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_39 
+ bl[37] br[37] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_40 
+ bl[38] br[38] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_41 
+ bl[39] br[39] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_42 
+ bl[40] br[40] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_43 
+ bl[41] br[41] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_44 
+ bl[42] br[42] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_45 
+ bl[43] br[43] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_46 
+ bl[44] br[44] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_47 
+ bl[45] br[45] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_48 
+ bl[46] br[46] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_49 
+ bl[47] br[47] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_50 
+ bl[48] br[48] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_51 
+ bl[49] br[49] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_52 
+ bl[50] br[50] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_53 
+ bl[51] br[51] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_54 
+ bl[52] br[52] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_55 
+ bl[53] br[53] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_56 
+ bl[54] br[54] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_57 
+ bl[55] br[55] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_58 
+ bl[56] br[56] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_59 
+ bl[57] br[57] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_60 
+ bl[58] br[58] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_61 
+ bl[59] br[59] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_62 
+ bl[60] br[60] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_63 
+ bl[61] br[61] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_64 
+ bl[62] br[62] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_65 
+ bl[63] br[63] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_66 
+ bl[64] br[64] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_67 
+ bl[65] br[65] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_68 
+ bl[66] br[66] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_69 
+ bl[67] br[67] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_70 
+ bl[68] br[68] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_71 
+ bl[69] br[69] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_72 
+ bl[70] br[70] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_73 
+ bl[71] br[71] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_74 
+ bl[72] br[72] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_75 
+ bl[73] br[73] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_76 
+ bl[74] br[74] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_77 
+ bl[75] br[75] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_78 
+ bl[76] br[76] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_79 
+ bl[77] br[77] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_80 
+ bl[78] br[78] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_81 
+ bl[79] br[79] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_82 
+ bl[80] br[80] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_83 
+ bl[81] br[81] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_84 
+ bl[82] br[82] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_85 
+ bl[83] br[83] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_86 
+ bl[84] br[84] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_87 
+ bl[85] br[85] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_88 
+ bl[86] br[86] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_89 
+ bl[87] br[87] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_90 
+ bl[88] br[88] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_91 
+ bl[89] br[89] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_92 
+ bl[90] br[90] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_93 
+ bl[91] br[91] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_94 
+ bl[92] br[92] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_95 
+ bl[93] br[93] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_96 
+ bl[94] br[94] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_97 
+ bl[95] br[95] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_98 
+ bl[96] br[96] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_99 
+ bl[97] br[97] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_100 
+ bl[98] br[98] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_101 
+ bl[99] br[99] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_102 
+ bl[100] br[100] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_103 
+ bl[101] br[101] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_104 
+ bl[102] br[102] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_105 
+ bl[103] br[103] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_106 
+ bl[104] br[104] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_107 
+ bl[105] br[105] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_108 
+ bl[106] br[106] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_109 
+ bl[107] br[107] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_110 
+ bl[108] br[108] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_111 
+ bl[109] br[109] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_112 
+ bl[110] br[110] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_113 
+ bl[111] br[111] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_114 
+ bl[112] br[112] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_115 
+ bl[113] br[113] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_116 
+ bl[114] br[114] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_117 
+ bl[115] br[115] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_118 
+ bl[116] br[116] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_119 
+ bl[117] br[117] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_120 
+ bl[118] br[118] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_121 
+ bl[119] br[119] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_122 
+ bl[120] br[120] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_123 
+ bl[121] br[121] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_124 
+ bl[122] br[122] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_125 
+ bl[123] br[123] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_126 
+ bl[124] br[124] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_127 
+ bl[125] br[125] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_128 
+ bl[126] br[126] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_129 
+ bl[127] br[127] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_130 
+ vdd vdd vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_131 
+ vdd vdd vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_0 
+ vdd vdd vss vdd vpb vnb wl[10] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_12_1 
+ rbl rbr vss vdd vpb vnb wl[10] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_12_2 
+ bl[0] br[0] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_3 
+ bl[1] br[1] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_4 
+ bl[2] br[2] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_5 
+ bl[3] br[3] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_6 
+ bl[4] br[4] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_7 
+ bl[5] br[5] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_8 
+ bl[6] br[6] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_9 
+ bl[7] br[7] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_10 
+ bl[8] br[8] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_11 
+ bl[9] br[9] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_12 
+ bl[10] br[10] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_13 
+ bl[11] br[11] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_14 
+ bl[12] br[12] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_15 
+ bl[13] br[13] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_16 
+ bl[14] br[14] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_17 
+ bl[15] br[15] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_18 
+ bl[16] br[16] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_19 
+ bl[17] br[17] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_20 
+ bl[18] br[18] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_21 
+ bl[19] br[19] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_22 
+ bl[20] br[20] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_23 
+ bl[21] br[21] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_24 
+ bl[22] br[22] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_25 
+ bl[23] br[23] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_26 
+ bl[24] br[24] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_27 
+ bl[25] br[25] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_28 
+ bl[26] br[26] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_29 
+ bl[27] br[27] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_30 
+ bl[28] br[28] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_31 
+ bl[29] br[29] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_32 
+ bl[30] br[30] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_33 
+ bl[31] br[31] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_34 
+ bl[32] br[32] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_35 
+ bl[33] br[33] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_36 
+ bl[34] br[34] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_37 
+ bl[35] br[35] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_38 
+ bl[36] br[36] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_39 
+ bl[37] br[37] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_40 
+ bl[38] br[38] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_41 
+ bl[39] br[39] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_42 
+ bl[40] br[40] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_43 
+ bl[41] br[41] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_44 
+ bl[42] br[42] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_45 
+ bl[43] br[43] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_46 
+ bl[44] br[44] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_47 
+ bl[45] br[45] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_48 
+ bl[46] br[46] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_49 
+ bl[47] br[47] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_50 
+ bl[48] br[48] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_51 
+ bl[49] br[49] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_52 
+ bl[50] br[50] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_53 
+ bl[51] br[51] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_54 
+ bl[52] br[52] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_55 
+ bl[53] br[53] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_56 
+ bl[54] br[54] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_57 
+ bl[55] br[55] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_58 
+ bl[56] br[56] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_59 
+ bl[57] br[57] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_60 
+ bl[58] br[58] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_61 
+ bl[59] br[59] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_62 
+ bl[60] br[60] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_63 
+ bl[61] br[61] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_64 
+ bl[62] br[62] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_65 
+ bl[63] br[63] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_66 
+ bl[64] br[64] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_67 
+ bl[65] br[65] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_68 
+ bl[66] br[66] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_69 
+ bl[67] br[67] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_70 
+ bl[68] br[68] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_71 
+ bl[69] br[69] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_72 
+ bl[70] br[70] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_73 
+ bl[71] br[71] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_74 
+ bl[72] br[72] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_75 
+ bl[73] br[73] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_76 
+ bl[74] br[74] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_77 
+ bl[75] br[75] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_78 
+ bl[76] br[76] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_79 
+ bl[77] br[77] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_80 
+ bl[78] br[78] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_81 
+ bl[79] br[79] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_82 
+ bl[80] br[80] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_83 
+ bl[81] br[81] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_84 
+ bl[82] br[82] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_85 
+ bl[83] br[83] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_86 
+ bl[84] br[84] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_87 
+ bl[85] br[85] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_88 
+ bl[86] br[86] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_89 
+ bl[87] br[87] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_90 
+ bl[88] br[88] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_91 
+ bl[89] br[89] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_92 
+ bl[90] br[90] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_93 
+ bl[91] br[91] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_94 
+ bl[92] br[92] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_95 
+ bl[93] br[93] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_96 
+ bl[94] br[94] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_97 
+ bl[95] br[95] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_98 
+ bl[96] br[96] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_99 
+ bl[97] br[97] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_100 
+ bl[98] br[98] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_101 
+ bl[99] br[99] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_102 
+ bl[100] br[100] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_103 
+ bl[101] br[101] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_104 
+ bl[102] br[102] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_105 
+ bl[103] br[103] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_106 
+ bl[104] br[104] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_107 
+ bl[105] br[105] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_108 
+ bl[106] br[106] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_109 
+ bl[107] br[107] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_110 
+ bl[108] br[108] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_111 
+ bl[109] br[109] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_112 
+ bl[110] br[110] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_113 
+ bl[111] br[111] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_114 
+ bl[112] br[112] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_115 
+ bl[113] br[113] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_116 
+ bl[114] br[114] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_117 
+ bl[115] br[115] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_118 
+ bl[116] br[116] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_119 
+ bl[117] br[117] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_120 
+ bl[118] br[118] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_121 
+ bl[119] br[119] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_122 
+ bl[120] br[120] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_123 
+ bl[121] br[121] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_124 
+ bl[122] br[122] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_125 
+ bl[123] br[123] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_126 
+ bl[124] br[124] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_127 
+ bl[125] br[125] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_128 
+ bl[126] br[126] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_129 
+ bl[127] br[127] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_130 
+ vdd vdd vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_131 
+ vdd vdd vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_0 
+ vdd vdd vss vdd vpb vnb wl[11] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_13_1 
+ rbl rbr vss vdd vpb vnb wl[11] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_13_2 
+ bl[0] br[0] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_3 
+ bl[1] br[1] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_4 
+ bl[2] br[2] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_5 
+ bl[3] br[3] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_6 
+ bl[4] br[4] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_7 
+ bl[5] br[5] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_8 
+ bl[6] br[6] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_9 
+ bl[7] br[7] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_10 
+ bl[8] br[8] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_11 
+ bl[9] br[9] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_12 
+ bl[10] br[10] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_13 
+ bl[11] br[11] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_14 
+ bl[12] br[12] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_15 
+ bl[13] br[13] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_16 
+ bl[14] br[14] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_17 
+ bl[15] br[15] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_18 
+ bl[16] br[16] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_19 
+ bl[17] br[17] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_20 
+ bl[18] br[18] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_21 
+ bl[19] br[19] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_22 
+ bl[20] br[20] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_23 
+ bl[21] br[21] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_24 
+ bl[22] br[22] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_25 
+ bl[23] br[23] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_26 
+ bl[24] br[24] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_27 
+ bl[25] br[25] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_28 
+ bl[26] br[26] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_29 
+ bl[27] br[27] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_30 
+ bl[28] br[28] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_31 
+ bl[29] br[29] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_32 
+ bl[30] br[30] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_33 
+ bl[31] br[31] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_34 
+ bl[32] br[32] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_35 
+ bl[33] br[33] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_36 
+ bl[34] br[34] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_37 
+ bl[35] br[35] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_38 
+ bl[36] br[36] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_39 
+ bl[37] br[37] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_40 
+ bl[38] br[38] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_41 
+ bl[39] br[39] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_42 
+ bl[40] br[40] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_43 
+ bl[41] br[41] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_44 
+ bl[42] br[42] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_45 
+ bl[43] br[43] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_46 
+ bl[44] br[44] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_47 
+ bl[45] br[45] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_48 
+ bl[46] br[46] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_49 
+ bl[47] br[47] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_50 
+ bl[48] br[48] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_51 
+ bl[49] br[49] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_52 
+ bl[50] br[50] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_53 
+ bl[51] br[51] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_54 
+ bl[52] br[52] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_55 
+ bl[53] br[53] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_56 
+ bl[54] br[54] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_57 
+ bl[55] br[55] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_58 
+ bl[56] br[56] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_59 
+ bl[57] br[57] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_60 
+ bl[58] br[58] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_61 
+ bl[59] br[59] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_62 
+ bl[60] br[60] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_63 
+ bl[61] br[61] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_64 
+ bl[62] br[62] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_65 
+ bl[63] br[63] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_66 
+ bl[64] br[64] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_67 
+ bl[65] br[65] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_68 
+ bl[66] br[66] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_69 
+ bl[67] br[67] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_70 
+ bl[68] br[68] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_71 
+ bl[69] br[69] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_72 
+ bl[70] br[70] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_73 
+ bl[71] br[71] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_74 
+ bl[72] br[72] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_75 
+ bl[73] br[73] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_76 
+ bl[74] br[74] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_77 
+ bl[75] br[75] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_78 
+ bl[76] br[76] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_79 
+ bl[77] br[77] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_80 
+ bl[78] br[78] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_81 
+ bl[79] br[79] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_82 
+ bl[80] br[80] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_83 
+ bl[81] br[81] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_84 
+ bl[82] br[82] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_85 
+ bl[83] br[83] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_86 
+ bl[84] br[84] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_87 
+ bl[85] br[85] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_88 
+ bl[86] br[86] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_89 
+ bl[87] br[87] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_90 
+ bl[88] br[88] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_91 
+ bl[89] br[89] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_92 
+ bl[90] br[90] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_93 
+ bl[91] br[91] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_94 
+ bl[92] br[92] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_95 
+ bl[93] br[93] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_96 
+ bl[94] br[94] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_97 
+ bl[95] br[95] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_98 
+ bl[96] br[96] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_99 
+ bl[97] br[97] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_100 
+ bl[98] br[98] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_101 
+ bl[99] br[99] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_102 
+ bl[100] br[100] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_103 
+ bl[101] br[101] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_104 
+ bl[102] br[102] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_105 
+ bl[103] br[103] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_106 
+ bl[104] br[104] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_107 
+ bl[105] br[105] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_108 
+ bl[106] br[106] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_109 
+ bl[107] br[107] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_110 
+ bl[108] br[108] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_111 
+ bl[109] br[109] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_112 
+ bl[110] br[110] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_113 
+ bl[111] br[111] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_114 
+ bl[112] br[112] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_115 
+ bl[113] br[113] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_116 
+ bl[114] br[114] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_117 
+ bl[115] br[115] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_118 
+ bl[116] br[116] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_119 
+ bl[117] br[117] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_120 
+ bl[118] br[118] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_121 
+ bl[119] br[119] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_122 
+ bl[120] br[120] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_123 
+ bl[121] br[121] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_124 
+ bl[122] br[122] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_125 
+ bl[123] br[123] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_126 
+ bl[124] br[124] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_127 
+ bl[125] br[125] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_128 
+ bl[126] br[126] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_129 
+ bl[127] br[127] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_130 
+ vdd vdd vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_131 
+ vdd vdd vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_0 
+ vdd vdd vss vdd vpb vnb wl[12] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_14_1 
+ rbl rbr vss vdd vpb vnb wl[12] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_14_2 
+ bl[0] br[0] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_3 
+ bl[1] br[1] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_4 
+ bl[2] br[2] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_5 
+ bl[3] br[3] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_6 
+ bl[4] br[4] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_7 
+ bl[5] br[5] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_8 
+ bl[6] br[6] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_9 
+ bl[7] br[7] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_10 
+ bl[8] br[8] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_11 
+ bl[9] br[9] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_12 
+ bl[10] br[10] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_13 
+ bl[11] br[11] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_14 
+ bl[12] br[12] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_15 
+ bl[13] br[13] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_16 
+ bl[14] br[14] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_17 
+ bl[15] br[15] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_18 
+ bl[16] br[16] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_19 
+ bl[17] br[17] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_20 
+ bl[18] br[18] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_21 
+ bl[19] br[19] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_22 
+ bl[20] br[20] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_23 
+ bl[21] br[21] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_24 
+ bl[22] br[22] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_25 
+ bl[23] br[23] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_26 
+ bl[24] br[24] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_27 
+ bl[25] br[25] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_28 
+ bl[26] br[26] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_29 
+ bl[27] br[27] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_30 
+ bl[28] br[28] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_31 
+ bl[29] br[29] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_32 
+ bl[30] br[30] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_33 
+ bl[31] br[31] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_34 
+ bl[32] br[32] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_35 
+ bl[33] br[33] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_36 
+ bl[34] br[34] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_37 
+ bl[35] br[35] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_38 
+ bl[36] br[36] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_39 
+ bl[37] br[37] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_40 
+ bl[38] br[38] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_41 
+ bl[39] br[39] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_42 
+ bl[40] br[40] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_43 
+ bl[41] br[41] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_44 
+ bl[42] br[42] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_45 
+ bl[43] br[43] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_46 
+ bl[44] br[44] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_47 
+ bl[45] br[45] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_48 
+ bl[46] br[46] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_49 
+ bl[47] br[47] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_50 
+ bl[48] br[48] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_51 
+ bl[49] br[49] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_52 
+ bl[50] br[50] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_53 
+ bl[51] br[51] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_54 
+ bl[52] br[52] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_55 
+ bl[53] br[53] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_56 
+ bl[54] br[54] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_57 
+ bl[55] br[55] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_58 
+ bl[56] br[56] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_59 
+ bl[57] br[57] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_60 
+ bl[58] br[58] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_61 
+ bl[59] br[59] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_62 
+ bl[60] br[60] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_63 
+ bl[61] br[61] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_64 
+ bl[62] br[62] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_65 
+ bl[63] br[63] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_66 
+ bl[64] br[64] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_67 
+ bl[65] br[65] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_68 
+ bl[66] br[66] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_69 
+ bl[67] br[67] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_70 
+ bl[68] br[68] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_71 
+ bl[69] br[69] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_72 
+ bl[70] br[70] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_73 
+ bl[71] br[71] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_74 
+ bl[72] br[72] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_75 
+ bl[73] br[73] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_76 
+ bl[74] br[74] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_77 
+ bl[75] br[75] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_78 
+ bl[76] br[76] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_79 
+ bl[77] br[77] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_80 
+ bl[78] br[78] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_81 
+ bl[79] br[79] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_82 
+ bl[80] br[80] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_83 
+ bl[81] br[81] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_84 
+ bl[82] br[82] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_85 
+ bl[83] br[83] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_86 
+ bl[84] br[84] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_87 
+ bl[85] br[85] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_88 
+ bl[86] br[86] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_89 
+ bl[87] br[87] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_90 
+ bl[88] br[88] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_91 
+ bl[89] br[89] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_92 
+ bl[90] br[90] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_93 
+ bl[91] br[91] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_94 
+ bl[92] br[92] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_95 
+ bl[93] br[93] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_96 
+ bl[94] br[94] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_97 
+ bl[95] br[95] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_98 
+ bl[96] br[96] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_99 
+ bl[97] br[97] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_100 
+ bl[98] br[98] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_101 
+ bl[99] br[99] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_102 
+ bl[100] br[100] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_103 
+ bl[101] br[101] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_104 
+ bl[102] br[102] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_105 
+ bl[103] br[103] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_106 
+ bl[104] br[104] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_107 
+ bl[105] br[105] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_108 
+ bl[106] br[106] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_109 
+ bl[107] br[107] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_110 
+ bl[108] br[108] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_111 
+ bl[109] br[109] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_112 
+ bl[110] br[110] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_113 
+ bl[111] br[111] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_114 
+ bl[112] br[112] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_115 
+ bl[113] br[113] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_116 
+ bl[114] br[114] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_117 
+ bl[115] br[115] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_118 
+ bl[116] br[116] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_119 
+ bl[117] br[117] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_120 
+ bl[118] br[118] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_121 
+ bl[119] br[119] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_122 
+ bl[120] br[120] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_123 
+ bl[121] br[121] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_124 
+ bl[122] br[122] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_125 
+ bl[123] br[123] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_126 
+ bl[124] br[124] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_127 
+ bl[125] br[125] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_128 
+ bl[126] br[126] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_129 
+ bl[127] br[127] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_130 
+ vdd vdd vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_131 
+ vdd vdd vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_0 
+ vdd vdd vss vdd vpb vnb wl[13] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_15_1 
+ rbl rbr vss vdd vpb vnb wl[13] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_15_2 
+ bl[0] br[0] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_3 
+ bl[1] br[1] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_4 
+ bl[2] br[2] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_5 
+ bl[3] br[3] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_6 
+ bl[4] br[4] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_7 
+ bl[5] br[5] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_8 
+ bl[6] br[6] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_9 
+ bl[7] br[7] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_10 
+ bl[8] br[8] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_11 
+ bl[9] br[9] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_12 
+ bl[10] br[10] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_13 
+ bl[11] br[11] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_14 
+ bl[12] br[12] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_15 
+ bl[13] br[13] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_16 
+ bl[14] br[14] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_17 
+ bl[15] br[15] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_18 
+ bl[16] br[16] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_19 
+ bl[17] br[17] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_20 
+ bl[18] br[18] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_21 
+ bl[19] br[19] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_22 
+ bl[20] br[20] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_23 
+ bl[21] br[21] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_24 
+ bl[22] br[22] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_25 
+ bl[23] br[23] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_26 
+ bl[24] br[24] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_27 
+ bl[25] br[25] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_28 
+ bl[26] br[26] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_29 
+ bl[27] br[27] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_30 
+ bl[28] br[28] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_31 
+ bl[29] br[29] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_32 
+ bl[30] br[30] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_33 
+ bl[31] br[31] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_34 
+ bl[32] br[32] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_35 
+ bl[33] br[33] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_36 
+ bl[34] br[34] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_37 
+ bl[35] br[35] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_38 
+ bl[36] br[36] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_39 
+ bl[37] br[37] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_40 
+ bl[38] br[38] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_41 
+ bl[39] br[39] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_42 
+ bl[40] br[40] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_43 
+ bl[41] br[41] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_44 
+ bl[42] br[42] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_45 
+ bl[43] br[43] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_46 
+ bl[44] br[44] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_47 
+ bl[45] br[45] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_48 
+ bl[46] br[46] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_49 
+ bl[47] br[47] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_50 
+ bl[48] br[48] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_51 
+ bl[49] br[49] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_52 
+ bl[50] br[50] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_53 
+ bl[51] br[51] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_54 
+ bl[52] br[52] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_55 
+ bl[53] br[53] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_56 
+ bl[54] br[54] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_57 
+ bl[55] br[55] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_58 
+ bl[56] br[56] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_59 
+ bl[57] br[57] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_60 
+ bl[58] br[58] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_61 
+ bl[59] br[59] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_62 
+ bl[60] br[60] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_63 
+ bl[61] br[61] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_64 
+ bl[62] br[62] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_65 
+ bl[63] br[63] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_66 
+ bl[64] br[64] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_67 
+ bl[65] br[65] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_68 
+ bl[66] br[66] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_69 
+ bl[67] br[67] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_70 
+ bl[68] br[68] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_71 
+ bl[69] br[69] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_72 
+ bl[70] br[70] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_73 
+ bl[71] br[71] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_74 
+ bl[72] br[72] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_75 
+ bl[73] br[73] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_76 
+ bl[74] br[74] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_77 
+ bl[75] br[75] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_78 
+ bl[76] br[76] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_79 
+ bl[77] br[77] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_80 
+ bl[78] br[78] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_81 
+ bl[79] br[79] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_82 
+ bl[80] br[80] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_83 
+ bl[81] br[81] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_84 
+ bl[82] br[82] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_85 
+ bl[83] br[83] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_86 
+ bl[84] br[84] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_87 
+ bl[85] br[85] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_88 
+ bl[86] br[86] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_89 
+ bl[87] br[87] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_90 
+ bl[88] br[88] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_91 
+ bl[89] br[89] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_92 
+ bl[90] br[90] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_93 
+ bl[91] br[91] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_94 
+ bl[92] br[92] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_95 
+ bl[93] br[93] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_96 
+ bl[94] br[94] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_97 
+ bl[95] br[95] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_98 
+ bl[96] br[96] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_99 
+ bl[97] br[97] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_100 
+ bl[98] br[98] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_101 
+ bl[99] br[99] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_102 
+ bl[100] br[100] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_103 
+ bl[101] br[101] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_104 
+ bl[102] br[102] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_105 
+ bl[103] br[103] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_106 
+ bl[104] br[104] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_107 
+ bl[105] br[105] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_108 
+ bl[106] br[106] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_109 
+ bl[107] br[107] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_110 
+ bl[108] br[108] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_111 
+ bl[109] br[109] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_112 
+ bl[110] br[110] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_113 
+ bl[111] br[111] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_114 
+ bl[112] br[112] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_115 
+ bl[113] br[113] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_116 
+ bl[114] br[114] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_117 
+ bl[115] br[115] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_118 
+ bl[116] br[116] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_119 
+ bl[117] br[117] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_120 
+ bl[118] br[118] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_121 
+ bl[119] br[119] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_122 
+ bl[120] br[120] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_123 
+ bl[121] br[121] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_124 
+ bl[122] br[122] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_125 
+ bl[123] br[123] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_126 
+ bl[124] br[124] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_127 
+ bl[125] br[125] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_128 
+ bl[126] br[126] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_129 
+ bl[127] br[127] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_130 
+ vdd vdd vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_131 
+ vdd vdd vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_0 
+ vdd vdd vss vdd vpb vnb wl[14] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_16_1 
+ rbl rbr vss vdd vpb vnb wl[14] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_16_2 
+ bl[0] br[0] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_3 
+ bl[1] br[1] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_4 
+ bl[2] br[2] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_5 
+ bl[3] br[3] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_6 
+ bl[4] br[4] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_7 
+ bl[5] br[5] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_8 
+ bl[6] br[6] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_9 
+ bl[7] br[7] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_10 
+ bl[8] br[8] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_11 
+ bl[9] br[9] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_12 
+ bl[10] br[10] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_13 
+ bl[11] br[11] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_14 
+ bl[12] br[12] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_15 
+ bl[13] br[13] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_16 
+ bl[14] br[14] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_17 
+ bl[15] br[15] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_18 
+ bl[16] br[16] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_19 
+ bl[17] br[17] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_20 
+ bl[18] br[18] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_21 
+ bl[19] br[19] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_22 
+ bl[20] br[20] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_23 
+ bl[21] br[21] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_24 
+ bl[22] br[22] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_25 
+ bl[23] br[23] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_26 
+ bl[24] br[24] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_27 
+ bl[25] br[25] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_28 
+ bl[26] br[26] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_29 
+ bl[27] br[27] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_30 
+ bl[28] br[28] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_31 
+ bl[29] br[29] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_32 
+ bl[30] br[30] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_33 
+ bl[31] br[31] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_34 
+ bl[32] br[32] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_35 
+ bl[33] br[33] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_36 
+ bl[34] br[34] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_37 
+ bl[35] br[35] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_38 
+ bl[36] br[36] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_39 
+ bl[37] br[37] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_40 
+ bl[38] br[38] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_41 
+ bl[39] br[39] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_42 
+ bl[40] br[40] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_43 
+ bl[41] br[41] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_44 
+ bl[42] br[42] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_45 
+ bl[43] br[43] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_46 
+ bl[44] br[44] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_47 
+ bl[45] br[45] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_48 
+ bl[46] br[46] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_49 
+ bl[47] br[47] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_50 
+ bl[48] br[48] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_51 
+ bl[49] br[49] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_52 
+ bl[50] br[50] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_53 
+ bl[51] br[51] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_54 
+ bl[52] br[52] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_55 
+ bl[53] br[53] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_56 
+ bl[54] br[54] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_57 
+ bl[55] br[55] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_58 
+ bl[56] br[56] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_59 
+ bl[57] br[57] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_60 
+ bl[58] br[58] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_61 
+ bl[59] br[59] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_62 
+ bl[60] br[60] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_63 
+ bl[61] br[61] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_64 
+ bl[62] br[62] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_65 
+ bl[63] br[63] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_66 
+ bl[64] br[64] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_67 
+ bl[65] br[65] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_68 
+ bl[66] br[66] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_69 
+ bl[67] br[67] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_70 
+ bl[68] br[68] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_71 
+ bl[69] br[69] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_72 
+ bl[70] br[70] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_73 
+ bl[71] br[71] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_74 
+ bl[72] br[72] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_75 
+ bl[73] br[73] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_76 
+ bl[74] br[74] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_77 
+ bl[75] br[75] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_78 
+ bl[76] br[76] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_79 
+ bl[77] br[77] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_80 
+ bl[78] br[78] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_81 
+ bl[79] br[79] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_82 
+ bl[80] br[80] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_83 
+ bl[81] br[81] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_84 
+ bl[82] br[82] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_85 
+ bl[83] br[83] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_86 
+ bl[84] br[84] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_87 
+ bl[85] br[85] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_88 
+ bl[86] br[86] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_89 
+ bl[87] br[87] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_90 
+ bl[88] br[88] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_91 
+ bl[89] br[89] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_92 
+ bl[90] br[90] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_93 
+ bl[91] br[91] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_94 
+ bl[92] br[92] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_95 
+ bl[93] br[93] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_96 
+ bl[94] br[94] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_97 
+ bl[95] br[95] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_98 
+ bl[96] br[96] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_99 
+ bl[97] br[97] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_100 
+ bl[98] br[98] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_101 
+ bl[99] br[99] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_102 
+ bl[100] br[100] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_103 
+ bl[101] br[101] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_104 
+ bl[102] br[102] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_105 
+ bl[103] br[103] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_106 
+ bl[104] br[104] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_107 
+ bl[105] br[105] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_108 
+ bl[106] br[106] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_109 
+ bl[107] br[107] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_110 
+ bl[108] br[108] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_111 
+ bl[109] br[109] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_112 
+ bl[110] br[110] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_113 
+ bl[111] br[111] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_114 
+ bl[112] br[112] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_115 
+ bl[113] br[113] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_116 
+ bl[114] br[114] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_117 
+ bl[115] br[115] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_118 
+ bl[116] br[116] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_119 
+ bl[117] br[117] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_120 
+ bl[118] br[118] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_121 
+ bl[119] br[119] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_122 
+ bl[120] br[120] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_123 
+ bl[121] br[121] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_124 
+ bl[122] br[122] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_125 
+ bl[123] br[123] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_126 
+ bl[124] br[124] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_127 
+ bl[125] br[125] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_128 
+ bl[126] br[126] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_129 
+ bl[127] br[127] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_130 
+ vdd vdd vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_131 
+ vdd vdd vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_0 
+ vdd vdd vss vdd vpb vnb wl[15] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_17_1 
+ rbl rbr vss vdd vpb vnb wl[15] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_17_2 
+ bl[0] br[0] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_3 
+ bl[1] br[1] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_4 
+ bl[2] br[2] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_5 
+ bl[3] br[3] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_6 
+ bl[4] br[4] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_7 
+ bl[5] br[5] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_8 
+ bl[6] br[6] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_9 
+ bl[7] br[7] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_10 
+ bl[8] br[8] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_11 
+ bl[9] br[9] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_12 
+ bl[10] br[10] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_13 
+ bl[11] br[11] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_14 
+ bl[12] br[12] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_15 
+ bl[13] br[13] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_16 
+ bl[14] br[14] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_17 
+ bl[15] br[15] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_18 
+ bl[16] br[16] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_19 
+ bl[17] br[17] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_20 
+ bl[18] br[18] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_21 
+ bl[19] br[19] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_22 
+ bl[20] br[20] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_23 
+ bl[21] br[21] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_24 
+ bl[22] br[22] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_25 
+ bl[23] br[23] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_26 
+ bl[24] br[24] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_27 
+ bl[25] br[25] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_28 
+ bl[26] br[26] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_29 
+ bl[27] br[27] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_30 
+ bl[28] br[28] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_31 
+ bl[29] br[29] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_32 
+ bl[30] br[30] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_33 
+ bl[31] br[31] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_34 
+ bl[32] br[32] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_35 
+ bl[33] br[33] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_36 
+ bl[34] br[34] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_37 
+ bl[35] br[35] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_38 
+ bl[36] br[36] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_39 
+ bl[37] br[37] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_40 
+ bl[38] br[38] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_41 
+ bl[39] br[39] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_42 
+ bl[40] br[40] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_43 
+ bl[41] br[41] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_44 
+ bl[42] br[42] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_45 
+ bl[43] br[43] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_46 
+ bl[44] br[44] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_47 
+ bl[45] br[45] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_48 
+ bl[46] br[46] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_49 
+ bl[47] br[47] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_50 
+ bl[48] br[48] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_51 
+ bl[49] br[49] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_52 
+ bl[50] br[50] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_53 
+ bl[51] br[51] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_54 
+ bl[52] br[52] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_55 
+ bl[53] br[53] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_56 
+ bl[54] br[54] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_57 
+ bl[55] br[55] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_58 
+ bl[56] br[56] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_59 
+ bl[57] br[57] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_60 
+ bl[58] br[58] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_61 
+ bl[59] br[59] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_62 
+ bl[60] br[60] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_63 
+ bl[61] br[61] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_64 
+ bl[62] br[62] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_65 
+ bl[63] br[63] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_66 
+ bl[64] br[64] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_67 
+ bl[65] br[65] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_68 
+ bl[66] br[66] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_69 
+ bl[67] br[67] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_70 
+ bl[68] br[68] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_71 
+ bl[69] br[69] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_72 
+ bl[70] br[70] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_73 
+ bl[71] br[71] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_74 
+ bl[72] br[72] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_75 
+ bl[73] br[73] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_76 
+ bl[74] br[74] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_77 
+ bl[75] br[75] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_78 
+ bl[76] br[76] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_79 
+ bl[77] br[77] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_80 
+ bl[78] br[78] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_81 
+ bl[79] br[79] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_82 
+ bl[80] br[80] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_83 
+ bl[81] br[81] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_84 
+ bl[82] br[82] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_85 
+ bl[83] br[83] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_86 
+ bl[84] br[84] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_87 
+ bl[85] br[85] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_88 
+ bl[86] br[86] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_89 
+ bl[87] br[87] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_90 
+ bl[88] br[88] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_91 
+ bl[89] br[89] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_92 
+ bl[90] br[90] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_93 
+ bl[91] br[91] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_94 
+ bl[92] br[92] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_95 
+ bl[93] br[93] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_96 
+ bl[94] br[94] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_97 
+ bl[95] br[95] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_98 
+ bl[96] br[96] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_99 
+ bl[97] br[97] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_100 
+ bl[98] br[98] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_101 
+ bl[99] br[99] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_102 
+ bl[100] br[100] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_103 
+ bl[101] br[101] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_104 
+ bl[102] br[102] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_105 
+ bl[103] br[103] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_106 
+ bl[104] br[104] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_107 
+ bl[105] br[105] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_108 
+ bl[106] br[106] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_109 
+ bl[107] br[107] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_110 
+ bl[108] br[108] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_111 
+ bl[109] br[109] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_112 
+ bl[110] br[110] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_113 
+ bl[111] br[111] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_114 
+ bl[112] br[112] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_115 
+ bl[113] br[113] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_116 
+ bl[114] br[114] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_117 
+ bl[115] br[115] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_118 
+ bl[116] br[116] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_119 
+ bl[117] br[117] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_120 
+ bl[118] br[118] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_121 
+ bl[119] br[119] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_122 
+ bl[120] br[120] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_123 
+ bl[121] br[121] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_124 
+ bl[122] br[122] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_125 
+ bl[123] br[123] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_126 
+ bl[124] br[124] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_127 
+ bl[125] br[125] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_128 
+ bl[126] br[126] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_129 
+ bl[127] br[127] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_130 
+ vdd vdd vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_131 
+ vdd vdd vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_0 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_1 
+ rbl rbr vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_2 
+ bl[0] br[0] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_3 
+ bl[1] br[1] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_4 
+ bl[2] br[2] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_5 
+ bl[3] br[3] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_6 
+ bl[4] br[4] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_7 
+ bl[5] br[5] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_8 
+ bl[6] br[6] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_9 
+ bl[7] br[7] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_10 
+ bl[8] br[8] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_11 
+ bl[9] br[9] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_12 
+ bl[10] br[10] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_13 
+ bl[11] br[11] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_14 
+ bl[12] br[12] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_15 
+ bl[13] br[13] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_16 
+ bl[14] br[14] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_17 
+ bl[15] br[15] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_18 
+ bl[16] br[16] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_19 
+ bl[17] br[17] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_20 
+ bl[18] br[18] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_21 
+ bl[19] br[19] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_22 
+ bl[20] br[20] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_23 
+ bl[21] br[21] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_24 
+ bl[22] br[22] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_25 
+ bl[23] br[23] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_26 
+ bl[24] br[24] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_27 
+ bl[25] br[25] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_28 
+ bl[26] br[26] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_29 
+ bl[27] br[27] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_30 
+ bl[28] br[28] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_31 
+ bl[29] br[29] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_32 
+ bl[30] br[30] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_33 
+ bl[31] br[31] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_34 
+ bl[32] br[32] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_35 
+ bl[33] br[33] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_36 
+ bl[34] br[34] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_37 
+ bl[35] br[35] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_38 
+ bl[36] br[36] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_39 
+ bl[37] br[37] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_40 
+ bl[38] br[38] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_41 
+ bl[39] br[39] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_42 
+ bl[40] br[40] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_43 
+ bl[41] br[41] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_44 
+ bl[42] br[42] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_45 
+ bl[43] br[43] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_46 
+ bl[44] br[44] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_47 
+ bl[45] br[45] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_48 
+ bl[46] br[46] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_49 
+ bl[47] br[47] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_50 
+ bl[48] br[48] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_51 
+ bl[49] br[49] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_52 
+ bl[50] br[50] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_53 
+ bl[51] br[51] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_54 
+ bl[52] br[52] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_55 
+ bl[53] br[53] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_56 
+ bl[54] br[54] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_57 
+ bl[55] br[55] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_58 
+ bl[56] br[56] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_59 
+ bl[57] br[57] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_60 
+ bl[58] br[58] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_61 
+ bl[59] br[59] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_62 
+ bl[60] br[60] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_63 
+ bl[61] br[61] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_64 
+ bl[62] br[62] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_65 
+ bl[63] br[63] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_66 
+ bl[64] br[64] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_67 
+ bl[65] br[65] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_68 
+ bl[66] br[66] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_69 
+ bl[67] br[67] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_70 
+ bl[68] br[68] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_71 
+ bl[69] br[69] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_72 
+ bl[70] br[70] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_73 
+ bl[71] br[71] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_74 
+ bl[72] br[72] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_75 
+ bl[73] br[73] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_76 
+ bl[74] br[74] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_77 
+ bl[75] br[75] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_78 
+ bl[76] br[76] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_79 
+ bl[77] br[77] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_80 
+ bl[78] br[78] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_81 
+ bl[79] br[79] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_82 
+ bl[80] br[80] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_83 
+ bl[81] br[81] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_84 
+ bl[82] br[82] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_85 
+ bl[83] br[83] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_86 
+ bl[84] br[84] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_87 
+ bl[85] br[85] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_88 
+ bl[86] br[86] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_89 
+ bl[87] br[87] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_90 
+ bl[88] br[88] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_91 
+ bl[89] br[89] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_92 
+ bl[90] br[90] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_93 
+ bl[91] br[91] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_94 
+ bl[92] br[92] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_95 
+ bl[93] br[93] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_96 
+ bl[94] br[94] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_97 
+ bl[95] br[95] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_98 
+ bl[96] br[96] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_99 
+ bl[97] br[97] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_100 
+ bl[98] br[98] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_101 
+ bl[99] br[99] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_102 
+ bl[100] br[100] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_103 
+ bl[101] br[101] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_104 
+ bl[102] br[102] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_105 
+ bl[103] br[103] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_106 
+ bl[104] br[104] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_107 
+ bl[105] br[105] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_108 
+ bl[106] br[106] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_109 
+ bl[107] br[107] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_110 
+ bl[108] br[108] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_111 
+ bl[109] br[109] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_112 
+ bl[110] br[110] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_113 
+ bl[111] br[111] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_114 
+ bl[112] br[112] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_115 
+ bl[113] br[113] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_116 
+ bl[114] br[114] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_117 
+ bl[115] br[115] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_118 
+ bl[116] br[116] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_119 
+ bl[117] br[117] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_120 
+ bl[118] br[118] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_121 
+ bl[119] br[119] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_122 
+ bl[120] br[120] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_123 
+ bl[121] br[121] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_124 
+ bl[122] br[122] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_125 
+ bl[123] br[123] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_126 
+ bl[124] br[124] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_127 
+ bl[125] br[125] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_128 
+ bl[126] br[126] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_129 
+ bl[127] br[127] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_130 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_131 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_0 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_1 
+ rbl rbr vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_2 
+ bl[0] br[0] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_3 
+ bl[1] br[1] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_4 
+ bl[2] br[2] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_5 
+ bl[3] br[3] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_6 
+ bl[4] br[4] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_7 
+ bl[5] br[5] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_8 
+ bl[6] br[6] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_9 
+ bl[7] br[7] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_10 
+ bl[8] br[8] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_11 
+ bl[9] br[9] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_12 
+ bl[10] br[10] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_13 
+ bl[11] br[11] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_14 
+ bl[12] br[12] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_15 
+ bl[13] br[13] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_16 
+ bl[14] br[14] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_17 
+ bl[15] br[15] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_18 
+ bl[16] br[16] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_19 
+ bl[17] br[17] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_20 
+ bl[18] br[18] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_21 
+ bl[19] br[19] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_22 
+ bl[20] br[20] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_23 
+ bl[21] br[21] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_24 
+ bl[22] br[22] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_25 
+ bl[23] br[23] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_26 
+ bl[24] br[24] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_27 
+ bl[25] br[25] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_28 
+ bl[26] br[26] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_29 
+ bl[27] br[27] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_30 
+ bl[28] br[28] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_31 
+ bl[29] br[29] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_32 
+ bl[30] br[30] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_33 
+ bl[31] br[31] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_34 
+ bl[32] br[32] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_35 
+ bl[33] br[33] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_36 
+ bl[34] br[34] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_37 
+ bl[35] br[35] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_38 
+ bl[36] br[36] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_39 
+ bl[37] br[37] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_40 
+ bl[38] br[38] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_41 
+ bl[39] br[39] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_42 
+ bl[40] br[40] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_43 
+ bl[41] br[41] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_44 
+ bl[42] br[42] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_45 
+ bl[43] br[43] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_46 
+ bl[44] br[44] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_47 
+ bl[45] br[45] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_48 
+ bl[46] br[46] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_49 
+ bl[47] br[47] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_50 
+ bl[48] br[48] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_51 
+ bl[49] br[49] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_52 
+ bl[50] br[50] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_53 
+ bl[51] br[51] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_54 
+ bl[52] br[52] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_55 
+ bl[53] br[53] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_56 
+ bl[54] br[54] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_57 
+ bl[55] br[55] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_58 
+ bl[56] br[56] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_59 
+ bl[57] br[57] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_60 
+ bl[58] br[58] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_61 
+ bl[59] br[59] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_62 
+ bl[60] br[60] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_63 
+ bl[61] br[61] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_64 
+ bl[62] br[62] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_65 
+ bl[63] br[63] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_66 
+ bl[64] br[64] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_67 
+ bl[65] br[65] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_68 
+ bl[66] br[66] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_69 
+ bl[67] br[67] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_70 
+ bl[68] br[68] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_71 
+ bl[69] br[69] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_72 
+ bl[70] br[70] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_73 
+ bl[71] br[71] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_74 
+ bl[72] br[72] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_75 
+ bl[73] br[73] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_76 
+ bl[74] br[74] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_77 
+ bl[75] br[75] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_78 
+ bl[76] br[76] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_79 
+ bl[77] br[77] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_80 
+ bl[78] br[78] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_81 
+ bl[79] br[79] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_82 
+ bl[80] br[80] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_83 
+ bl[81] br[81] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_84 
+ bl[82] br[82] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_85 
+ bl[83] br[83] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_86 
+ bl[84] br[84] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_87 
+ bl[85] br[85] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_88 
+ bl[86] br[86] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_89 
+ bl[87] br[87] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_90 
+ bl[88] br[88] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_91 
+ bl[89] br[89] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_92 
+ bl[90] br[90] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_93 
+ bl[91] br[91] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_94 
+ bl[92] br[92] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_95 
+ bl[93] br[93] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_96 
+ bl[94] br[94] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_97 
+ bl[95] br[95] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_98 
+ bl[96] br[96] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_99 
+ bl[97] br[97] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_100 
+ bl[98] br[98] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_101 
+ bl[99] br[99] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_102 
+ bl[100] br[100] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_103 
+ bl[101] br[101] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_104 
+ bl[102] br[102] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_105 
+ bl[103] br[103] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_106 
+ bl[104] br[104] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_107 
+ bl[105] br[105] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_108 
+ bl[106] br[106] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_109 
+ bl[107] br[107] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_110 
+ bl[108] br[108] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_111 
+ bl[109] br[109] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_112 
+ bl[110] br[110] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_113 
+ bl[111] br[111] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_114 
+ bl[112] br[112] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_115 
+ bl[113] br[113] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_116 
+ bl[114] br[114] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_117 
+ bl[115] br[115] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_118 
+ bl[116] br[116] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_119 
+ bl[117] br[117] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_120 
+ bl[118] br[118] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_121 
+ bl[119] br[119] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_122 
+ bl[120] br[120] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_123 
+ bl[121] br[121] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_124 
+ bl[122] br[122] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_125 
+ bl[123] br[123] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_126 
+ bl[124] br[124] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_127 
+ bl[125] br[125] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_128 
+ bl[126] br[126] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_129 
+ bl[127] br[127] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_130 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_131 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xcolend_0_bot 
+ vdd vdd vss vdd vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_0_top 
+ vdd vdd vss vdd vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_1_bot 
+ rbr vdd vss rbl vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_1_top 
+ rbr vdd vss rbl vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_2_bot 
+ br[0] vdd vss bl[0] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_2_top 
+ br[0] vdd vss bl[0] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_3_bot 
+ br[1] vdd vss bl[1] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_3_top 
+ br[1] vdd vss bl[1] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_4_bot 
+ br[2] vdd vss bl[2] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_4_top 
+ br[2] vdd vss bl[2] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_5_bot 
+ br[3] vdd vss bl[3] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_5_top 
+ br[3] vdd vss bl[3] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_6_bot 
+ br[4] vdd vss bl[4] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_6_top 
+ br[4] vdd vss bl[4] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_7_bot 
+ br[5] vdd vss bl[5] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_7_top 
+ br[5] vdd vss bl[5] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_8_bot 
+ br[6] vdd vss bl[6] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_8_top 
+ br[6] vdd vss bl[6] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_9_bot 
+ br[7] vdd vss bl[7] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_9_top 
+ br[7] vdd vss bl[7] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_10_bot 
+ br[8] vdd vss bl[8] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_10_top 
+ br[8] vdd vss bl[8] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_11_bot 
+ br[9] vdd vss bl[9] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_11_top 
+ br[9] vdd vss bl[9] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_12_bot 
+ br[10] vdd vss bl[10] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_12_top 
+ br[10] vdd vss bl[10] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_13_bot 
+ br[11] vdd vss bl[11] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_13_top 
+ br[11] vdd vss bl[11] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_14_bot 
+ br[12] vdd vss bl[12] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_14_top 
+ br[12] vdd vss bl[12] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_15_bot 
+ br[13] vdd vss bl[13] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_15_top 
+ br[13] vdd vss bl[13] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_16_bot 
+ br[14] vdd vss bl[14] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_16_top 
+ br[14] vdd vss bl[14] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_17_bot 
+ br[15] vdd vss bl[15] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_17_top 
+ br[15] vdd vss bl[15] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_18_bot 
+ br[16] vdd vss bl[16] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_18_top 
+ br[16] vdd vss bl[16] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_19_bot 
+ br[17] vdd vss bl[17] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_19_top 
+ br[17] vdd vss bl[17] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_20_bot 
+ br[18] vdd vss bl[18] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_20_top 
+ br[18] vdd vss bl[18] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_21_bot 
+ br[19] vdd vss bl[19] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_21_top 
+ br[19] vdd vss bl[19] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_22_bot 
+ br[20] vdd vss bl[20] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_22_top 
+ br[20] vdd vss bl[20] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_23_bot 
+ br[21] vdd vss bl[21] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_23_top 
+ br[21] vdd vss bl[21] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_24_bot 
+ br[22] vdd vss bl[22] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_24_top 
+ br[22] vdd vss bl[22] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_25_bot 
+ br[23] vdd vss bl[23] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_25_top 
+ br[23] vdd vss bl[23] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_26_bot 
+ br[24] vdd vss bl[24] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_26_top 
+ br[24] vdd vss bl[24] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_27_bot 
+ br[25] vdd vss bl[25] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_27_top 
+ br[25] vdd vss bl[25] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_28_bot 
+ br[26] vdd vss bl[26] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_28_top 
+ br[26] vdd vss bl[26] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_29_bot 
+ br[27] vdd vss bl[27] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_29_top 
+ br[27] vdd vss bl[27] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_30_bot 
+ br[28] vdd vss bl[28] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_30_top 
+ br[28] vdd vss bl[28] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_31_bot 
+ br[29] vdd vss bl[29] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_31_top 
+ br[29] vdd vss bl[29] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_32_bot 
+ br[30] vdd vss bl[30] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_32_top 
+ br[30] vdd vss bl[30] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_33_bot 
+ br[31] vdd vss bl[31] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_33_top 
+ br[31] vdd vss bl[31] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_34_bot 
+ br[32] vdd vss bl[32] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_34_top 
+ br[32] vdd vss bl[32] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_35_bot 
+ br[33] vdd vss bl[33] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_35_top 
+ br[33] vdd vss bl[33] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_36_bot 
+ br[34] vdd vss bl[34] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_36_top 
+ br[34] vdd vss bl[34] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_37_bot 
+ br[35] vdd vss bl[35] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_37_top 
+ br[35] vdd vss bl[35] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_38_bot 
+ br[36] vdd vss bl[36] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_38_top 
+ br[36] vdd vss bl[36] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_39_bot 
+ br[37] vdd vss bl[37] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_39_top 
+ br[37] vdd vss bl[37] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_40_bot 
+ br[38] vdd vss bl[38] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_40_top 
+ br[38] vdd vss bl[38] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_41_bot 
+ br[39] vdd vss bl[39] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_41_top 
+ br[39] vdd vss bl[39] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_42_bot 
+ br[40] vdd vss bl[40] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_42_top 
+ br[40] vdd vss bl[40] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_43_bot 
+ br[41] vdd vss bl[41] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_43_top 
+ br[41] vdd vss bl[41] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_44_bot 
+ br[42] vdd vss bl[42] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_44_top 
+ br[42] vdd vss bl[42] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_45_bot 
+ br[43] vdd vss bl[43] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_45_top 
+ br[43] vdd vss bl[43] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_46_bot 
+ br[44] vdd vss bl[44] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_46_top 
+ br[44] vdd vss bl[44] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_47_bot 
+ br[45] vdd vss bl[45] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_47_top 
+ br[45] vdd vss bl[45] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_48_bot 
+ br[46] vdd vss bl[46] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_48_top 
+ br[46] vdd vss bl[46] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_49_bot 
+ br[47] vdd vss bl[47] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_49_top 
+ br[47] vdd vss bl[47] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_50_bot 
+ br[48] vdd vss bl[48] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_50_top 
+ br[48] vdd vss bl[48] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_51_bot 
+ br[49] vdd vss bl[49] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_51_top 
+ br[49] vdd vss bl[49] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_52_bot 
+ br[50] vdd vss bl[50] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_52_top 
+ br[50] vdd vss bl[50] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_53_bot 
+ br[51] vdd vss bl[51] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_53_top 
+ br[51] vdd vss bl[51] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_54_bot 
+ br[52] vdd vss bl[52] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_54_top 
+ br[52] vdd vss bl[52] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_55_bot 
+ br[53] vdd vss bl[53] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_55_top 
+ br[53] vdd vss bl[53] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_56_bot 
+ br[54] vdd vss bl[54] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_56_top 
+ br[54] vdd vss bl[54] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_57_bot 
+ br[55] vdd vss bl[55] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_57_top 
+ br[55] vdd vss bl[55] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_58_bot 
+ br[56] vdd vss bl[56] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_58_top 
+ br[56] vdd vss bl[56] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_59_bot 
+ br[57] vdd vss bl[57] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_59_top 
+ br[57] vdd vss bl[57] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_60_bot 
+ br[58] vdd vss bl[58] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_60_top 
+ br[58] vdd vss bl[58] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_61_bot 
+ br[59] vdd vss bl[59] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_61_top 
+ br[59] vdd vss bl[59] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_62_bot 
+ br[60] vdd vss bl[60] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_62_top 
+ br[60] vdd vss bl[60] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_63_bot 
+ br[61] vdd vss bl[61] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_63_top 
+ br[61] vdd vss bl[61] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_64_bot 
+ br[62] vdd vss bl[62] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_64_top 
+ br[62] vdd vss bl[62] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_65_bot 
+ br[63] vdd vss bl[63] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_65_top 
+ br[63] vdd vss bl[63] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_66_bot 
+ br[64] vdd vss bl[64] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_66_top 
+ br[64] vdd vss bl[64] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_67_bot 
+ br[65] vdd vss bl[65] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_67_top 
+ br[65] vdd vss bl[65] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_68_bot 
+ br[66] vdd vss bl[66] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_68_top 
+ br[66] vdd vss bl[66] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_69_bot 
+ br[67] vdd vss bl[67] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_69_top 
+ br[67] vdd vss bl[67] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_70_bot 
+ br[68] vdd vss bl[68] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_70_top 
+ br[68] vdd vss bl[68] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_71_bot 
+ br[69] vdd vss bl[69] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_71_top 
+ br[69] vdd vss bl[69] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_72_bot 
+ br[70] vdd vss bl[70] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_72_top 
+ br[70] vdd vss bl[70] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_73_bot 
+ br[71] vdd vss bl[71] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_73_top 
+ br[71] vdd vss bl[71] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_74_bot 
+ br[72] vdd vss bl[72] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_74_top 
+ br[72] vdd vss bl[72] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_75_bot 
+ br[73] vdd vss bl[73] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_75_top 
+ br[73] vdd vss bl[73] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_76_bot 
+ br[74] vdd vss bl[74] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_76_top 
+ br[74] vdd vss bl[74] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_77_bot 
+ br[75] vdd vss bl[75] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_77_top 
+ br[75] vdd vss bl[75] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_78_bot 
+ br[76] vdd vss bl[76] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_78_top 
+ br[76] vdd vss bl[76] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_79_bot 
+ br[77] vdd vss bl[77] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_79_top 
+ br[77] vdd vss bl[77] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_80_bot 
+ br[78] vdd vss bl[78] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_80_top 
+ br[78] vdd vss bl[78] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_81_bot 
+ br[79] vdd vss bl[79] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_81_top 
+ br[79] vdd vss bl[79] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_82_bot 
+ br[80] vdd vss bl[80] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_82_top 
+ br[80] vdd vss bl[80] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_83_bot 
+ br[81] vdd vss bl[81] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_83_top 
+ br[81] vdd vss bl[81] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_84_bot 
+ br[82] vdd vss bl[82] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_84_top 
+ br[82] vdd vss bl[82] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_85_bot 
+ br[83] vdd vss bl[83] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_85_top 
+ br[83] vdd vss bl[83] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_86_bot 
+ br[84] vdd vss bl[84] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_86_top 
+ br[84] vdd vss bl[84] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_87_bot 
+ br[85] vdd vss bl[85] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_87_top 
+ br[85] vdd vss bl[85] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_88_bot 
+ br[86] vdd vss bl[86] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_88_top 
+ br[86] vdd vss bl[86] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_89_bot 
+ br[87] vdd vss bl[87] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_89_top 
+ br[87] vdd vss bl[87] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_90_bot 
+ br[88] vdd vss bl[88] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_90_top 
+ br[88] vdd vss bl[88] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_91_bot 
+ br[89] vdd vss bl[89] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_91_top 
+ br[89] vdd vss bl[89] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_92_bot 
+ br[90] vdd vss bl[90] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_92_top 
+ br[90] vdd vss bl[90] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_93_bot 
+ br[91] vdd vss bl[91] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_93_top 
+ br[91] vdd vss bl[91] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_94_bot 
+ br[92] vdd vss bl[92] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_94_top 
+ br[92] vdd vss bl[92] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_95_bot 
+ br[93] vdd vss bl[93] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_95_top 
+ br[93] vdd vss bl[93] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_96_bot 
+ br[94] vdd vss bl[94] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_96_top 
+ br[94] vdd vss bl[94] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_97_bot 
+ br[95] vdd vss bl[95] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_97_top 
+ br[95] vdd vss bl[95] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_98_bot 
+ br[96] vdd vss bl[96] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_98_top 
+ br[96] vdd vss bl[96] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_99_bot 
+ br[97] vdd vss bl[97] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_99_top 
+ br[97] vdd vss bl[97] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_100_bot 
+ br[98] vdd vss bl[98] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_100_top 
+ br[98] vdd vss bl[98] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_101_bot 
+ br[99] vdd vss bl[99] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_101_top 
+ br[99] vdd vss bl[99] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_102_bot 
+ br[100] vdd vss bl[100] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_102_top 
+ br[100] vdd vss bl[100] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_103_bot 
+ br[101] vdd vss bl[101] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_103_top 
+ br[101] vdd vss bl[101] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_104_bot 
+ br[102] vdd vss bl[102] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_104_top 
+ br[102] vdd vss bl[102] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_105_bot 
+ br[103] vdd vss bl[103] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_105_top 
+ br[103] vdd vss bl[103] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_106_bot 
+ br[104] vdd vss bl[104] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_106_top 
+ br[104] vdd vss bl[104] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_107_bot 
+ br[105] vdd vss bl[105] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_107_top 
+ br[105] vdd vss bl[105] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_108_bot 
+ br[106] vdd vss bl[106] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_108_top 
+ br[106] vdd vss bl[106] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_109_bot 
+ br[107] vdd vss bl[107] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_109_top 
+ br[107] vdd vss bl[107] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_110_bot 
+ br[108] vdd vss bl[108] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_110_top 
+ br[108] vdd vss bl[108] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_111_bot 
+ br[109] vdd vss bl[109] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_111_top 
+ br[109] vdd vss bl[109] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_112_bot 
+ br[110] vdd vss bl[110] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_112_top 
+ br[110] vdd vss bl[110] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_113_bot 
+ br[111] vdd vss bl[111] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_113_top 
+ br[111] vdd vss bl[111] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_114_bot 
+ br[112] vdd vss bl[112] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_114_top 
+ br[112] vdd vss bl[112] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_115_bot 
+ br[113] vdd vss bl[113] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_115_top 
+ br[113] vdd vss bl[113] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_116_bot 
+ br[114] vdd vss bl[114] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_116_top 
+ br[114] vdd vss bl[114] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_117_bot 
+ br[115] vdd vss bl[115] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_117_top 
+ br[115] vdd vss bl[115] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_118_bot 
+ br[116] vdd vss bl[116] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_118_top 
+ br[116] vdd vss bl[116] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_119_bot 
+ br[117] vdd vss bl[117] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_119_top 
+ br[117] vdd vss bl[117] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_120_bot 
+ br[118] vdd vss bl[118] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_120_top 
+ br[118] vdd vss bl[118] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_121_bot 
+ br[119] vdd vss bl[119] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_121_top 
+ br[119] vdd vss bl[119] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_122_bot 
+ br[120] vdd vss bl[120] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_122_top 
+ br[120] vdd vss bl[120] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_123_bot 
+ br[121] vdd vss bl[121] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_123_top 
+ br[121] vdd vss bl[121] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_124_bot 
+ br[122] vdd vss bl[122] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_124_top 
+ br[122] vdd vss bl[122] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_125_bot 
+ br[123] vdd vss bl[123] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_125_top 
+ br[123] vdd vss bl[123] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_126_bot 
+ br[124] vdd vss bl[124] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_126_top 
+ br[124] vdd vss bl[124] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_127_bot 
+ br[125] vdd vss bl[125] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_127_top 
+ br[125] vdd vss bl[125] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_128_bot 
+ br[126] vdd vss bl[126] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_128_top 
+ br[126] vdd vss bl[126] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_129_bot 
+ br[127] vdd vss bl[127] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_129_top 
+ br[127] vdd vss bl[127] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_130_bot 
+ vdd vdd vss vdd vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_130_top 
+ vdd vdd vss vdd vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_131_bot 
+ vdd vdd vss vdd vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_131_top 
+ vdd vdd vss vdd vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

.ENDS

.SUBCKT precharge 
+ vdd bl br en_b 

xbl_pull_up 
+ bl en_b vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='1.0' l='0.15' 

xbr_pull_up 
+ br en_b vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='1.0' l='0.15' 

xequalizer 
+ bl en_b br vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='1.0' l='0.15' 

.ENDS

.SUBCKT precharge_array 
+ vdd en_b bl[128] bl[127] bl[126] bl[125] bl[124] bl[123] bl[122] bl[121] bl[120] bl[119] bl[118] bl[117] bl[116] bl[115] bl[114] bl[113] bl[112] bl[111] bl[110] bl[109] bl[108] bl[107] bl[106] bl[105] bl[104] bl[103] bl[102] bl[101] bl[100] bl[99] bl[98] bl[97] bl[96] bl[95] bl[94] bl[93] bl[92] bl[91] bl[90] bl[89] bl[88] bl[87] bl[86] bl[85] bl[84] bl[83] bl[82] bl[81] bl[80] bl[79] bl[78] bl[77] bl[76] bl[75] bl[74] bl[73] bl[72] bl[71] bl[70] bl[69] bl[68] bl[67] bl[66] bl[65] bl[64] bl[63] bl[62] bl[61] bl[60] bl[59] bl[58] bl[57] bl[56] bl[55] bl[54] bl[53] bl[52] bl[51] bl[50] bl[49] bl[48] bl[47] bl[46] bl[45] bl[44] bl[43] bl[42] bl[41] bl[40] bl[39] bl[38] bl[37] bl[36] bl[35] bl[34] bl[33] bl[32] bl[31] bl[30] bl[29] bl[28] bl[27] bl[26] bl[25] bl[24] bl[23] bl[22] bl[21] bl[20] bl[19] bl[18] bl[17] bl[16] bl[15] bl[14] bl[13] bl[12] bl[11] bl[10] bl[9] bl[8] bl[7] bl[6] bl[5] bl[4] bl[3] bl[2] bl[1] bl[0] br[128] br[127] br[126] br[125] br[124] br[123] br[122] br[121] br[120] br[119] br[118] br[117] br[116] br[115] br[114] br[113] br[112] br[111] br[110] br[109] br[108] br[107] br[106] br[105] br[104] br[103] br[102] br[101] br[100] br[99] br[98] br[97] br[96] br[95] br[94] br[93] br[92] br[91] br[90] br[89] br[88] br[87] br[86] br[85] br[84] br[83] br[82] br[81] br[80] br[79] br[78] br[77] br[76] br[75] br[74] br[73] br[72] br[71] br[70] br[69] br[68] br[67] br[66] br[65] br[64] br[63] br[62] br[61] br[60] br[59] br[58] br[57] br[56] br[55] br[54] br[53] br[52] br[51] br[50] br[49] br[48] br[47] br[46] br[45] br[44] br[43] br[42] br[41] br[40] br[39] br[38] br[37] br[36] br[35] br[34] br[33] br[32] br[31] br[30] br[29] br[28] br[27] br[26] br[25] br[24] br[23] br[22] br[21] br[20] br[19] br[18] br[17] br[16] br[15] br[14] br[13] br[12] br[11] br[10] br[9] br[8] br[7] br[6] br[5] br[4] br[3] br[2] br[1] br[0] 

xprecharge_0 
+ vdd bl[0] br[0] en_b 
+ precharge 
* No parameters

xprecharge_1 
+ vdd bl[1] br[1] en_b 
+ precharge 
* No parameters

xprecharge_2 
+ vdd bl[2] br[2] en_b 
+ precharge 
* No parameters

xprecharge_3 
+ vdd bl[3] br[3] en_b 
+ precharge 
* No parameters

xprecharge_4 
+ vdd bl[4] br[4] en_b 
+ precharge 
* No parameters

xprecharge_5 
+ vdd bl[5] br[5] en_b 
+ precharge 
* No parameters

xprecharge_6 
+ vdd bl[6] br[6] en_b 
+ precharge 
* No parameters

xprecharge_7 
+ vdd bl[7] br[7] en_b 
+ precharge 
* No parameters

xprecharge_8 
+ vdd bl[8] br[8] en_b 
+ precharge 
* No parameters

xprecharge_9 
+ vdd bl[9] br[9] en_b 
+ precharge 
* No parameters

xprecharge_10 
+ vdd bl[10] br[10] en_b 
+ precharge 
* No parameters

xprecharge_11 
+ vdd bl[11] br[11] en_b 
+ precharge 
* No parameters

xprecharge_12 
+ vdd bl[12] br[12] en_b 
+ precharge 
* No parameters

xprecharge_13 
+ vdd bl[13] br[13] en_b 
+ precharge 
* No parameters

xprecharge_14 
+ vdd bl[14] br[14] en_b 
+ precharge 
* No parameters

xprecharge_15 
+ vdd bl[15] br[15] en_b 
+ precharge 
* No parameters

xprecharge_16 
+ vdd bl[16] br[16] en_b 
+ precharge 
* No parameters

xprecharge_17 
+ vdd bl[17] br[17] en_b 
+ precharge 
* No parameters

xprecharge_18 
+ vdd bl[18] br[18] en_b 
+ precharge 
* No parameters

xprecharge_19 
+ vdd bl[19] br[19] en_b 
+ precharge 
* No parameters

xprecharge_20 
+ vdd bl[20] br[20] en_b 
+ precharge 
* No parameters

xprecharge_21 
+ vdd bl[21] br[21] en_b 
+ precharge 
* No parameters

xprecharge_22 
+ vdd bl[22] br[22] en_b 
+ precharge 
* No parameters

xprecharge_23 
+ vdd bl[23] br[23] en_b 
+ precharge 
* No parameters

xprecharge_24 
+ vdd bl[24] br[24] en_b 
+ precharge 
* No parameters

xprecharge_25 
+ vdd bl[25] br[25] en_b 
+ precharge 
* No parameters

xprecharge_26 
+ vdd bl[26] br[26] en_b 
+ precharge 
* No parameters

xprecharge_27 
+ vdd bl[27] br[27] en_b 
+ precharge 
* No parameters

xprecharge_28 
+ vdd bl[28] br[28] en_b 
+ precharge 
* No parameters

xprecharge_29 
+ vdd bl[29] br[29] en_b 
+ precharge 
* No parameters

xprecharge_30 
+ vdd bl[30] br[30] en_b 
+ precharge 
* No parameters

xprecharge_31 
+ vdd bl[31] br[31] en_b 
+ precharge 
* No parameters

xprecharge_32 
+ vdd bl[32] br[32] en_b 
+ precharge 
* No parameters

xprecharge_33 
+ vdd bl[33] br[33] en_b 
+ precharge 
* No parameters

xprecharge_34 
+ vdd bl[34] br[34] en_b 
+ precharge 
* No parameters

xprecharge_35 
+ vdd bl[35] br[35] en_b 
+ precharge 
* No parameters

xprecharge_36 
+ vdd bl[36] br[36] en_b 
+ precharge 
* No parameters

xprecharge_37 
+ vdd bl[37] br[37] en_b 
+ precharge 
* No parameters

xprecharge_38 
+ vdd bl[38] br[38] en_b 
+ precharge 
* No parameters

xprecharge_39 
+ vdd bl[39] br[39] en_b 
+ precharge 
* No parameters

xprecharge_40 
+ vdd bl[40] br[40] en_b 
+ precharge 
* No parameters

xprecharge_41 
+ vdd bl[41] br[41] en_b 
+ precharge 
* No parameters

xprecharge_42 
+ vdd bl[42] br[42] en_b 
+ precharge 
* No parameters

xprecharge_43 
+ vdd bl[43] br[43] en_b 
+ precharge 
* No parameters

xprecharge_44 
+ vdd bl[44] br[44] en_b 
+ precharge 
* No parameters

xprecharge_45 
+ vdd bl[45] br[45] en_b 
+ precharge 
* No parameters

xprecharge_46 
+ vdd bl[46] br[46] en_b 
+ precharge 
* No parameters

xprecharge_47 
+ vdd bl[47] br[47] en_b 
+ precharge 
* No parameters

xprecharge_48 
+ vdd bl[48] br[48] en_b 
+ precharge 
* No parameters

xprecharge_49 
+ vdd bl[49] br[49] en_b 
+ precharge 
* No parameters

xprecharge_50 
+ vdd bl[50] br[50] en_b 
+ precharge 
* No parameters

xprecharge_51 
+ vdd bl[51] br[51] en_b 
+ precharge 
* No parameters

xprecharge_52 
+ vdd bl[52] br[52] en_b 
+ precharge 
* No parameters

xprecharge_53 
+ vdd bl[53] br[53] en_b 
+ precharge 
* No parameters

xprecharge_54 
+ vdd bl[54] br[54] en_b 
+ precharge 
* No parameters

xprecharge_55 
+ vdd bl[55] br[55] en_b 
+ precharge 
* No parameters

xprecharge_56 
+ vdd bl[56] br[56] en_b 
+ precharge 
* No parameters

xprecharge_57 
+ vdd bl[57] br[57] en_b 
+ precharge 
* No parameters

xprecharge_58 
+ vdd bl[58] br[58] en_b 
+ precharge 
* No parameters

xprecharge_59 
+ vdd bl[59] br[59] en_b 
+ precharge 
* No parameters

xprecharge_60 
+ vdd bl[60] br[60] en_b 
+ precharge 
* No parameters

xprecharge_61 
+ vdd bl[61] br[61] en_b 
+ precharge 
* No parameters

xprecharge_62 
+ vdd bl[62] br[62] en_b 
+ precharge 
* No parameters

xprecharge_63 
+ vdd bl[63] br[63] en_b 
+ precharge 
* No parameters

xprecharge_64 
+ vdd bl[64] br[64] en_b 
+ precharge 
* No parameters

xprecharge_65 
+ vdd bl[65] br[65] en_b 
+ precharge 
* No parameters

xprecharge_66 
+ vdd bl[66] br[66] en_b 
+ precharge 
* No parameters

xprecharge_67 
+ vdd bl[67] br[67] en_b 
+ precharge 
* No parameters

xprecharge_68 
+ vdd bl[68] br[68] en_b 
+ precharge 
* No parameters

xprecharge_69 
+ vdd bl[69] br[69] en_b 
+ precharge 
* No parameters

xprecharge_70 
+ vdd bl[70] br[70] en_b 
+ precharge 
* No parameters

xprecharge_71 
+ vdd bl[71] br[71] en_b 
+ precharge 
* No parameters

xprecharge_72 
+ vdd bl[72] br[72] en_b 
+ precharge 
* No parameters

xprecharge_73 
+ vdd bl[73] br[73] en_b 
+ precharge 
* No parameters

xprecharge_74 
+ vdd bl[74] br[74] en_b 
+ precharge 
* No parameters

xprecharge_75 
+ vdd bl[75] br[75] en_b 
+ precharge 
* No parameters

xprecharge_76 
+ vdd bl[76] br[76] en_b 
+ precharge 
* No parameters

xprecharge_77 
+ vdd bl[77] br[77] en_b 
+ precharge 
* No parameters

xprecharge_78 
+ vdd bl[78] br[78] en_b 
+ precharge 
* No parameters

xprecharge_79 
+ vdd bl[79] br[79] en_b 
+ precharge 
* No parameters

xprecharge_80 
+ vdd bl[80] br[80] en_b 
+ precharge 
* No parameters

xprecharge_81 
+ vdd bl[81] br[81] en_b 
+ precharge 
* No parameters

xprecharge_82 
+ vdd bl[82] br[82] en_b 
+ precharge 
* No parameters

xprecharge_83 
+ vdd bl[83] br[83] en_b 
+ precharge 
* No parameters

xprecharge_84 
+ vdd bl[84] br[84] en_b 
+ precharge 
* No parameters

xprecharge_85 
+ vdd bl[85] br[85] en_b 
+ precharge 
* No parameters

xprecharge_86 
+ vdd bl[86] br[86] en_b 
+ precharge 
* No parameters

xprecharge_87 
+ vdd bl[87] br[87] en_b 
+ precharge 
* No parameters

xprecharge_88 
+ vdd bl[88] br[88] en_b 
+ precharge 
* No parameters

xprecharge_89 
+ vdd bl[89] br[89] en_b 
+ precharge 
* No parameters

xprecharge_90 
+ vdd bl[90] br[90] en_b 
+ precharge 
* No parameters

xprecharge_91 
+ vdd bl[91] br[91] en_b 
+ precharge 
* No parameters

xprecharge_92 
+ vdd bl[92] br[92] en_b 
+ precharge 
* No parameters

xprecharge_93 
+ vdd bl[93] br[93] en_b 
+ precharge 
* No parameters

xprecharge_94 
+ vdd bl[94] br[94] en_b 
+ precharge 
* No parameters

xprecharge_95 
+ vdd bl[95] br[95] en_b 
+ precharge 
* No parameters

xprecharge_96 
+ vdd bl[96] br[96] en_b 
+ precharge 
* No parameters

xprecharge_97 
+ vdd bl[97] br[97] en_b 
+ precharge 
* No parameters

xprecharge_98 
+ vdd bl[98] br[98] en_b 
+ precharge 
* No parameters

xprecharge_99 
+ vdd bl[99] br[99] en_b 
+ precharge 
* No parameters

xprecharge_100 
+ vdd bl[100] br[100] en_b 
+ precharge 
* No parameters

xprecharge_101 
+ vdd bl[101] br[101] en_b 
+ precharge 
* No parameters

xprecharge_102 
+ vdd bl[102] br[102] en_b 
+ precharge 
* No parameters

xprecharge_103 
+ vdd bl[103] br[103] en_b 
+ precharge 
* No parameters

xprecharge_104 
+ vdd bl[104] br[104] en_b 
+ precharge 
* No parameters

xprecharge_105 
+ vdd bl[105] br[105] en_b 
+ precharge 
* No parameters

xprecharge_106 
+ vdd bl[106] br[106] en_b 
+ precharge 
* No parameters

xprecharge_107 
+ vdd bl[107] br[107] en_b 
+ precharge 
* No parameters

xprecharge_108 
+ vdd bl[108] br[108] en_b 
+ precharge 
* No parameters

xprecharge_109 
+ vdd bl[109] br[109] en_b 
+ precharge 
* No parameters

xprecharge_110 
+ vdd bl[110] br[110] en_b 
+ precharge 
* No parameters

xprecharge_111 
+ vdd bl[111] br[111] en_b 
+ precharge 
* No parameters

xprecharge_112 
+ vdd bl[112] br[112] en_b 
+ precharge 
* No parameters

xprecharge_113 
+ vdd bl[113] br[113] en_b 
+ precharge 
* No parameters

xprecharge_114 
+ vdd bl[114] br[114] en_b 
+ precharge 
* No parameters

xprecharge_115 
+ vdd bl[115] br[115] en_b 
+ precharge 
* No parameters

xprecharge_116 
+ vdd bl[116] br[116] en_b 
+ precharge 
* No parameters

xprecharge_117 
+ vdd bl[117] br[117] en_b 
+ precharge 
* No parameters

xprecharge_118 
+ vdd bl[118] br[118] en_b 
+ precharge 
* No parameters

xprecharge_119 
+ vdd bl[119] br[119] en_b 
+ precharge 
* No parameters

xprecharge_120 
+ vdd bl[120] br[120] en_b 
+ precharge 
* No parameters

xprecharge_121 
+ vdd bl[121] br[121] en_b 
+ precharge 
* No parameters

xprecharge_122 
+ vdd bl[122] br[122] en_b 
+ precharge 
* No parameters

xprecharge_123 
+ vdd bl[123] br[123] en_b 
+ precharge 
* No parameters

xprecharge_124 
+ vdd bl[124] br[124] en_b 
+ precharge 
* No parameters

xprecharge_125 
+ vdd bl[125] br[125] en_b 
+ precharge 
* No parameters

xprecharge_126 
+ vdd bl[126] br[126] en_b 
+ precharge 
* No parameters

xprecharge_127 
+ vdd bl[127] br[127] en_b 
+ precharge 
* No parameters

xprecharge_128 
+ vdd bl[128] br[128] en_b 
+ precharge 
* No parameters

.ENDS

.SUBCKT read_mux 
+ sel_b bl br bl_out br_out vdd 

xMBL 
+ bl_out sel_b bl vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='1.2' l='0.15' 

xMBR 
+ br_out sel_b br vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='1.2' l='0.15' 

.ENDS

.SUBCKT read_mux_array 
+ sel_b[3] sel_b[2] sel_b[1] sel_b[0] bl[127] bl[126] bl[125] bl[124] bl[123] bl[122] bl[121] bl[120] bl[119] bl[118] bl[117] bl[116] bl[115] bl[114] bl[113] bl[112] bl[111] bl[110] bl[109] bl[108] bl[107] bl[106] bl[105] bl[104] bl[103] bl[102] bl[101] bl[100] bl[99] bl[98] bl[97] bl[96] bl[95] bl[94] bl[93] bl[92] bl[91] bl[90] bl[89] bl[88] bl[87] bl[86] bl[85] bl[84] bl[83] bl[82] bl[81] bl[80] bl[79] bl[78] bl[77] bl[76] bl[75] bl[74] bl[73] bl[72] bl[71] bl[70] bl[69] bl[68] bl[67] bl[66] bl[65] bl[64] bl[63] bl[62] bl[61] bl[60] bl[59] bl[58] bl[57] bl[56] bl[55] bl[54] bl[53] bl[52] bl[51] bl[50] bl[49] bl[48] bl[47] bl[46] bl[45] bl[44] bl[43] bl[42] bl[41] bl[40] bl[39] bl[38] bl[37] bl[36] bl[35] bl[34] bl[33] bl[32] bl[31] bl[30] bl[29] bl[28] bl[27] bl[26] bl[25] bl[24] bl[23] bl[22] bl[21] bl[20] bl[19] bl[18] bl[17] bl[16] bl[15] bl[14] bl[13] bl[12] bl[11] bl[10] bl[9] bl[8] bl[7] bl[6] bl[5] bl[4] bl[3] bl[2] bl[1] bl[0] br[127] br[126] br[125] br[124] br[123] br[122] br[121] br[120] br[119] br[118] br[117] br[116] br[115] br[114] br[113] br[112] br[111] br[110] br[109] br[108] br[107] br[106] br[105] br[104] br[103] br[102] br[101] br[100] br[99] br[98] br[97] br[96] br[95] br[94] br[93] br[92] br[91] br[90] br[89] br[88] br[87] br[86] br[85] br[84] br[83] br[82] br[81] br[80] br[79] br[78] br[77] br[76] br[75] br[74] br[73] br[72] br[71] br[70] br[69] br[68] br[67] br[66] br[65] br[64] br[63] br[62] br[61] br[60] br[59] br[58] br[57] br[56] br[55] br[54] br[53] br[52] br[51] br[50] br[49] br[48] br[47] br[46] br[45] br[44] br[43] br[42] br[41] br[40] br[39] br[38] br[37] br[36] br[35] br[34] br[33] br[32] br[31] br[30] br[29] br[28] br[27] br[26] br[25] br[24] br[23] br[22] br[21] br[20] br[19] br[18] br[17] br[16] br[15] br[14] br[13] br[12] br[11] br[10] br[9] br[8] br[7] br[6] br[5] br[4] br[3] br[2] br[1] br[0] bl_out[31] bl_out[30] bl_out[29] bl_out[28] bl_out[27] bl_out[26] bl_out[25] bl_out[24] bl_out[23] bl_out[22] bl_out[21] bl_out[20] bl_out[19] bl_out[18] bl_out[17] bl_out[16] bl_out[15] bl_out[14] bl_out[13] bl_out[12] bl_out[11] bl_out[10] bl_out[9] bl_out[8] bl_out[7] bl_out[6] bl_out[5] bl_out[4] bl_out[3] bl_out[2] bl_out[1] bl_out[0] br_out[31] br_out[30] br_out[29] br_out[28] br_out[27] br_out[26] br_out[25] br_out[24] br_out[23] br_out[22] br_out[21] br_out[20] br_out[19] br_out[18] br_out[17] br_out[16] br_out[15] br_out[14] br_out[13] br_out[12] br_out[11] br_out[10] br_out[9] br_out[8] br_out[7] br_out[6] br_out[5] br_out[4] br_out[3] br_out[2] br_out[1] br_out[0] vdd 

xmux_0 
+ sel_b[0] bl[0] br[0] bl_out[0] br_out[0] vdd 
+ read_mux 
* No parameters

xmux_1 
+ sel_b[1] bl[1] br[1] bl_out[0] br_out[0] vdd 
+ read_mux 
* No parameters

xmux_2 
+ sel_b[2] bl[2] br[2] bl_out[0] br_out[0] vdd 
+ read_mux 
* No parameters

xmux_3 
+ sel_b[3] bl[3] br[3] bl_out[0] br_out[0] vdd 
+ read_mux 
* No parameters

xmux_4 
+ sel_b[0] bl[4] br[4] bl_out[1] br_out[1] vdd 
+ read_mux 
* No parameters

xmux_5 
+ sel_b[1] bl[5] br[5] bl_out[1] br_out[1] vdd 
+ read_mux 
* No parameters

xmux_6 
+ sel_b[2] bl[6] br[6] bl_out[1] br_out[1] vdd 
+ read_mux 
* No parameters

xmux_7 
+ sel_b[3] bl[7] br[7] bl_out[1] br_out[1] vdd 
+ read_mux 
* No parameters

xmux_8 
+ sel_b[0] bl[8] br[8] bl_out[2] br_out[2] vdd 
+ read_mux 
* No parameters

xmux_9 
+ sel_b[1] bl[9] br[9] bl_out[2] br_out[2] vdd 
+ read_mux 
* No parameters

xmux_10 
+ sel_b[2] bl[10] br[10] bl_out[2] br_out[2] vdd 
+ read_mux 
* No parameters

xmux_11 
+ sel_b[3] bl[11] br[11] bl_out[2] br_out[2] vdd 
+ read_mux 
* No parameters

xmux_12 
+ sel_b[0] bl[12] br[12] bl_out[3] br_out[3] vdd 
+ read_mux 
* No parameters

xmux_13 
+ sel_b[1] bl[13] br[13] bl_out[3] br_out[3] vdd 
+ read_mux 
* No parameters

xmux_14 
+ sel_b[2] bl[14] br[14] bl_out[3] br_out[3] vdd 
+ read_mux 
* No parameters

xmux_15 
+ sel_b[3] bl[15] br[15] bl_out[3] br_out[3] vdd 
+ read_mux 
* No parameters

xmux_16 
+ sel_b[0] bl[16] br[16] bl_out[4] br_out[4] vdd 
+ read_mux 
* No parameters

xmux_17 
+ sel_b[1] bl[17] br[17] bl_out[4] br_out[4] vdd 
+ read_mux 
* No parameters

xmux_18 
+ sel_b[2] bl[18] br[18] bl_out[4] br_out[4] vdd 
+ read_mux 
* No parameters

xmux_19 
+ sel_b[3] bl[19] br[19] bl_out[4] br_out[4] vdd 
+ read_mux 
* No parameters

xmux_20 
+ sel_b[0] bl[20] br[20] bl_out[5] br_out[5] vdd 
+ read_mux 
* No parameters

xmux_21 
+ sel_b[1] bl[21] br[21] bl_out[5] br_out[5] vdd 
+ read_mux 
* No parameters

xmux_22 
+ sel_b[2] bl[22] br[22] bl_out[5] br_out[5] vdd 
+ read_mux 
* No parameters

xmux_23 
+ sel_b[3] bl[23] br[23] bl_out[5] br_out[5] vdd 
+ read_mux 
* No parameters

xmux_24 
+ sel_b[0] bl[24] br[24] bl_out[6] br_out[6] vdd 
+ read_mux 
* No parameters

xmux_25 
+ sel_b[1] bl[25] br[25] bl_out[6] br_out[6] vdd 
+ read_mux 
* No parameters

xmux_26 
+ sel_b[2] bl[26] br[26] bl_out[6] br_out[6] vdd 
+ read_mux 
* No parameters

xmux_27 
+ sel_b[3] bl[27] br[27] bl_out[6] br_out[6] vdd 
+ read_mux 
* No parameters

xmux_28 
+ sel_b[0] bl[28] br[28] bl_out[7] br_out[7] vdd 
+ read_mux 
* No parameters

xmux_29 
+ sel_b[1] bl[29] br[29] bl_out[7] br_out[7] vdd 
+ read_mux 
* No parameters

xmux_30 
+ sel_b[2] bl[30] br[30] bl_out[7] br_out[7] vdd 
+ read_mux 
* No parameters

xmux_31 
+ sel_b[3] bl[31] br[31] bl_out[7] br_out[7] vdd 
+ read_mux 
* No parameters

xmux_32 
+ sel_b[0] bl[32] br[32] bl_out[8] br_out[8] vdd 
+ read_mux 
* No parameters

xmux_33 
+ sel_b[1] bl[33] br[33] bl_out[8] br_out[8] vdd 
+ read_mux 
* No parameters

xmux_34 
+ sel_b[2] bl[34] br[34] bl_out[8] br_out[8] vdd 
+ read_mux 
* No parameters

xmux_35 
+ sel_b[3] bl[35] br[35] bl_out[8] br_out[8] vdd 
+ read_mux 
* No parameters

xmux_36 
+ sel_b[0] bl[36] br[36] bl_out[9] br_out[9] vdd 
+ read_mux 
* No parameters

xmux_37 
+ sel_b[1] bl[37] br[37] bl_out[9] br_out[9] vdd 
+ read_mux 
* No parameters

xmux_38 
+ sel_b[2] bl[38] br[38] bl_out[9] br_out[9] vdd 
+ read_mux 
* No parameters

xmux_39 
+ sel_b[3] bl[39] br[39] bl_out[9] br_out[9] vdd 
+ read_mux 
* No parameters

xmux_40 
+ sel_b[0] bl[40] br[40] bl_out[10] br_out[10] vdd 
+ read_mux 
* No parameters

xmux_41 
+ sel_b[1] bl[41] br[41] bl_out[10] br_out[10] vdd 
+ read_mux 
* No parameters

xmux_42 
+ sel_b[2] bl[42] br[42] bl_out[10] br_out[10] vdd 
+ read_mux 
* No parameters

xmux_43 
+ sel_b[3] bl[43] br[43] bl_out[10] br_out[10] vdd 
+ read_mux 
* No parameters

xmux_44 
+ sel_b[0] bl[44] br[44] bl_out[11] br_out[11] vdd 
+ read_mux 
* No parameters

xmux_45 
+ sel_b[1] bl[45] br[45] bl_out[11] br_out[11] vdd 
+ read_mux 
* No parameters

xmux_46 
+ sel_b[2] bl[46] br[46] bl_out[11] br_out[11] vdd 
+ read_mux 
* No parameters

xmux_47 
+ sel_b[3] bl[47] br[47] bl_out[11] br_out[11] vdd 
+ read_mux 
* No parameters

xmux_48 
+ sel_b[0] bl[48] br[48] bl_out[12] br_out[12] vdd 
+ read_mux 
* No parameters

xmux_49 
+ sel_b[1] bl[49] br[49] bl_out[12] br_out[12] vdd 
+ read_mux 
* No parameters

xmux_50 
+ sel_b[2] bl[50] br[50] bl_out[12] br_out[12] vdd 
+ read_mux 
* No parameters

xmux_51 
+ sel_b[3] bl[51] br[51] bl_out[12] br_out[12] vdd 
+ read_mux 
* No parameters

xmux_52 
+ sel_b[0] bl[52] br[52] bl_out[13] br_out[13] vdd 
+ read_mux 
* No parameters

xmux_53 
+ sel_b[1] bl[53] br[53] bl_out[13] br_out[13] vdd 
+ read_mux 
* No parameters

xmux_54 
+ sel_b[2] bl[54] br[54] bl_out[13] br_out[13] vdd 
+ read_mux 
* No parameters

xmux_55 
+ sel_b[3] bl[55] br[55] bl_out[13] br_out[13] vdd 
+ read_mux 
* No parameters

xmux_56 
+ sel_b[0] bl[56] br[56] bl_out[14] br_out[14] vdd 
+ read_mux 
* No parameters

xmux_57 
+ sel_b[1] bl[57] br[57] bl_out[14] br_out[14] vdd 
+ read_mux 
* No parameters

xmux_58 
+ sel_b[2] bl[58] br[58] bl_out[14] br_out[14] vdd 
+ read_mux 
* No parameters

xmux_59 
+ sel_b[3] bl[59] br[59] bl_out[14] br_out[14] vdd 
+ read_mux 
* No parameters

xmux_60 
+ sel_b[0] bl[60] br[60] bl_out[15] br_out[15] vdd 
+ read_mux 
* No parameters

xmux_61 
+ sel_b[1] bl[61] br[61] bl_out[15] br_out[15] vdd 
+ read_mux 
* No parameters

xmux_62 
+ sel_b[2] bl[62] br[62] bl_out[15] br_out[15] vdd 
+ read_mux 
* No parameters

xmux_63 
+ sel_b[3] bl[63] br[63] bl_out[15] br_out[15] vdd 
+ read_mux 
* No parameters

xmux_64 
+ sel_b[0] bl[64] br[64] bl_out[16] br_out[16] vdd 
+ read_mux 
* No parameters

xmux_65 
+ sel_b[1] bl[65] br[65] bl_out[16] br_out[16] vdd 
+ read_mux 
* No parameters

xmux_66 
+ sel_b[2] bl[66] br[66] bl_out[16] br_out[16] vdd 
+ read_mux 
* No parameters

xmux_67 
+ sel_b[3] bl[67] br[67] bl_out[16] br_out[16] vdd 
+ read_mux 
* No parameters

xmux_68 
+ sel_b[0] bl[68] br[68] bl_out[17] br_out[17] vdd 
+ read_mux 
* No parameters

xmux_69 
+ sel_b[1] bl[69] br[69] bl_out[17] br_out[17] vdd 
+ read_mux 
* No parameters

xmux_70 
+ sel_b[2] bl[70] br[70] bl_out[17] br_out[17] vdd 
+ read_mux 
* No parameters

xmux_71 
+ sel_b[3] bl[71] br[71] bl_out[17] br_out[17] vdd 
+ read_mux 
* No parameters

xmux_72 
+ sel_b[0] bl[72] br[72] bl_out[18] br_out[18] vdd 
+ read_mux 
* No parameters

xmux_73 
+ sel_b[1] bl[73] br[73] bl_out[18] br_out[18] vdd 
+ read_mux 
* No parameters

xmux_74 
+ sel_b[2] bl[74] br[74] bl_out[18] br_out[18] vdd 
+ read_mux 
* No parameters

xmux_75 
+ sel_b[3] bl[75] br[75] bl_out[18] br_out[18] vdd 
+ read_mux 
* No parameters

xmux_76 
+ sel_b[0] bl[76] br[76] bl_out[19] br_out[19] vdd 
+ read_mux 
* No parameters

xmux_77 
+ sel_b[1] bl[77] br[77] bl_out[19] br_out[19] vdd 
+ read_mux 
* No parameters

xmux_78 
+ sel_b[2] bl[78] br[78] bl_out[19] br_out[19] vdd 
+ read_mux 
* No parameters

xmux_79 
+ sel_b[3] bl[79] br[79] bl_out[19] br_out[19] vdd 
+ read_mux 
* No parameters

xmux_80 
+ sel_b[0] bl[80] br[80] bl_out[20] br_out[20] vdd 
+ read_mux 
* No parameters

xmux_81 
+ sel_b[1] bl[81] br[81] bl_out[20] br_out[20] vdd 
+ read_mux 
* No parameters

xmux_82 
+ sel_b[2] bl[82] br[82] bl_out[20] br_out[20] vdd 
+ read_mux 
* No parameters

xmux_83 
+ sel_b[3] bl[83] br[83] bl_out[20] br_out[20] vdd 
+ read_mux 
* No parameters

xmux_84 
+ sel_b[0] bl[84] br[84] bl_out[21] br_out[21] vdd 
+ read_mux 
* No parameters

xmux_85 
+ sel_b[1] bl[85] br[85] bl_out[21] br_out[21] vdd 
+ read_mux 
* No parameters

xmux_86 
+ sel_b[2] bl[86] br[86] bl_out[21] br_out[21] vdd 
+ read_mux 
* No parameters

xmux_87 
+ sel_b[3] bl[87] br[87] bl_out[21] br_out[21] vdd 
+ read_mux 
* No parameters

xmux_88 
+ sel_b[0] bl[88] br[88] bl_out[22] br_out[22] vdd 
+ read_mux 
* No parameters

xmux_89 
+ sel_b[1] bl[89] br[89] bl_out[22] br_out[22] vdd 
+ read_mux 
* No parameters

xmux_90 
+ sel_b[2] bl[90] br[90] bl_out[22] br_out[22] vdd 
+ read_mux 
* No parameters

xmux_91 
+ sel_b[3] bl[91] br[91] bl_out[22] br_out[22] vdd 
+ read_mux 
* No parameters

xmux_92 
+ sel_b[0] bl[92] br[92] bl_out[23] br_out[23] vdd 
+ read_mux 
* No parameters

xmux_93 
+ sel_b[1] bl[93] br[93] bl_out[23] br_out[23] vdd 
+ read_mux 
* No parameters

xmux_94 
+ sel_b[2] bl[94] br[94] bl_out[23] br_out[23] vdd 
+ read_mux 
* No parameters

xmux_95 
+ sel_b[3] bl[95] br[95] bl_out[23] br_out[23] vdd 
+ read_mux 
* No parameters

xmux_96 
+ sel_b[0] bl[96] br[96] bl_out[24] br_out[24] vdd 
+ read_mux 
* No parameters

xmux_97 
+ sel_b[1] bl[97] br[97] bl_out[24] br_out[24] vdd 
+ read_mux 
* No parameters

xmux_98 
+ sel_b[2] bl[98] br[98] bl_out[24] br_out[24] vdd 
+ read_mux 
* No parameters

xmux_99 
+ sel_b[3] bl[99] br[99] bl_out[24] br_out[24] vdd 
+ read_mux 
* No parameters

xmux_100 
+ sel_b[0] bl[100] br[100] bl_out[25] br_out[25] vdd 
+ read_mux 
* No parameters

xmux_101 
+ sel_b[1] bl[101] br[101] bl_out[25] br_out[25] vdd 
+ read_mux 
* No parameters

xmux_102 
+ sel_b[2] bl[102] br[102] bl_out[25] br_out[25] vdd 
+ read_mux 
* No parameters

xmux_103 
+ sel_b[3] bl[103] br[103] bl_out[25] br_out[25] vdd 
+ read_mux 
* No parameters

xmux_104 
+ sel_b[0] bl[104] br[104] bl_out[26] br_out[26] vdd 
+ read_mux 
* No parameters

xmux_105 
+ sel_b[1] bl[105] br[105] bl_out[26] br_out[26] vdd 
+ read_mux 
* No parameters

xmux_106 
+ sel_b[2] bl[106] br[106] bl_out[26] br_out[26] vdd 
+ read_mux 
* No parameters

xmux_107 
+ sel_b[3] bl[107] br[107] bl_out[26] br_out[26] vdd 
+ read_mux 
* No parameters

xmux_108 
+ sel_b[0] bl[108] br[108] bl_out[27] br_out[27] vdd 
+ read_mux 
* No parameters

xmux_109 
+ sel_b[1] bl[109] br[109] bl_out[27] br_out[27] vdd 
+ read_mux 
* No parameters

xmux_110 
+ sel_b[2] bl[110] br[110] bl_out[27] br_out[27] vdd 
+ read_mux 
* No parameters

xmux_111 
+ sel_b[3] bl[111] br[111] bl_out[27] br_out[27] vdd 
+ read_mux 
* No parameters

xmux_112 
+ sel_b[0] bl[112] br[112] bl_out[28] br_out[28] vdd 
+ read_mux 
* No parameters

xmux_113 
+ sel_b[1] bl[113] br[113] bl_out[28] br_out[28] vdd 
+ read_mux 
* No parameters

xmux_114 
+ sel_b[2] bl[114] br[114] bl_out[28] br_out[28] vdd 
+ read_mux 
* No parameters

xmux_115 
+ sel_b[3] bl[115] br[115] bl_out[28] br_out[28] vdd 
+ read_mux 
* No parameters

xmux_116 
+ sel_b[0] bl[116] br[116] bl_out[29] br_out[29] vdd 
+ read_mux 
* No parameters

xmux_117 
+ sel_b[1] bl[117] br[117] bl_out[29] br_out[29] vdd 
+ read_mux 
* No parameters

xmux_118 
+ sel_b[2] bl[118] br[118] bl_out[29] br_out[29] vdd 
+ read_mux 
* No parameters

xmux_119 
+ sel_b[3] bl[119] br[119] bl_out[29] br_out[29] vdd 
+ read_mux 
* No parameters

xmux_120 
+ sel_b[0] bl[120] br[120] bl_out[30] br_out[30] vdd 
+ read_mux 
* No parameters

xmux_121 
+ sel_b[1] bl[121] br[121] bl_out[30] br_out[30] vdd 
+ read_mux 
* No parameters

xmux_122 
+ sel_b[2] bl[122] br[122] bl_out[30] br_out[30] vdd 
+ read_mux 
* No parameters

xmux_123 
+ sel_b[3] bl[123] br[123] bl_out[30] br_out[30] vdd 
+ read_mux 
* No parameters

xmux_124 
+ sel_b[0] bl[124] br[124] bl_out[31] br_out[31] vdd 
+ read_mux 
* No parameters

xmux_125 
+ sel_b[1] bl[125] br[125] bl_out[31] br_out[31] vdd 
+ read_mux 
* No parameters

xmux_126 
+ sel_b[2] bl[126] br[126] bl_out[31] br_out[31] vdd 
+ read_mux 
* No parameters

xmux_127 
+ sel_b[3] bl[127] br[127] bl_out[31] br_out[31] vdd 
+ read_mux 
* No parameters

.ENDS

.SUBCKT write_mux 
+ we data data_b bl br vss 

xMMUXBR 
+ br data x vss 
+ sky130_fd_pr__nfet_01v8 
+ w='2.0' l='0.15' 

xMMUXBL 
+ bl data_b x vss 
+ sky130_fd_pr__nfet_01v8 
+ w='2.0' l='0.15' 

xMPD 
+ x we vss vss 
+ sky130_fd_pr__nfet_01v8 
+ w='2.0' l='0.15' 

.ENDS

.SUBCKT write_mux_array 
+ we[3] we[2] we[1] we[0] data[31] data[30] data[29] data[28] data[27] data[26] data[25] data[24] data[23] data[22] data[21] data[20] data[19] data[18] data[17] data[16] data[15] data[14] data[13] data[12] data[11] data[10] data[9] data[8] data[7] data[6] data[5] data[4] data[3] data[2] data[1] data[0] data_b[31] data_b[30] data_b[29] data_b[28] data_b[27] data_b[26] data_b[25] data_b[24] data_b[23] data_b[22] data_b[21] data_b[20] data_b[19] data_b[18] data_b[17] data_b[16] data_b[15] data_b[14] data_b[13] data_b[12] data_b[11] data_b[10] data_b[9] data_b[8] data_b[7] data_b[6] data_b[5] data_b[4] data_b[3] data_b[2] data_b[1] data_b[0] bl[127] bl[126] bl[125] bl[124] bl[123] bl[122] bl[121] bl[120] bl[119] bl[118] bl[117] bl[116] bl[115] bl[114] bl[113] bl[112] bl[111] bl[110] bl[109] bl[108] bl[107] bl[106] bl[105] bl[104] bl[103] bl[102] bl[101] bl[100] bl[99] bl[98] bl[97] bl[96] bl[95] bl[94] bl[93] bl[92] bl[91] bl[90] bl[89] bl[88] bl[87] bl[86] bl[85] bl[84] bl[83] bl[82] bl[81] bl[80] bl[79] bl[78] bl[77] bl[76] bl[75] bl[74] bl[73] bl[72] bl[71] bl[70] bl[69] bl[68] bl[67] bl[66] bl[65] bl[64] bl[63] bl[62] bl[61] bl[60] bl[59] bl[58] bl[57] bl[56] bl[55] bl[54] bl[53] bl[52] bl[51] bl[50] bl[49] bl[48] bl[47] bl[46] bl[45] bl[44] bl[43] bl[42] bl[41] bl[40] bl[39] bl[38] bl[37] bl[36] bl[35] bl[34] bl[33] bl[32] bl[31] bl[30] bl[29] bl[28] bl[27] bl[26] bl[25] bl[24] bl[23] bl[22] bl[21] bl[20] bl[19] bl[18] bl[17] bl[16] bl[15] bl[14] bl[13] bl[12] bl[11] bl[10] bl[9] bl[8] bl[7] bl[6] bl[5] bl[4] bl[3] bl[2] bl[1] bl[0] br[127] br[126] br[125] br[124] br[123] br[122] br[121] br[120] br[119] br[118] br[117] br[116] br[115] br[114] br[113] br[112] br[111] br[110] br[109] br[108] br[107] br[106] br[105] br[104] br[103] br[102] br[101] br[100] br[99] br[98] br[97] br[96] br[95] br[94] br[93] br[92] br[91] br[90] br[89] br[88] br[87] br[86] br[85] br[84] br[83] br[82] br[81] br[80] br[79] br[78] br[77] br[76] br[75] br[74] br[73] br[72] br[71] br[70] br[69] br[68] br[67] br[66] br[65] br[64] br[63] br[62] br[61] br[60] br[59] br[58] br[57] br[56] br[55] br[54] br[53] br[52] br[51] br[50] br[49] br[48] br[47] br[46] br[45] br[44] br[43] br[42] br[41] br[40] br[39] br[38] br[37] br[36] br[35] br[34] br[33] br[32] br[31] br[30] br[29] br[28] br[27] br[26] br[25] br[24] br[23] br[22] br[21] br[20] br[19] br[18] br[17] br[16] br[15] br[14] br[13] br[12] br[11] br[10] br[9] br[8] br[7] br[6] br[5] br[4] br[3] br[2] br[1] br[0] vss 

xmux_0 
+ we[0] data[0] data_b[0] bl[0] br[0] vss 
+ write_mux 
* No parameters

xmux_1 
+ we[1] data[0] data_b[0] bl[1] br[1] vss 
+ write_mux 
* No parameters

xmux_2 
+ we[2] data[0] data_b[0] bl[2] br[2] vss 
+ write_mux 
* No parameters

xmux_3 
+ we[3] data[0] data_b[0] bl[3] br[3] vss 
+ write_mux 
* No parameters

xmux_4 
+ we[0] data[1] data_b[1] bl[4] br[4] vss 
+ write_mux 
* No parameters

xmux_5 
+ we[1] data[1] data_b[1] bl[5] br[5] vss 
+ write_mux 
* No parameters

xmux_6 
+ we[2] data[1] data_b[1] bl[6] br[6] vss 
+ write_mux 
* No parameters

xmux_7 
+ we[3] data[1] data_b[1] bl[7] br[7] vss 
+ write_mux 
* No parameters

xmux_8 
+ we[0] data[2] data_b[2] bl[8] br[8] vss 
+ write_mux 
* No parameters

xmux_9 
+ we[1] data[2] data_b[2] bl[9] br[9] vss 
+ write_mux 
* No parameters

xmux_10 
+ we[2] data[2] data_b[2] bl[10] br[10] vss 
+ write_mux 
* No parameters

xmux_11 
+ we[3] data[2] data_b[2] bl[11] br[11] vss 
+ write_mux 
* No parameters

xmux_12 
+ we[0] data[3] data_b[3] bl[12] br[12] vss 
+ write_mux 
* No parameters

xmux_13 
+ we[1] data[3] data_b[3] bl[13] br[13] vss 
+ write_mux 
* No parameters

xmux_14 
+ we[2] data[3] data_b[3] bl[14] br[14] vss 
+ write_mux 
* No parameters

xmux_15 
+ we[3] data[3] data_b[3] bl[15] br[15] vss 
+ write_mux 
* No parameters

xmux_16 
+ we[0] data[4] data_b[4] bl[16] br[16] vss 
+ write_mux 
* No parameters

xmux_17 
+ we[1] data[4] data_b[4] bl[17] br[17] vss 
+ write_mux 
* No parameters

xmux_18 
+ we[2] data[4] data_b[4] bl[18] br[18] vss 
+ write_mux 
* No parameters

xmux_19 
+ we[3] data[4] data_b[4] bl[19] br[19] vss 
+ write_mux 
* No parameters

xmux_20 
+ we[0] data[5] data_b[5] bl[20] br[20] vss 
+ write_mux 
* No parameters

xmux_21 
+ we[1] data[5] data_b[5] bl[21] br[21] vss 
+ write_mux 
* No parameters

xmux_22 
+ we[2] data[5] data_b[5] bl[22] br[22] vss 
+ write_mux 
* No parameters

xmux_23 
+ we[3] data[5] data_b[5] bl[23] br[23] vss 
+ write_mux 
* No parameters

xmux_24 
+ we[0] data[6] data_b[6] bl[24] br[24] vss 
+ write_mux 
* No parameters

xmux_25 
+ we[1] data[6] data_b[6] bl[25] br[25] vss 
+ write_mux 
* No parameters

xmux_26 
+ we[2] data[6] data_b[6] bl[26] br[26] vss 
+ write_mux 
* No parameters

xmux_27 
+ we[3] data[6] data_b[6] bl[27] br[27] vss 
+ write_mux 
* No parameters

xmux_28 
+ we[0] data[7] data_b[7] bl[28] br[28] vss 
+ write_mux 
* No parameters

xmux_29 
+ we[1] data[7] data_b[7] bl[29] br[29] vss 
+ write_mux 
* No parameters

xmux_30 
+ we[2] data[7] data_b[7] bl[30] br[30] vss 
+ write_mux 
* No parameters

xmux_31 
+ we[3] data[7] data_b[7] bl[31] br[31] vss 
+ write_mux 
* No parameters

xmux_32 
+ we[0] data[8] data_b[8] bl[32] br[32] vss 
+ write_mux 
* No parameters

xmux_33 
+ we[1] data[8] data_b[8] bl[33] br[33] vss 
+ write_mux 
* No parameters

xmux_34 
+ we[2] data[8] data_b[8] bl[34] br[34] vss 
+ write_mux 
* No parameters

xmux_35 
+ we[3] data[8] data_b[8] bl[35] br[35] vss 
+ write_mux 
* No parameters

xmux_36 
+ we[0] data[9] data_b[9] bl[36] br[36] vss 
+ write_mux 
* No parameters

xmux_37 
+ we[1] data[9] data_b[9] bl[37] br[37] vss 
+ write_mux 
* No parameters

xmux_38 
+ we[2] data[9] data_b[9] bl[38] br[38] vss 
+ write_mux 
* No parameters

xmux_39 
+ we[3] data[9] data_b[9] bl[39] br[39] vss 
+ write_mux 
* No parameters

xmux_40 
+ we[0] data[10] data_b[10] bl[40] br[40] vss 
+ write_mux 
* No parameters

xmux_41 
+ we[1] data[10] data_b[10] bl[41] br[41] vss 
+ write_mux 
* No parameters

xmux_42 
+ we[2] data[10] data_b[10] bl[42] br[42] vss 
+ write_mux 
* No parameters

xmux_43 
+ we[3] data[10] data_b[10] bl[43] br[43] vss 
+ write_mux 
* No parameters

xmux_44 
+ we[0] data[11] data_b[11] bl[44] br[44] vss 
+ write_mux 
* No parameters

xmux_45 
+ we[1] data[11] data_b[11] bl[45] br[45] vss 
+ write_mux 
* No parameters

xmux_46 
+ we[2] data[11] data_b[11] bl[46] br[46] vss 
+ write_mux 
* No parameters

xmux_47 
+ we[3] data[11] data_b[11] bl[47] br[47] vss 
+ write_mux 
* No parameters

xmux_48 
+ we[0] data[12] data_b[12] bl[48] br[48] vss 
+ write_mux 
* No parameters

xmux_49 
+ we[1] data[12] data_b[12] bl[49] br[49] vss 
+ write_mux 
* No parameters

xmux_50 
+ we[2] data[12] data_b[12] bl[50] br[50] vss 
+ write_mux 
* No parameters

xmux_51 
+ we[3] data[12] data_b[12] bl[51] br[51] vss 
+ write_mux 
* No parameters

xmux_52 
+ we[0] data[13] data_b[13] bl[52] br[52] vss 
+ write_mux 
* No parameters

xmux_53 
+ we[1] data[13] data_b[13] bl[53] br[53] vss 
+ write_mux 
* No parameters

xmux_54 
+ we[2] data[13] data_b[13] bl[54] br[54] vss 
+ write_mux 
* No parameters

xmux_55 
+ we[3] data[13] data_b[13] bl[55] br[55] vss 
+ write_mux 
* No parameters

xmux_56 
+ we[0] data[14] data_b[14] bl[56] br[56] vss 
+ write_mux 
* No parameters

xmux_57 
+ we[1] data[14] data_b[14] bl[57] br[57] vss 
+ write_mux 
* No parameters

xmux_58 
+ we[2] data[14] data_b[14] bl[58] br[58] vss 
+ write_mux 
* No parameters

xmux_59 
+ we[3] data[14] data_b[14] bl[59] br[59] vss 
+ write_mux 
* No parameters

xmux_60 
+ we[0] data[15] data_b[15] bl[60] br[60] vss 
+ write_mux 
* No parameters

xmux_61 
+ we[1] data[15] data_b[15] bl[61] br[61] vss 
+ write_mux 
* No parameters

xmux_62 
+ we[2] data[15] data_b[15] bl[62] br[62] vss 
+ write_mux 
* No parameters

xmux_63 
+ we[3] data[15] data_b[15] bl[63] br[63] vss 
+ write_mux 
* No parameters

xmux_64 
+ we[0] data[16] data_b[16] bl[64] br[64] vss 
+ write_mux 
* No parameters

xmux_65 
+ we[1] data[16] data_b[16] bl[65] br[65] vss 
+ write_mux 
* No parameters

xmux_66 
+ we[2] data[16] data_b[16] bl[66] br[66] vss 
+ write_mux 
* No parameters

xmux_67 
+ we[3] data[16] data_b[16] bl[67] br[67] vss 
+ write_mux 
* No parameters

xmux_68 
+ we[0] data[17] data_b[17] bl[68] br[68] vss 
+ write_mux 
* No parameters

xmux_69 
+ we[1] data[17] data_b[17] bl[69] br[69] vss 
+ write_mux 
* No parameters

xmux_70 
+ we[2] data[17] data_b[17] bl[70] br[70] vss 
+ write_mux 
* No parameters

xmux_71 
+ we[3] data[17] data_b[17] bl[71] br[71] vss 
+ write_mux 
* No parameters

xmux_72 
+ we[0] data[18] data_b[18] bl[72] br[72] vss 
+ write_mux 
* No parameters

xmux_73 
+ we[1] data[18] data_b[18] bl[73] br[73] vss 
+ write_mux 
* No parameters

xmux_74 
+ we[2] data[18] data_b[18] bl[74] br[74] vss 
+ write_mux 
* No parameters

xmux_75 
+ we[3] data[18] data_b[18] bl[75] br[75] vss 
+ write_mux 
* No parameters

xmux_76 
+ we[0] data[19] data_b[19] bl[76] br[76] vss 
+ write_mux 
* No parameters

xmux_77 
+ we[1] data[19] data_b[19] bl[77] br[77] vss 
+ write_mux 
* No parameters

xmux_78 
+ we[2] data[19] data_b[19] bl[78] br[78] vss 
+ write_mux 
* No parameters

xmux_79 
+ we[3] data[19] data_b[19] bl[79] br[79] vss 
+ write_mux 
* No parameters

xmux_80 
+ we[0] data[20] data_b[20] bl[80] br[80] vss 
+ write_mux 
* No parameters

xmux_81 
+ we[1] data[20] data_b[20] bl[81] br[81] vss 
+ write_mux 
* No parameters

xmux_82 
+ we[2] data[20] data_b[20] bl[82] br[82] vss 
+ write_mux 
* No parameters

xmux_83 
+ we[3] data[20] data_b[20] bl[83] br[83] vss 
+ write_mux 
* No parameters

xmux_84 
+ we[0] data[21] data_b[21] bl[84] br[84] vss 
+ write_mux 
* No parameters

xmux_85 
+ we[1] data[21] data_b[21] bl[85] br[85] vss 
+ write_mux 
* No parameters

xmux_86 
+ we[2] data[21] data_b[21] bl[86] br[86] vss 
+ write_mux 
* No parameters

xmux_87 
+ we[3] data[21] data_b[21] bl[87] br[87] vss 
+ write_mux 
* No parameters

xmux_88 
+ we[0] data[22] data_b[22] bl[88] br[88] vss 
+ write_mux 
* No parameters

xmux_89 
+ we[1] data[22] data_b[22] bl[89] br[89] vss 
+ write_mux 
* No parameters

xmux_90 
+ we[2] data[22] data_b[22] bl[90] br[90] vss 
+ write_mux 
* No parameters

xmux_91 
+ we[3] data[22] data_b[22] bl[91] br[91] vss 
+ write_mux 
* No parameters

xmux_92 
+ we[0] data[23] data_b[23] bl[92] br[92] vss 
+ write_mux 
* No parameters

xmux_93 
+ we[1] data[23] data_b[23] bl[93] br[93] vss 
+ write_mux 
* No parameters

xmux_94 
+ we[2] data[23] data_b[23] bl[94] br[94] vss 
+ write_mux 
* No parameters

xmux_95 
+ we[3] data[23] data_b[23] bl[95] br[95] vss 
+ write_mux 
* No parameters

xmux_96 
+ we[0] data[24] data_b[24] bl[96] br[96] vss 
+ write_mux 
* No parameters

xmux_97 
+ we[1] data[24] data_b[24] bl[97] br[97] vss 
+ write_mux 
* No parameters

xmux_98 
+ we[2] data[24] data_b[24] bl[98] br[98] vss 
+ write_mux 
* No parameters

xmux_99 
+ we[3] data[24] data_b[24] bl[99] br[99] vss 
+ write_mux 
* No parameters

xmux_100 
+ we[0] data[25] data_b[25] bl[100] br[100] vss 
+ write_mux 
* No parameters

xmux_101 
+ we[1] data[25] data_b[25] bl[101] br[101] vss 
+ write_mux 
* No parameters

xmux_102 
+ we[2] data[25] data_b[25] bl[102] br[102] vss 
+ write_mux 
* No parameters

xmux_103 
+ we[3] data[25] data_b[25] bl[103] br[103] vss 
+ write_mux 
* No parameters

xmux_104 
+ we[0] data[26] data_b[26] bl[104] br[104] vss 
+ write_mux 
* No parameters

xmux_105 
+ we[1] data[26] data_b[26] bl[105] br[105] vss 
+ write_mux 
* No parameters

xmux_106 
+ we[2] data[26] data_b[26] bl[106] br[106] vss 
+ write_mux 
* No parameters

xmux_107 
+ we[3] data[26] data_b[26] bl[107] br[107] vss 
+ write_mux 
* No parameters

xmux_108 
+ we[0] data[27] data_b[27] bl[108] br[108] vss 
+ write_mux 
* No parameters

xmux_109 
+ we[1] data[27] data_b[27] bl[109] br[109] vss 
+ write_mux 
* No parameters

xmux_110 
+ we[2] data[27] data_b[27] bl[110] br[110] vss 
+ write_mux 
* No parameters

xmux_111 
+ we[3] data[27] data_b[27] bl[111] br[111] vss 
+ write_mux 
* No parameters

xmux_112 
+ we[0] data[28] data_b[28] bl[112] br[112] vss 
+ write_mux 
* No parameters

xmux_113 
+ we[1] data[28] data_b[28] bl[113] br[113] vss 
+ write_mux 
* No parameters

xmux_114 
+ we[2] data[28] data_b[28] bl[114] br[114] vss 
+ write_mux 
* No parameters

xmux_115 
+ we[3] data[28] data_b[28] bl[115] br[115] vss 
+ write_mux 
* No parameters

xmux_116 
+ we[0] data[29] data_b[29] bl[116] br[116] vss 
+ write_mux 
* No parameters

xmux_117 
+ we[1] data[29] data_b[29] bl[117] br[117] vss 
+ write_mux 
* No parameters

xmux_118 
+ we[2] data[29] data_b[29] bl[118] br[118] vss 
+ write_mux 
* No parameters

xmux_119 
+ we[3] data[29] data_b[29] bl[119] br[119] vss 
+ write_mux 
* No parameters

xmux_120 
+ we[0] data[30] data_b[30] bl[120] br[120] vss 
+ write_mux 
* No parameters

xmux_121 
+ we[1] data[30] data_b[30] bl[121] br[121] vss 
+ write_mux 
* No parameters

xmux_122 
+ we[2] data[30] data_b[30] bl[122] br[122] vss 
+ write_mux 
* No parameters

xmux_123 
+ we[3] data[30] data_b[30] bl[123] br[123] vss 
+ write_mux 
* No parameters

xmux_124 
+ we[0] data[31] data_b[31] bl[124] br[124] vss 
+ write_mux 
* No parameters

xmux_125 
+ we[1] data[31] data_b[31] bl[125] br[125] vss 
+ write_mux 
* No parameters

xmux_126 
+ we[2] data[31] data_b[31] bl[126] br[126] vss 
+ write_mux 
* No parameters

xmux_127 
+ we[3] data[31] data_b[31] bl[127] br[127] vss 
+ write_mux 
* No parameters

.ENDS

.SUBCKT data_dff_array 
+ vdd vss clk d[31] d[30] d[29] d[28] d[27] d[26] d[25] d[24] d[23] d[22] d[21] d[20] d[19] d[18] d[17] d[16] d[15] d[14] d[13] d[12] d[11] d[10] d[9] d[8] d[7] d[6] d[5] d[4] d[3] d[2] d[1] d[0] q[31] q[30] q[29] q[28] q[27] q[26] q[25] q[24] q[23] q[22] q[21] q[20] q[19] q[18] q[17] q[16] q[15] q[14] q[13] q[12] q[11] q[10] q[9] q[8] q[7] q[6] q[5] q[4] q[3] q[2] q[1] q[0] q_b[31] q_b[30] q_b[29] q_b[28] q_b[27] q_b[26] q_b[25] q_b[24] q_b[23] q_b[22] q_b[21] q_b[20] q_b[19] q_b[18] q_b[17] q_b[16] q_b[15] q_b[14] q_b[13] q_b[12] q_b[11] q_b[10] q_b[9] q_b[8] q_b[7] q_b[6] q_b[5] q_b[4] q_b[3] q_b[2] q_b[1] q_b[0] 

xdff_0 
+ vdd vss clk d[0] q[0] q_b[0] 
+ openram_dff 
* No parameters

xdff_1 
+ vdd vss clk d[1] q[1] q_b[1] 
+ openram_dff 
* No parameters

xdff_2 
+ vdd vss clk d[2] q[2] q_b[2] 
+ openram_dff 
* No parameters

xdff_3 
+ vdd vss clk d[3] q[3] q_b[3] 
+ openram_dff 
* No parameters

xdff_4 
+ vdd vss clk d[4] q[4] q_b[4] 
+ openram_dff 
* No parameters

xdff_5 
+ vdd vss clk d[5] q[5] q_b[5] 
+ openram_dff 
* No parameters

xdff_6 
+ vdd vss clk d[6] q[6] q_b[6] 
+ openram_dff 
* No parameters

xdff_7 
+ vdd vss clk d[7] q[7] q_b[7] 
+ openram_dff 
* No parameters

xdff_8 
+ vdd vss clk d[8] q[8] q_b[8] 
+ openram_dff 
* No parameters

xdff_9 
+ vdd vss clk d[9] q[9] q_b[9] 
+ openram_dff 
* No parameters

xdff_10 
+ vdd vss clk d[10] q[10] q_b[10] 
+ openram_dff 
* No parameters

xdff_11 
+ vdd vss clk d[11] q[11] q_b[11] 
+ openram_dff 
* No parameters

xdff_12 
+ vdd vss clk d[12] q[12] q_b[12] 
+ openram_dff 
* No parameters

xdff_13 
+ vdd vss clk d[13] q[13] q_b[13] 
+ openram_dff 
* No parameters

xdff_14 
+ vdd vss clk d[14] q[14] q_b[14] 
+ openram_dff 
* No parameters

xdff_15 
+ vdd vss clk d[15] q[15] q_b[15] 
+ openram_dff 
* No parameters

xdff_16 
+ vdd vss clk d[16] q[16] q_b[16] 
+ openram_dff 
* No parameters

xdff_17 
+ vdd vss clk d[17] q[17] q_b[17] 
+ openram_dff 
* No parameters

xdff_18 
+ vdd vss clk d[18] q[18] q_b[18] 
+ openram_dff 
* No parameters

xdff_19 
+ vdd vss clk d[19] q[19] q_b[19] 
+ openram_dff 
* No parameters

xdff_20 
+ vdd vss clk d[20] q[20] q_b[20] 
+ openram_dff 
* No parameters

xdff_21 
+ vdd vss clk d[21] q[21] q_b[21] 
+ openram_dff 
* No parameters

xdff_22 
+ vdd vss clk d[22] q[22] q_b[22] 
+ openram_dff 
* No parameters

xdff_23 
+ vdd vss clk d[23] q[23] q_b[23] 
+ openram_dff 
* No parameters

xdff_24 
+ vdd vss clk d[24] q[24] q_b[24] 
+ openram_dff 
* No parameters

xdff_25 
+ vdd vss clk d[25] q[25] q_b[25] 
+ openram_dff 
* No parameters

xdff_26 
+ vdd vss clk d[26] q[26] q_b[26] 
+ openram_dff 
* No parameters

xdff_27 
+ vdd vss clk d[27] q[27] q_b[27] 
+ openram_dff 
* No parameters

xdff_28 
+ vdd vss clk d[28] q[28] q_b[28] 
+ openram_dff 
* No parameters

xdff_29 
+ vdd vss clk d[29] q[29] q_b[29] 
+ openram_dff 
* No parameters

xdff_30 
+ vdd vss clk d[30] q[30] q_b[30] 
+ openram_dff 
* No parameters

xdff_31 
+ vdd vss clk d[31] q[31] q_b[31] 
+ openram_dff 
* No parameters

.ENDS

.SUBCKT addr_dff_array 
+ vdd vss clk d[5] d[4] d[3] d[2] d[1] d[0] q[5] q[4] q[3] q[2] q[1] q[0] q_b[5] q_b[4] q_b[3] q_b[2] q_b[1] q_b[0] 

xdff_0 
+ vdd vss clk d[0] q[0] q_b[0] 
+ openram_dff 
* No parameters

xdff_1 
+ vdd vss clk d[1] q[1] q_b[1] 
+ openram_dff 
* No parameters

xdff_2 
+ vdd vss clk d[2] q[2] q_b[2] 
+ openram_dff 
* No parameters

xdff_3 
+ vdd vss clk d[3] q[3] q_b[3] 
+ openram_dff 
* No parameters

xdff_4 
+ vdd vss clk d[4] q[4] q_b[4] 
+ openram_dff 
* No parameters

xdff_5 
+ vdd vss clk d[5] q[5] q_b[5] 
+ openram_dff 
* No parameters

.ENDS

.SUBCKT col_data_inv 
+ din din_b vdd vss 

xMP0 
+ din_b din vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.6' l='0.15' 

xMN0 
+ din_b din vss vss 
+ sky130_fd_pr__nfet_01v8 
+ w='1.4' l='0.15' 

.ENDS

.SUBCKT col_inv_array 
+ din[31] din[30] din[29] din[28] din[27] din[26] din[25] din[24] din[23] din[22] din[21] din[20] din[19] din[18] din[17] din[16] din[15] din[14] din[13] din[12] din[11] din[10] din[9] din[8] din[7] din[6] din[5] din[4] din[3] din[2] din[1] din[0] din_b[31] din_b[30] din_b[29] din_b[28] din_b[27] din_b[26] din_b[25] din_b[24] din_b[23] din_b[22] din_b[21] din_b[20] din_b[19] din_b[18] din_b[17] din_b[16] din_b[15] din_b[14] din_b[13] din_b[12] din_b[11] din_b[10] din_b[9] din_b[8] din_b[7] din_b[6] din_b[5] din_b[4] din_b[3] din_b[2] din_b[1] din_b[0] vdd vss 

xinv_0 
+ din[0] din_b[0] vdd vss 
+ col_data_inv 
* No parameters

xinv_1 
+ din[1] din_b[1] vdd vss 
+ col_data_inv 
* No parameters

xinv_2 
+ din[2] din_b[2] vdd vss 
+ col_data_inv 
* No parameters

xinv_3 
+ din[3] din_b[3] vdd vss 
+ col_data_inv 
* No parameters

xinv_4 
+ din[4] din_b[4] vdd vss 
+ col_data_inv 
* No parameters

xinv_5 
+ din[5] din_b[5] vdd vss 
+ col_data_inv 
* No parameters

xinv_6 
+ din[6] din_b[6] vdd vss 
+ col_data_inv 
* No parameters

xinv_7 
+ din[7] din_b[7] vdd vss 
+ col_data_inv 
* No parameters

xinv_8 
+ din[8] din_b[8] vdd vss 
+ col_data_inv 
* No parameters

xinv_9 
+ din[9] din_b[9] vdd vss 
+ col_data_inv 
* No parameters

xinv_10 
+ din[10] din_b[10] vdd vss 
+ col_data_inv 
* No parameters

xinv_11 
+ din[11] din_b[11] vdd vss 
+ col_data_inv 
* No parameters

xinv_12 
+ din[12] din_b[12] vdd vss 
+ col_data_inv 
* No parameters

xinv_13 
+ din[13] din_b[13] vdd vss 
+ col_data_inv 
* No parameters

xinv_14 
+ din[14] din_b[14] vdd vss 
+ col_data_inv 
* No parameters

xinv_15 
+ din[15] din_b[15] vdd vss 
+ col_data_inv 
* No parameters

xinv_16 
+ din[16] din_b[16] vdd vss 
+ col_data_inv 
* No parameters

xinv_17 
+ din[17] din_b[17] vdd vss 
+ col_data_inv 
* No parameters

xinv_18 
+ din[18] din_b[18] vdd vss 
+ col_data_inv 
* No parameters

xinv_19 
+ din[19] din_b[19] vdd vss 
+ col_data_inv 
* No parameters

xinv_20 
+ din[20] din_b[20] vdd vss 
+ col_data_inv 
* No parameters

xinv_21 
+ din[21] din_b[21] vdd vss 
+ col_data_inv 
* No parameters

xinv_22 
+ din[22] din_b[22] vdd vss 
+ col_data_inv 
* No parameters

xinv_23 
+ din[23] din_b[23] vdd vss 
+ col_data_inv 
* No parameters

xinv_24 
+ din[24] din_b[24] vdd vss 
+ col_data_inv 
* No parameters

xinv_25 
+ din[25] din_b[25] vdd vss 
+ col_data_inv 
* No parameters

xinv_26 
+ din[26] din_b[26] vdd vss 
+ col_data_inv 
* No parameters

xinv_27 
+ din[27] din_b[27] vdd vss 
+ col_data_inv 
* No parameters

xinv_28 
+ din[28] din_b[28] vdd vss 
+ col_data_inv 
* No parameters

xinv_29 
+ din[29] din_b[29] vdd vss 
+ col_data_inv 
* No parameters

xinv_30 
+ din[30] din_b[30] vdd vss 
+ col_data_inv 
* No parameters

xinv_31 
+ din[31] din_b[31] vdd vss 
+ col_data_inv 
* No parameters

.ENDS

.SUBCKT sense_amp_array 
+ vdd vss clk bl[31] bl[30] bl[29] bl[28] bl[27] bl[26] bl[25] bl[24] bl[23] bl[22] bl[21] bl[20] bl[19] bl[18] bl[17] bl[16] bl[15] bl[14] bl[13] bl[12] bl[11] bl[10] bl[9] bl[8] bl[7] bl[6] bl[5] bl[4] bl[3] bl[2] bl[1] bl[0] br[31] br[30] br[29] br[28] br[27] br[26] br[25] br[24] br[23] br[22] br[21] br[20] br[19] br[18] br[17] br[16] br[15] br[14] br[13] br[12] br[11] br[10] br[9] br[8] br[7] br[6] br[5] br[4] br[3] br[2] br[1] br[0] data[31] data[30] data[29] data[28] data[27] data[26] data[25] data[24] data[23] data[22] data[21] data[20] data[19] data[18] data[17] data[16] data[15] data[14] data[13] data[12] data[11] data[10] data[9] data[8] data[7] data[6] data[5] data[4] data[3] data[2] data[1] data[0] data_b[31] data_b[30] data_b[29] data_b[28] data_b[27] data_b[26] data_b[25] data_b[24] data_b[23] data_b[22] data_b[21] data_b[20] data_b[19] data_b[18] data_b[17] data_b[16] data_b[15] data_b[14] data_b[13] data_b[12] data_b[11] data_b[10] data_b[9] data_b[8] data_b[7] data_b[6] data_b[5] data_b[4] data_b[3] data_b[2] data_b[1] data_b[0] 

xsense_amp_0 
+ clk br[0] bl[0] data_b[0] data[0] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_1 
+ clk br[1] bl[1] data_b[1] data[1] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_2 
+ clk br[2] bl[2] data_b[2] data[2] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_3 
+ clk br[3] bl[3] data_b[3] data[3] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_4 
+ clk br[4] bl[4] data_b[4] data[4] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_5 
+ clk br[5] bl[5] data_b[5] data[5] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_6 
+ clk br[6] bl[6] data_b[6] data[6] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_7 
+ clk br[7] bl[7] data_b[7] data[7] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_8 
+ clk br[8] bl[8] data_b[8] data[8] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_9 
+ clk br[9] bl[9] data_b[9] data[9] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_10 
+ clk br[10] bl[10] data_b[10] data[10] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_11 
+ clk br[11] bl[11] data_b[11] data[11] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_12 
+ clk br[12] bl[12] data_b[12] data[12] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_13 
+ clk br[13] bl[13] data_b[13] data[13] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_14 
+ clk br[14] bl[14] data_b[14] data[14] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_15 
+ clk br[15] bl[15] data_b[15] data[15] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_16 
+ clk br[16] bl[16] data_b[16] data[16] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_17 
+ clk br[17] bl[17] data_b[17] data[17] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_18 
+ clk br[18] bl[18] data_b[18] data[18] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_19 
+ clk br[19] bl[19] data_b[19] data[19] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_20 
+ clk br[20] bl[20] data_b[20] data[20] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_21 
+ clk br[21] bl[21] data_b[21] data[21] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_22 
+ clk br[22] bl[22] data_b[22] data[22] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_23 
+ clk br[23] bl[23] data_b[23] data[23] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_24 
+ clk br[24] bl[24] data_b[24] data[24] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_25 
+ clk br[25] bl[25] data_b[25] data[25] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_26 
+ clk br[26] bl[26] data_b[26] data[26] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_27 
+ clk br[27] bl[27] data_b[27] data[27] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_28 
+ clk br[28] bl[28] data_b[28] data[28] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_29 
+ clk br[29] bl[29] data_b[29] data[29] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_30 
+ clk br[30] bl[30] data_b[30] data[30] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_31 
+ clk br[31] bl[31] data_b[31] data[31] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

.ENDS

.SUBCKT dout_buf 
+ din1 din2 dout1 dout2 vdd vss 

xMP11 
+ x1 din1 vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='1.6' l='0.15' 

xMN11 
+ x1 din1 vss vss 
+ sky130_fd_pr__nfet_01v8 
+ w='1.0' l='0.15' 

xMP21 
+ dout1 x1 vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='3.2' l='0.15' 

xMN21 
+ dout1 x1 vss vss 
+ sky130_fd_pr__nfet_01v8 
+ w='2.0' l='0.15' 

xMP12 
+ x2 din2 vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='1.6' l='0.15' 

xMN12 
+ x2 din2 vss vss 
+ sky130_fd_pr__nfet_01v8 
+ w='1.0' l='0.15' 

xMP22 
+ dout2 x2 vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='3.2' l='0.15' 

xMN22 
+ dout2 x2 vss vss 
+ sky130_fd_pr__nfet_01v8 
+ w='2.0' l='0.15' 

.ENDS

.SUBCKT dout_buf_array 
+ din1[31] din1[30] din1[29] din1[28] din1[27] din1[26] din1[25] din1[24] din1[23] din1[22] din1[21] din1[20] din1[19] din1[18] din1[17] din1[16] din1[15] din1[14] din1[13] din1[12] din1[11] din1[10] din1[9] din1[8] din1[7] din1[6] din1[5] din1[4] din1[3] din1[2] din1[1] din1[0] din2[31] din2[30] din2[29] din2[28] din2[27] din2[26] din2[25] din2[24] din2[23] din2[22] din2[21] din2[20] din2[19] din2[18] din2[17] din2[16] din2[15] din2[14] din2[13] din2[12] din2[11] din2[10] din2[9] din2[8] din2[7] din2[6] din2[5] din2[4] din2[3] din2[2] din2[1] din2[0] dout1[31] dout1[30] dout1[29] dout1[28] dout1[27] dout1[26] dout1[25] dout1[24] dout1[23] dout1[22] dout1[21] dout1[20] dout1[19] dout1[18] dout1[17] dout1[16] dout1[15] dout1[14] dout1[13] dout1[12] dout1[11] dout1[10] dout1[9] dout1[8] dout1[7] dout1[6] dout1[5] dout1[4] dout1[3] dout1[2] dout1[1] dout1[0] dout2[31] dout2[30] dout2[29] dout2[28] dout2[27] dout2[26] dout2[25] dout2[24] dout2[23] dout2[22] dout2[21] dout2[20] dout2[19] dout2[18] dout2[17] dout2[16] dout2[15] dout2[14] dout2[13] dout2[12] dout2[11] dout2[10] dout2[9] dout2[8] dout2[7] dout2[6] dout2[5] dout2[4] dout2[3] dout2[2] dout2[1] dout2[0] vdd vss 

xbuf_0 
+ din1[0] din2[0] dout1[0] dout2[0] vdd vss 
+ dout_buf 
* No parameters

xbuf_1 
+ din1[1] din2[1] dout1[1] dout2[1] vdd vss 
+ dout_buf 
* No parameters

xbuf_2 
+ din1[2] din2[2] dout1[2] dout2[2] vdd vss 
+ dout_buf 
* No parameters

xbuf_3 
+ din1[3] din2[3] dout1[3] dout2[3] vdd vss 
+ dout_buf 
* No parameters

xbuf_4 
+ din1[4] din2[4] dout1[4] dout2[4] vdd vss 
+ dout_buf 
* No parameters

xbuf_5 
+ din1[5] din2[5] dout1[5] dout2[5] vdd vss 
+ dout_buf 
* No parameters

xbuf_6 
+ din1[6] din2[6] dout1[6] dout2[6] vdd vss 
+ dout_buf 
* No parameters

xbuf_7 
+ din1[7] din2[7] dout1[7] dout2[7] vdd vss 
+ dout_buf 
* No parameters

xbuf_8 
+ din1[8] din2[8] dout1[8] dout2[8] vdd vss 
+ dout_buf 
* No parameters

xbuf_9 
+ din1[9] din2[9] dout1[9] dout2[9] vdd vss 
+ dout_buf 
* No parameters

xbuf_10 
+ din1[10] din2[10] dout1[10] dout2[10] vdd vss 
+ dout_buf 
* No parameters

xbuf_11 
+ din1[11] din2[11] dout1[11] dout2[11] vdd vss 
+ dout_buf 
* No parameters

xbuf_12 
+ din1[12] din2[12] dout1[12] dout2[12] vdd vss 
+ dout_buf 
* No parameters

xbuf_13 
+ din1[13] din2[13] dout1[13] dout2[13] vdd vss 
+ dout_buf 
* No parameters

xbuf_14 
+ din1[14] din2[14] dout1[14] dout2[14] vdd vss 
+ dout_buf 
* No parameters

xbuf_15 
+ din1[15] din2[15] dout1[15] dout2[15] vdd vss 
+ dout_buf 
* No parameters

xbuf_16 
+ din1[16] din2[16] dout1[16] dout2[16] vdd vss 
+ dout_buf 
* No parameters

xbuf_17 
+ din1[17] din2[17] dout1[17] dout2[17] vdd vss 
+ dout_buf 
* No parameters

xbuf_18 
+ din1[18] din2[18] dout1[18] dout2[18] vdd vss 
+ dout_buf 
* No parameters

xbuf_19 
+ din1[19] din2[19] dout1[19] dout2[19] vdd vss 
+ dout_buf 
* No parameters

xbuf_20 
+ din1[20] din2[20] dout1[20] dout2[20] vdd vss 
+ dout_buf 
* No parameters

xbuf_21 
+ din1[21] din2[21] dout1[21] dout2[21] vdd vss 
+ dout_buf 
* No parameters

xbuf_22 
+ din1[22] din2[22] dout1[22] dout2[22] vdd vss 
+ dout_buf 
* No parameters

xbuf_23 
+ din1[23] din2[23] dout1[23] dout2[23] vdd vss 
+ dout_buf 
* No parameters

xbuf_24 
+ din1[24] din2[24] dout1[24] dout2[24] vdd vss 
+ dout_buf 
* No parameters

xbuf_25 
+ din1[25] din2[25] dout1[25] dout2[25] vdd vss 
+ dout_buf 
* No parameters

xbuf_26 
+ din1[26] din2[26] dout1[26] dout2[26] vdd vss 
+ dout_buf 
* No parameters

xbuf_27 
+ din1[27] din2[27] dout1[27] dout2[27] vdd vss 
+ dout_buf 
* No parameters

xbuf_28 
+ din1[28] din2[28] dout1[28] dout2[28] vdd vss 
+ dout_buf 
* No parameters

xbuf_29 
+ din1[29] din2[29] dout1[29] dout2[29] vdd vss 
+ dout_buf 
* No parameters

xbuf_30 
+ din1[30] din2[30] dout1[30] dout2[30] vdd vss 
+ dout_buf 
* No parameters

xbuf_31 
+ din1[31] din2[31] dout1[31] dout2[31] vdd vss 
+ dout_buf 
* No parameters

.ENDS

.SUBCKT we_control_and2_nand 
+ gnd vdd a b y 

xn1 
+ x a gnd gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='3.0' l='0.15' 

xn2 
+ y b x gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='3.0' l='0.15' 

xp1 
+ y a vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='4.0' l='0.15' 

xp2 
+ y b vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='4.0' l='0.15' 

.ENDS

.SUBCKT we_control_and2_inv 
+ gnd vdd din din_b 

xn 
+ din_b din gnd gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='8.0' l='0.15' 

xp 
+ din_b din vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='12.0' l='0.15' 

.ENDS

.SUBCKT we_control_and2 
+ a b y vdd vss 

xnand 
+ vss vdd a b tmp 
+ we_control_and2_nand 
* No parameters

xinv 
+ vss vdd tmp y 
+ we_control_and2_inv 
* No parameters

.ENDS

.SUBCKT we_control 
+ wr_en sel[3] sel[2] sel[1] sel[0] write_driver_en[3] write_driver_en[2] write_driver_en[1] write_driver_en[0] vdd vss 

xand2_0 
+ sel[0] wr_en write_driver_en[0] vdd vss 
+ we_control_and2 
* No parameters

xand2_1 
+ sel[1] wr_en write_driver_en[1] vdd vss 
+ we_control_and2 
* No parameters

xand2_2 
+ sel[2] wr_en write_driver_en[2] vdd vss 
+ we_control_and2 
* No parameters

xand2_3 
+ sel[3] wr_en write_driver_en[3] vdd vss 
+ we_control_and2 
* No parameters

.ENDS

.SUBCKT control_logic_delay_chain 
+ din dout vdd vss 

xinv_0 
+ din int[0] vdd vss 
+ control_logic_inv 
* No parameters

xinv_1 
+ int[0] int[1] vdd vss 
+ control_logic_inv 
* No parameters

xinv_2 
+ int[1] int[2] vdd vss 
+ control_logic_inv 
* No parameters

xinv_3 
+ int[2] int[3] vdd vss 
+ control_logic_inv 
* No parameters

xinv_4 
+ int[3] int[4] vdd vss 
+ control_logic_inv 
* No parameters

xinv_5 
+ int[4] int[5] vdd vss 
+ control_logic_inv 
* No parameters

xinv_6 
+ int[5] int[6] vdd vss 
+ control_logic_inv 
* No parameters

xinv_7 
+ int[6] int[7] vdd vss 
+ control_logic_inv 
* No parameters

xinv_8 
+ int[7] int[8] vdd vss 
+ control_logic_inv 
* No parameters

xinv_9 
+ int[8] int[9] vdd vss 
+ control_logic_inv 
* No parameters

xinv_10 
+ int[9] int[10] vdd vss 
+ control_logic_inv 
* No parameters

xinv_11 
+ int[10] int[11] vdd vss 
+ control_logic_inv 
* No parameters

xinv_12 
+ int[11] int[12] vdd vss 
+ control_logic_inv 
* No parameters

xinv_13 
+ int[12] int[13] vdd vss 
+ control_logic_inv 
* No parameters

xinv_14 
+ int[13] int[14] vdd vss 
+ control_logic_inv 
* No parameters

xinv_15 
+ int[14] int[15] vdd vss 
+ control_logic_inv 
* No parameters

xinv_16 
+ int[15] int[16] vdd vss 
+ control_logic_inv 
* No parameters

xinv_17 
+ int[16] int[17] vdd vss 
+ control_logic_inv 
* No parameters

xinv_18 
+ int[17] int[18] vdd vss 
+ control_logic_inv 
* No parameters

xinv_19 
+ int[18] int[19] vdd vss 
+ control_logic_inv 
* No parameters

xinv_20 
+ int[19] int[20] vdd vss 
+ control_logic_inv 
* No parameters

xinv_21 
+ int[20] int[21] vdd vss 
+ control_logic_inv 
* No parameters

xinv_22 
+ int[21] int[22] vdd vss 
+ control_logic_inv 
* No parameters

xinv_23 
+ int[22] int[23] vdd vss 
+ control_logic_inv 
* No parameters

xinv_24 
+ int[23] int[24] vdd vss 
+ control_logic_inv 
* No parameters

xinv_25 
+ int[24] int[25] vdd vss 
+ control_logic_inv 
* No parameters

xinv_26 
+ int[25] int[26] vdd vss 
+ control_logic_inv 
* No parameters

xinv_27 
+ int[26] int[27] vdd vss 
+ control_logic_inv 
* No parameters

xinv_28 
+ int[27] int[28] vdd vss 
+ control_logic_inv 
* No parameters

xinv_29 
+ int[28] int[29] vdd vss 
+ control_logic_inv 
* No parameters

xinv_30 
+ int[29] int[30] vdd vss 
+ control_logic_inv 
* No parameters

xinv_31 
+ int[30] int[31] vdd vss 
+ control_logic_inv 
* No parameters

xinv_32 
+ int[31] int[32] vdd vss 
+ control_logic_inv 
* No parameters

xinv_33 
+ int[32] int[33] vdd vss 
+ control_logic_inv 
* No parameters

xinv_34 
+ int[33] int[34] vdd vss 
+ control_logic_inv 
* No parameters

xinv_35 
+ int[34] int[35] vdd vss 
+ control_logic_inv 
* No parameters

xinv_36 
+ int[35] int[36] vdd vss 
+ control_logic_inv 
* No parameters

xinv_37 
+ int[36] int[37] vdd vss 
+ control_logic_inv 
* No parameters

xinv_38 
+ int[37] int[38] vdd vss 
+ control_logic_inv 
* No parameters

xinv_39 
+ int[38] int[39] vdd vss 
+ control_logic_inv 
* No parameters

xinv_40 
+ int[39] int[40] vdd vss 
+ control_logic_inv 
* No parameters

xinv_41 
+ int[40] int[41] vdd vss 
+ control_logic_inv 
* No parameters

xinv_42 
+ int[41] int[42] vdd vss 
+ control_logic_inv 
* No parameters

xinv_43 
+ int[42] int[43] vdd vss 
+ control_logic_inv 
* No parameters

xinv_44 
+ int[43] dout vdd vss 
+ control_logic_inv 
* No parameters

.ENDS

.SUBCKT sramgen_sram_64x32m4w32_replica_v1 
+ vdd vss clk din[31] din[30] din[29] din[28] din[27] din[26] din[25] din[24] din[23] din[22] din[21] din[20] din[19] din[18] din[17] din[16] din[15] din[14] din[13] din[12] din[11] din[10] din[9] din[8] din[7] din[6] din[5] din[4] din[3] din[2] din[1] din[0] dout[31] dout[30] dout[29] dout[28] dout[27] dout[26] dout[25] dout[24] dout[23] dout[22] dout[21] dout[20] dout[19] dout[18] dout[17] dout[16] dout[15] dout[14] dout[13] dout[12] dout[11] dout[10] dout[9] dout[8] dout[7] dout[6] dout[5] dout[4] dout[3] dout[2] dout[1] dout[0] we addr[5] addr[4] addr[3] addr[2] addr[1] addr[0] 

xdin_dffs 
+ vdd vss clk din[31] din[30] din[29] din[28] din[27] din[26] din[25] din[24] din[23] din[22] din[21] din[20] din[19] din[18] din[17] din[16] din[15] din[14] din[13] din[12] din[11] din[10] din[9] din[8] din[7] din[6] din[5] din[4] din[3] din[2] din[1] din[0] bank_din[31] bank_din[30] bank_din[29] bank_din[28] bank_din[27] bank_din[26] bank_din[25] bank_din[24] bank_din[23] bank_din[22] bank_din[21] bank_din[20] bank_din[19] bank_din[18] bank_din[17] bank_din[16] bank_din[15] bank_din[14] bank_din[13] bank_din[12] bank_din[11] bank_din[10] bank_din[9] bank_din[8] bank_din[7] bank_din[6] bank_din[5] bank_din[4] bank_din[3] bank_din[2] bank_din[1] bank_din[0] dff_din_b[31] dff_din_b[30] dff_din_b[29] dff_din_b[28] dff_din_b[27] dff_din_b[26] dff_din_b[25] dff_din_b[24] dff_din_b[23] dff_din_b[22] dff_din_b[21] dff_din_b[20] dff_din_b[19] dff_din_b[18] dff_din_b[17] dff_din_b[16] dff_din_b[15] dff_din_b[14] dff_din_b[13] dff_din_b[12] dff_din_b[11] dff_din_b[10] dff_din_b[9] dff_din_b[8] dff_din_b[7] dff_din_b[6] dff_din_b[5] dff_din_b[4] dff_din_b[3] dff_din_b[2] dff_din_b[1] dff_din_b[0] 
+ data_dff_array 
* No parameters

xaddr_dffs 
+ vdd vss clk addr[5] addr[4] addr[3] addr[2] addr[1] addr[0] bank_addr[5] bank_addr[4] bank_addr[3] bank_addr[2] bank_addr[1] bank_addr[0] bank_addr_b[5] bank_addr_b[4] bank_addr_b[3] bank_addr_b[2] bank_addr_b[1] bank_addr_b[0] 
+ addr_dff_array 
* No parameters

xwe_dff 
+ vdd vss clk we bank_we bank_we_b 
+ openram_dff 
* No parameters

xdecoder 
+ vdd vss bank_addr[5] bank_addr[4] bank_addr[3] bank_addr[2] bank_addr_b[5] bank_addr_b[4] bank_addr_b[3] bank_addr_b[2] wl_data[15] wl_data[14] wl_data[13] wl_data[12] wl_data[11] wl_data[10] wl_data[9] wl_data[8] wl_data[7] wl_data[6] wl_data[5] wl_data[4] wl_data[3] wl_data[2] wl_data[1] wl_data[0] wl_data_b[15] wl_data_b[14] wl_data_b[13] wl_data_b[12] wl_data_b[11] wl_data_b[10] wl_data_b[9] wl_data_b[8] wl_data_b[7] wl_data_b[6] wl_data_b[5] wl_data_b[4] wl_data_b[3] wl_data_b[2] wl_data_b[1] wl_data_b[0] 
+ hierarchical_decoder 
* No parameters

xwl_driver_array 
+ vdd vss wl_data[15] wl_data[14] wl_data[13] wl_data[12] wl_data[11] wl_data[10] wl_data[9] wl_data[8] wl_data[7] wl_data[6] wl_data[5] wl_data[4] wl_data[3] wl_data[2] wl_data[1] wl_data[0] wl_en wl[15] wl[14] wl[13] wl[12] wl[11] wl[10] wl[9] wl[8] wl[7] wl[6] wl[5] wl[4] wl[3] wl[2] wl[1] wl[0] 
+ wordline_driver_array 
* No parameters

xbitcells 
+ vdd vss bl[127] bl[126] bl[125] bl[124] bl[123] bl[122] bl[121] bl[120] bl[119] bl[118] bl[117] bl[116] bl[115] bl[114] bl[113] bl[112] bl[111] bl[110] bl[109] bl[108] bl[107] bl[106] bl[105] bl[104] bl[103] bl[102] bl[101] bl[100] bl[99] bl[98] bl[97] bl[96] bl[95] bl[94] bl[93] bl[92] bl[91] bl[90] bl[89] bl[88] bl[87] bl[86] bl[85] bl[84] bl[83] bl[82] bl[81] bl[80] bl[79] bl[78] bl[77] bl[76] bl[75] bl[74] bl[73] bl[72] bl[71] bl[70] bl[69] bl[68] bl[67] bl[66] bl[65] bl[64] bl[63] bl[62] bl[61] bl[60] bl[59] bl[58] bl[57] bl[56] bl[55] bl[54] bl[53] bl[52] bl[51] bl[50] bl[49] bl[48] bl[47] bl[46] bl[45] bl[44] bl[43] bl[42] bl[41] bl[40] bl[39] bl[38] bl[37] bl[36] bl[35] bl[34] bl[33] bl[32] bl[31] bl[30] bl[29] bl[28] bl[27] bl[26] bl[25] bl[24] bl[23] bl[22] bl[21] bl[20] bl[19] bl[18] bl[17] bl[16] bl[15] bl[14] bl[13] bl[12] bl[11] bl[10] bl[9] bl[8] bl[7] bl[6] bl[5] bl[4] bl[3] bl[2] bl[1] bl[0] br[127] br[126] br[125] br[124] br[123] br[122] br[121] br[120] br[119] br[118] br[117] br[116] br[115] br[114] br[113] br[112] br[111] br[110] br[109] br[108] br[107] br[106] br[105] br[104] br[103] br[102] br[101] br[100] br[99] br[98] br[97] br[96] br[95] br[94] br[93] br[92] br[91] br[90] br[89] br[88] br[87] br[86] br[85] br[84] br[83] br[82] br[81] br[80] br[79] br[78] br[77] br[76] br[75] br[74] br[73] br[72] br[71] br[70] br[69] br[68] br[67] br[66] br[65] br[64] br[63] br[62] br[61] br[60] br[59] br[58] br[57] br[56] br[55] br[54] br[53] br[52] br[51] br[50] br[49] br[48] br[47] br[46] br[45] br[44] br[43] br[42] br[41] br[40] br[39] br[38] br[37] br[36] br[35] br[34] br[33] br[32] br[31] br[30] br[29] br[28] br[27] br[26] br[25] br[24] br[23] br[22] br[21] br[20] br[19] br[18] br[17] br[16] br[15] br[14] br[13] br[12] br[11] br[10] br[9] br[8] br[7] br[6] br[5] br[4] br[3] br[2] br[1] br[0] wl[15] wl[14] wl[13] wl[12] wl[11] wl[10] wl[9] wl[8] wl[7] wl[6] wl[5] wl[4] wl[3] wl[2] wl[1] wl[0] vss vdd rbl rbr 
+ bitcell_array 
* No parameters

xprecharge_array 
+ vdd pc_b rbl bl[127] bl[126] bl[125] bl[124] bl[123] bl[122] bl[121] bl[120] bl[119] bl[118] bl[117] bl[116] bl[115] bl[114] bl[113] bl[112] bl[111] bl[110] bl[109] bl[108] bl[107] bl[106] bl[105] bl[104] bl[103] bl[102] bl[101] bl[100] bl[99] bl[98] bl[97] bl[96] bl[95] bl[94] bl[93] bl[92] bl[91] bl[90] bl[89] bl[88] bl[87] bl[86] bl[85] bl[84] bl[83] bl[82] bl[81] bl[80] bl[79] bl[78] bl[77] bl[76] bl[75] bl[74] bl[73] bl[72] bl[71] bl[70] bl[69] bl[68] bl[67] bl[66] bl[65] bl[64] bl[63] bl[62] bl[61] bl[60] bl[59] bl[58] bl[57] bl[56] bl[55] bl[54] bl[53] bl[52] bl[51] bl[50] bl[49] bl[48] bl[47] bl[46] bl[45] bl[44] bl[43] bl[42] bl[41] bl[40] bl[39] bl[38] bl[37] bl[36] bl[35] bl[34] bl[33] bl[32] bl[31] bl[30] bl[29] bl[28] bl[27] bl[26] bl[25] bl[24] bl[23] bl[22] bl[21] bl[20] bl[19] bl[18] bl[17] bl[16] bl[15] bl[14] bl[13] bl[12] bl[11] bl[10] bl[9] bl[8] bl[7] bl[6] bl[5] bl[4] bl[3] bl[2] bl[1] bl[0]  rbr br[127] br[126] br[125] br[124] br[123] br[122] br[121] br[120] br[119] br[118] br[117] br[116] br[115] br[114] br[113] br[112] br[111] br[110] br[109] br[108] br[107] br[106] br[105] br[104] br[103] br[102] br[101] br[100] br[99] br[98] br[97] br[96] br[95] br[94] br[93] br[92] br[91] br[90] br[89] br[88] br[87] br[86] br[85] br[84] br[83] br[82] br[81] br[80] br[79] br[78] br[77] br[76] br[75] br[74] br[73] br[72] br[71] br[70] br[69] br[68] br[67] br[66] br[65] br[64] br[63] br[62] br[61] br[60] br[59] br[58] br[57] br[56] br[55] br[54] br[53] br[52] br[51] br[50] br[49] br[48] br[47] br[46] br[45] br[44] br[43] br[42] br[41] br[40] br[39] br[38] br[37] br[36] br[35] br[34] br[33] br[32] br[31] br[30] br[29] br[28] br[27] br[26] br[25] br[24] br[23] br[22] br[21] br[20] br[19] br[18] br[17] br[16] br[15] br[14] br[13] br[12] br[11] br[10] br[9] br[8] br[7] br[6] br[5] br[4] br[3] br[2] br[1] br[0]  
+ precharge_array 
* No parameters

xwrite_mux_array 
+ write_driver_en[3] write_driver_en[2] write_driver_en[1] write_driver_en[0] bank_din[31] bank_din[30] bank_din[29] bank_din[28] bank_din[27] bank_din[26] bank_din[25] bank_din[24] bank_din[23] bank_din[22] bank_din[21] bank_din[20] bank_din[19] bank_din[18] bank_din[17] bank_din[16] bank_din[15] bank_din[14] bank_din[13] bank_din[12] bank_din[11] bank_din[10] bank_din[9] bank_din[8] bank_din[7] bank_din[6] bank_din[5] bank_din[4] bank_din[3] bank_din[2] bank_din[1] bank_din[0] bank_din_b[31] bank_din_b[30] bank_din_b[29] bank_din_b[28] bank_din_b[27] bank_din_b[26] bank_din_b[25] bank_din_b[24] bank_din_b[23] bank_din_b[22] bank_din_b[21] bank_din_b[20] bank_din_b[19] bank_din_b[18] bank_din_b[17] bank_din_b[16] bank_din_b[15] bank_din_b[14] bank_din_b[13] bank_din_b[12] bank_din_b[11] bank_din_b[10] bank_din_b[9] bank_din_b[8] bank_din_b[7] bank_din_b[6] bank_din_b[5] bank_din_b[4] bank_din_b[3] bank_din_b[2] bank_din_b[1] bank_din_b[0] bl[127] bl[126] bl[125] bl[124] bl[123] bl[122] bl[121] bl[120] bl[119] bl[118] bl[117] bl[116] bl[115] bl[114] bl[113] bl[112] bl[111] bl[110] bl[109] bl[108] bl[107] bl[106] bl[105] bl[104] bl[103] bl[102] bl[101] bl[100] bl[99] bl[98] bl[97] bl[96] bl[95] bl[94] bl[93] bl[92] bl[91] bl[90] bl[89] bl[88] bl[87] bl[86] bl[85] bl[84] bl[83] bl[82] bl[81] bl[80] bl[79] bl[78] bl[77] bl[76] bl[75] bl[74] bl[73] bl[72] bl[71] bl[70] bl[69] bl[68] bl[67] bl[66] bl[65] bl[64] bl[63] bl[62] bl[61] bl[60] bl[59] bl[58] bl[57] bl[56] bl[55] bl[54] bl[53] bl[52] bl[51] bl[50] bl[49] bl[48] bl[47] bl[46] bl[45] bl[44] bl[43] bl[42] bl[41] bl[40] bl[39] bl[38] bl[37] bl[36] bl[35] bl[34] bl[33] bl[32] bl[31] bl[30] bl[29] bl[28] bl[27] bl[26] bl[25] bl[24] bl[23] bl[22] bl[21] bl[20] bl[19] bl[18] bl[17] bl[16] bl[15] bl[14] bl[13] bl[12] bl[11] bl[10] bl[9] bl[8] bl[7] bl[6] bl[5] bl[4] bl[3] bl[2] bl[1] bl[0] br[127] br[126] br[125] br[124] br[123] br[122] br[121] br[120] br[119] br[118] br[117] br[116] br[115] br[114] br[113] br[112] br[111] br[110] br[109] br[108] br[107] br[106] br[105] br[104] br[103] br[102] br[101] br[100] br[99] br[98] br[97] br[96] br[95] br[94] br[93] br[92] br[91] br[90] br[89] br[88] br[87] br[86] br[85] br[84] br[83] br[82] br[81] br[80] br[79] br[78] br[77] br[76] br[75] br[74] br[73] br[72] br[71] br[70] br[69] br[68] br[67] br[66] br[65] br[64] br[63] br[62] br[61] br[60] br[59] br[58] br[57] br[56] br[55] br[54] br[53] br[52] br[51] br[50] br[49] br[48] br[47] br[46] br[45] br[44] br[43] br[42] br[41] br[40] br[39] br[38] br[37] br[36] br[35] br[34] br[33] br[32] br[31] br[30] br[29] br[28] br[27] br[26] br[25] br[24] br[23] br[22] br[21] br[20] br[19] br[18] br[17] br[16] br[15] br[14] br[13] br[12] br[11] br[10] br[9] br[8] br[7] br[6] br[5] br[4] br[3] br[2] br[1] br[0] vss 
+ write_mux_array 
* No parameters

xread_mux_array 
+ col_sel_b[3] col_sel_b[2] col_sel_b[1] col_sel_b[0] bl[127] bl[126] bl[125] bl[124] bl[123] bl[122] bl[121] bl[120] bl[119] bl[118] bl[117] bl[116] bl[115] bl[114] bl[113] bl[112] bl[111] bl[110] bl[109] bl[108] bl[107] bl[106] bl[105] bl[104] bl[103] bl[102] bl[101] bl[100] bl[99] bl[98] bl[97] bl[96] bl[95] bl[94] bl[93] bl[92] bl[91] bl[90] bl[89] bl[88] bl[87] bl[86] bl[85] bl[84] bl[83] bl[82] bl[81] bl[80] bl[79] bl[78] bl[77] bl[76] bl[75] bl[74] bl[73] bl[72] bl[71] bl[70] bl[69] bl[68] bl[67] bl[66] bl[65] bl[64] bl[63] bl[62] bl[61] bl[60] bl[59] bl[58] bl[57] bl[56] bl[55] bl[54] bl[53] bl[52] bl[51] bl[50] bl[49] bl[48] bl[47] bl[46] bl[45] bl[44] bl[43] bl[42] bl[41] bl[40] bl[39] bl[38] bl[37] bl[36] bl[35] bl[34] bl[33] bl[32] bl[31] bl[30] bl[29] bl[28] bl[27] bl[26] bl[25] bl[24] bl[23] bl[22] bl[21] bl[20] bl[19] bl[18] bl[17] bl[16] bl[15] bl[14] bl[13] bl[12] bl[11] bl[10] bl[9] bl[8] bl[7] bl[6] bl[5] bl[4] bl[3] bl[2] bl[1] bl[0] br[127] br[126] br[125] br[124] br[123] br[122] br[121] br[120] br[119] br[118] br[117] br[116] br[115] br[114] br[113] br[112] br[111] br[110] br[109] br[108] br[107] br[106] br[105] br[104] br[103] br[102] br[101] br[100] br[99] br[98] br[97] br[96] br[95] br[94] br[93] br[92] br[91] br[90] br[89] br[88] br[87] br[86] br[85] br[84] br[83] br[82] br[81] br[80] br[79] br[78] br[77] br[76] br[75] br[74] br[73] br[72] br[71] br[70] br[69] br[68] br[67] br[66] br[65] br[64] br[63] br[62] br[61] br[60] br[59] br[58] br[57] br[56] br[55] br[54] br[53] br[52] br[51] br[50] br[49] br[48] br[47] br[46] br[45] br[44] br[43] br[42] br[41] br[40] br[39] br[38] br[37] br[36] br[35] br[34] br[33] br[32] br[31] br[30] br[29] br[28] br[27] br[26] br[25] br[24] br[23] br[22] br[21] br[20] br[19] br[18] br[17] br[16] br[15] br[14] br[13] br[12] br[11] br[10] br[9] br[8] br[7] br[6] br[5] br[4] br[3] br[2] br[1] br[0] bl_read[31] bl_read[30] bl_read[29] bl_read[28] bl_read[27] bl_read[26] bl_read[25] bl_read[24] bl_read[23] bl_read[22] bl_read[21] bl_read[20] bl_read[19] bl_read[18] bl_read[17] bl_read[16] bl_read[15] bl_read[14] bl_read[13] bl_read[12] bl_read[11] bl_read[10] bl_read[9] bl_read[8] bl_read[7] bl_read[6] bl_read[5] bl_read[4] bl_read[3] bl_read[2] bl_read[1] bl_read[0] br_read[31] br_read[30] br_read[29] br_read[28] br_read[27] br_read[26] br_read[25] br_read[24] br_read[23] br_read[22] br_read[21] br_read[20] br_read[19] br_read[18] br_read[17] br_read[16] br_read[15] br_read[14] br_read[13] br_read[12] br_read[11] br_read[10] br_read[9] br_read[8] br_read[7] br_read[6] br_read[5] br_read[4] br_read[3] br_read[2] br_read[1] br_read[0] vdd 
+ read_mux_array 
* No parameters

xcol_inv_array 
+ bank_din[31] bank_din[30] bank_din[29] bank_din[28] bank_din[27] bank_din[26] bank_din[25] bank_din[24] bank_din[23] bank_din[22] bank_din[21] bank_din[20] bank_din[19] bank_din[18] bank_din[17] bank_din[16] bank_din[15] bank_din[14] bank_din[13] bank_din[12] bank_din[11] bank_din[10] bank_din[9] bank_din[8] bank_din[7] bank_din[6] bank_din[5] bank_din[4] bank_din[3] bank_din[2] bank_din[1] bank_din[0] bank_din_b[31] bank_din_b[30] bank_din_b[29] bank_din_b[28] bank_din_b[27] bank_din_b[26] bank_din_b[25] bank_din_b[24] bank_din_b[23] bank_din_b[22] bank_din_b[21] bank_din_b[20] bank_din_b[19] bank_din_b[18] bank_din_b[17] bank_din_b[16] bank_din_b[15] bank_din_b[14] bank_din_b[13] bank_din_b[12] bank_din_b[11] bank_din_b[10] bank_din_b[9] bank_din_b[8] bank_din_b[7] bank_din_b[6] bank_din_b[5] bank_din_b[4] bank_din_b[3] bank_din_b[2] bank_din_b[1] bank_din_b[0] vdd vss 
+ col_inv_array 
* No parameters

xsense_amp_array 
+ vdd vss sense_amp_en bl_read[31] bl_read[30] bl_read[29] bl_read[28] bl_read[27] bl_read[26] bl_read[25] bl_read[24] bl_read[23] bl_read[22] bl_read[21] bl_read[20] bl_read[19] bl_read[18] bl_read[17] bl_read[16] bl_read[15] bl_read[14] bl_read[13] bl_read[12] bl_read[11] bl_read[10] bl_read[9] bl_read[8] bl_read[7] bl_read[6] bl_read[5] bl_read[4] bl_read[3] bl_read[2] bl_read[1] bl_read[0] br_read[31] br_read[30] br_read[29] br_read[28] br_read[27] br_read[26] br_read[25] br_read[24] br_read[23] br_read[22] br_read[21] br_read[20] br_read[19] br_read[18] br_read[17] br_read[16] br_read[15] br_read[14] br_read[13] br_read[12] br_read[11] br_read[10] br_read[9] br_read[8] br_read[7] br_read[6] br_read[5] br_read[4] br_read[3] br_read[2] br_read[1] br_read[0] sa_outp[31] sa_outp[30] sa_outp[29] sa_outp[28] sa_outp[27] sa_outp[26] sa_outp[25] sa_outp[24] sa_outp[23] sa_outp[22] sa_outp[21] sa_outp[20] sa_outp[19] sa_outp[18] sa_outp[17] sa_outp[16] sa_outp[15] sa_outp[14] sa_outp[13] sa_outp[12] sa_outp[11] sa_outp[10] sa_outp[9] sa_outp[8] sa_outp[7] sa_outp[6] sa_outp[5] sa_outp[4] sa_outp[3] sa_outp[2] sa_outp[1] sa_outp[0] sa_outn[31] sa_outn[30] sa_outn[29] sa_outn[28] sa_outn[27] sa_outn[26] sa_outn[25] sa_outn[24] sa_outn[23] sa_outn[22] sa_outn[21] sa_outn[20] sa_outn[19] sa_outn[18] sa_outn[17] sa_outn[16] sa_outn[15] sa_outn[14] sa_outn[13] sa_outn[12] sa_outn[11] sa_outn[10] sa_outn[9] sa_outn[8] sa_outn[7] sa_outn[6] sa_outn[5] sa_outn[4] sa_outn[3] sa_outn[2] sa_outn[1] sa_outn[0] 
+ sense_amp_array 
* No parameters

xdout_buf_array 
+ sa_outp[31] sa_outp[30] sa_outp[29] sa_outp[28] sa_outp[27] sa_outp[26] sa_outp[25] sa_outp[24] sa_outp[23] sa_outp[22] sa_outp[21] sa_outp[20] sa_outp[19] sa_outp[18] sa_outp[17] sa_outp[16] sa_outp[15] sa_outp[14] sa_outp[13] sa_outp[12] sa_outp[11] sa_outp[10] sa_outp[9] sa_outp[8] sa_outp[7] sa_outp[6] sa_outp[5] sa_outp[4] sa_outp[3] sa_outp[2] sa_outp[1] sa_outp[0] sa_outn[31] sa_outn[30] sa_outn[29] sa_outn[28] sa_outn[27] sa_outn[26] sa_outn[25] sa_outn[24] sa_outn[23] sa_outn[22] sa_outn[21] sa_outn[20] sa_outn[19] sa_outn[18] sa_outn[17] sa_outn[16] sa_outn[15] sa_outn[14] sa_outn[13] sa_outn[12] sa_outn[11] sa_outn[10] sa_outn[9] sa_outn[8] sa_outn[7] sa_outn[6] sa_outn[5] sa_outn[4] sa_outn[3] sa_outn[2] sa_outn[1] sa_outn[0] dout[31] dout[30] dout[29] dout[28] dout[27] dout[26] dout[25] dout[24] dout[23] dout[22] dout[21] dout[20] dout[19] dout[18] dout[17] dout[16] dout[15] dout[14] dout[13] dout[12] dout[11] dout[10] dout[9] dout[8] dout[7] dout[6] dout[5] dout[4] dout[3] dout[2] dout[1] dout[0] dout_b[31] dout_b[30] dout_b[29] dout_b[28] dout_b[27] dout_b[26] dout_b[25] dout_b[24] dout_b[23] dout_b[22] dout_b[21] dout_b[20] dout_b[19] dout_b[18] dout_b[17] dout_b[16] dout_b[15] dout_b[14] dout_b[13] dout_b[12] dout_b[11] dout_b[10] dout_b[9] dout_b[8] dout_b[7] dout_b[6] dout_b[5] dout_b[4] dout_b[3] dout_b[2] dout_b[1] dout_b[0] vdd vss 
+ dout_buf_array 
* No parameters

xcontrol_logic 
+ clk bank_we rbl pc_b wl_en wr_en sense_amp_en vdd vss 
+ sramgen_control_replica_v1 
* No parameters

xcolumn_decoder 
+ vdd vss bank_addr[1] bank_addr[0] bank_addr_b[1] bank_addr_b[0] col_sel[3] col_sel[2] col_sel[1] col_sel[0] col_sel_b[3] col_sel_b[2] col_sel_b[1] col_sel_b[0] 
+ column_decoder 
* No parameters

xwe_control 
+ wr_en col_sel[3] col_sel[2] col_sel[1] col_sel[0] write_driver_en[3] write_driver_en[2] write_driver_en[1] write_driver_en[0] vdd vss 
+ we_control 
* No parameters

.ENDS

