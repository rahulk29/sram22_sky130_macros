* circuit.Package sramgen_sramgen_sram_1024x32m8w8_replica_v1
* Written by SpiceNetlister
* 

.SUBCKT hierarchical_decoder_nand_2 
+ gnd vdd a b c y 

xn1 
+ x1 a gnd gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='3.2' l='0.15' 

xn2 
+ x2 b x1 gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='3.2' l='0.15' 

xn3 
+ y c x2 gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='3.2' l='0.15' 

xp1 
+ y a vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.4' l='0.15' 

xp2 
+ y b vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.4' l='0.15' 

xp3 
+ y c vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.4' l='0.15' 

.ENDS

.SUBCKT hierarchical_decoder_inv_3 
+ gnd vdd din din_b 

xn 
+ din_b din gnd gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='1.6' l='0.15' 

xp 
+ din_b din vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.4' l='0.15' 

.ENDS

.SUBCKT hierarchical_decoder_nand_29 
+ gnd vdd a b y 

xn1 
+ x a gnd gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='3.2' l='0.15' 

xn2 
+ y b x gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='3.2' l='0.15' 

xp1 
+ y a vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.4' l='0.15' 

xp2 
+ y b vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.4' l='0.15' 

.ENDS

.SUBCKT hierarchical_decoder 
+ vdd gnd addr[6] addr[5] addr[4] addr[3] addr[2] addr[1] addr[0] addr_b[6] addr_b[5] addr_b[4] addr_b[3] addr_b[2] addr_b[1] addr_b[0] decode[127] decode[126] decode[125] decode[124] decode[123] decode[122] decode[121] decode[120] decode[119] decode[118] decode[117] decode[116] decode[115] decode[114] decode[113] decode[112] decode[111] decode[110] decode[109] decode[108] decode[107] decode[106] decode[105] decode[104] decode[103] decode[102] decode[101] decode[100] decode[99] decode[98] decode[97] decode[96] decode[95] decode[94] decode[93] decode[92] decode[91] decode[90] decode[89] decode[88] decode[87] decode[86] decode[85] decode[84] decode[83] decode[82] decode[81] decode[80] decode[79] decode[78] decode[77] decode[76] decode[75] decode[74] decode[73] decode[72] decode[71] decode[70] decode[69] decode[68] decode[67] decode[66] decode[65] decode[64] decode[63] decode[62] decode[61] decode[60] decode[59] decode[58] decode[57] decode[56] decode[55] decode[54] decode[53] decode[52] decode[51] decode[50] decode[49] decode[48] decode[47] decode[46] decode[45] decode[44] decode[43] decode[42] decode[41] decode[40] decode[39] decode[38] decode[37] decode[36] decode[35] decode[34] decode[33] decode[32] decode[31] decode[30] decode[29] decode[28] decode[27] decode[26] decode[25] decode[24] decode[23] decode[22] decode[21] decode[20] decode[19] decode[18] decode[17] decode[16] decode[15] decode[14] decode[13] decode[12] decode[11] decode[10] decode[9] decode[8] decode[7] decode[6] decode[5] decode[4] decode[3] decode[2] decode[1] decode[0] decode_b[127] decode_b[126] decode_b[125] decode_b[124] decode_b[123] decode_b[122] decode_b[121] decode_b[120] decode_b[119] decode_b[118] decode_b[117] decode_b[116] decode_b[115] decode_b[114] decode_b[113] decode_b[112] decode_b[111] decode_b[110] decode_b[109] decode_b[108] decode_b[107] decode_b[106] decode_b[105] decode_b[104] decode_b[103] decode_b[102] decode_b[101] decode_b[100] decode_b[99] decode_b[98] decode_b[97] decode_b[96] decode_b[95] decode_b[94] decode_b[93] decode_b[92] decode_b[91] decode_b[90] decode_b[89] decode_b[88] decode_b[87] decode_b[86] decode_b[85] decode_b[84] decode_b[83] decode_b[82] decode_b[81] decode_b[80] decode_b[79] decode_b[78] decode_b[77] decode_b[76] decode_b[75] decode_b[74] decode_b[73] decode_b[72] decode_b[71] decode_b[70] decode_b[69] decode_b[68] decode_b[67] decode_b[66] decode_b[65] decode_b[64] decode_b[63] decode_b[62] decode_b[61] decode_b[60] decode_b[59] decode_b[58] decode_b[57] decode_b[56] decode_b[55] decode_b[54] decode_b[53] decode_b[52] decode_b[51] decode_b[50] decode_b[49] decode_b[48] decode_b[47] decode_b[46] decode_b[45] decode_b[44] decode_b[43] decode_b[42] decode_b[41] decode_b[40] decode_b[39] decode_b[38] decode_b[37] decode_b[36] decode_b[35] decode_b[34] decode_b[33] decode_b[32] decode_b[31] decode_b[30] decode_b[29] decode_b[28] decode_b[27] decode_b[26] decode_b[25] decode_b[24] decode_b[23] decode_b[22] decode_b[21] decode_b[20] decode_b[19] decode_b[18] decode_b[17] decode_b[16] decode_b[15] decode_b[14] decode_b[13] decode_b[12] decode_b[11] decode_b[10] decode_b[9] decode_b[8] decode_b[7] decode_b[6] decode_b[5] decode_b[4] decode_b[3] decode_b[2] decode_b[1] decode_b[0] 

xnand_5 
+ gnd vdd addr_b[6] addr_b[5] addr_b[4] net_4 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_6 
+ gnd vdd net_4 predecode_1[0] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_8 
+ gnd vdd addr_b[6] addr_b[5] addr[4] net_7 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_9 
+ gnd vdd net_7 predecode_1[1] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_11 
+ gnd vdd addr_b[6] addr[5] addr_b[4] net_10 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_12 
+ gnd vdd net_10 predecode_1[2] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_14 
+ gnd vdd addr_b[6] addr[5] addr[4] net_13 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_15 
+ gnd vdd net_13 predecode_1[3] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_17 
+ gnd vdd addr[6] addr_b[5] addr_b[4] net_16 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_18 
+ gnd vdd net_16 predecode_1[4] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_20 
+ gnd vdd addr[6] addr_b[5] addr[4] net_19 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_21 
+ gnd vdd net_19 predecode_1[5] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_23 
+ gnd vdd addr[6] addr[5] addr_b[4] net_22 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_24 
+ gnd vdd net_22 predecode_1[6] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_26 
+ gnd vdd addr[6] addr[5] addr[4] net_25 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_27 
+ gnd vdd net_25 predecode_1[7] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_31 
+ gnd vdd addr_b[3] addr_b[2] net_30 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_32 
+ gnd vdd net_30 predecode_28[0] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_34 
+ gnd vdd addr_b[3] addr[2] net_33 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_35 
+ gnd vdd net_33 predecode_28[1] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_37 
+ gnd vdd addr[3] addr_b[2] net_36 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_38 
+ gnd vdd net_36 predecode_28[2] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_40 
+ gnd vdd addr[3] addr[2] net_39 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_41 
+ gnd vdd net_39 predecode_28[3] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_44 
+ gnd vdd addr_b[1] addr_b[0] net_43 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_45 
+ gnd vdd net_43 predecode_42[0] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_47 
+ gnd vdd addr_b[1] addr[0] net_46 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_48 
+ gnd vdd net_46 predecode_42[1] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_50 
+ gnd vdd addr[1] addr_b[0] net_49 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_51 
+ gnd vdd net_49 predecode_42[2] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_53 
+ gnd vdd addr[1] addr[0] net_52 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_54 
+ gnd vdd net_52 predecode_42[3] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_57 
+ gnd vdd predecode_28[0] predecode_42[0] net_56 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_58 
+ gnd vdd net_56 predecode_55[0] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_60 
+ gnd vdd predecode_28[0] predecode_42[1] net_59 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_61 
+ gnd vdd net_59 predecode_55[1] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_63 
+ gnd vdd predecode_28[0] predecode_42[2] net_62 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_64 
+ gnd vdd net_62 predecode_55[2] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_66 
+ gnd vdd predecode_28[0] predecode_42[3] net_65 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_67 
+ gnd vdd net_65 predecode_55[3] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_69 
+ gnd vdd predecode_28[1] predecode_42[0] net_68 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_70 
+ gnd vdd net_68 predecode_55[4] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_72 
+ gnd vdd predecode_28[1] predecode_42[1] net_71 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_73 
+ gnd vdd net_71 predecode_55[5] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_75 
+ gnd vdd predecode_28[1] predecode_42[2] net_74 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_76 
+ gnd vdd net_74 predecode_55[6] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_78 
+ gnd vdd predecode_28[1] predecode_42[3] net_77 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_79 
+ gnd vdd net_77 predecode_55[7] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_81 
+ gnd vdd predecode_28[2] predecode_42[0] net_80 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_82 
+ gnd vdd net_80 predecode_55[8] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_84 
+ gnd vdd predecode_28[2] predecode_42[1] net_83 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_85 
+ gnd vdd net_83 predecode_55[9] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_87 
+ gnd vdd predecode_28[2] predecode_42[2] net_86 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_88 
+ gnd vdd net_86 predecode_55[10] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_90 
+ gnd vdd predecode_28[2] predecode_42[3] net_89 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_91 
+ gnd vdd net_89 predecode_55[11] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_93 
+ gnd vdd predecode_28[3] predecode_42[0] net_92 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_94 
+ gnd vdd net_92 predecode_55[12] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_96 
+ gnd vdd predecode_28[3] predecode_42[1] net_95 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_97 
+ gnd vdd net_95 predecode_55[13] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_99 
+ gnd vdd predecode_28[3] predecode_42[2] net_98 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_100 
+ gnd vdd net_98 predecode_55[14] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_102 
+ gnd vdd predecode_28[3] predecode_42[3] net_101 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_103 
+ gnd vdd net_101 predecode_55[15] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_104 
+ gnd vdd predecode_1[0] predecode_55[0] decode_b[0] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_105 
+ gnd vdd decode_b[0] decode[0] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_106 
+ gnd vdd predecode_1[0] predecode_55[1] decode_b[1] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_107 
+ gnd vdd decode_b[1] decode[1] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_108 
+ gnd vdd predecode_1[0] predecode_55[2] decode_b[2] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_109 
+ gnd vdd decode_b[2] decode[2] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_110 
+ gnd vdd predecode_1[0] predecode_55[3] decode_b[3] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_111 
+ gnd vdd decode_b[3] decode[3] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_112 
+ gnd vdd predecode_1[0] predecode_55[4] decode_b[4] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_113 
+ gnd vdd decode_b[4] decode[4] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_114 
+ gnd vdd predecode_1[0] predecode_55[5] decode_b[5] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_115 
+ gnd vdd decode_b[5] decode[5] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_116 
+ gnd vdd predecode_1[0] predecode_55[6] decode_b[6] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_117 
+ gnd vdd decode_b[6] decode[6] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_118 
+ gnd vdd predecode_1[0] predecode_55[7] decode_b[7] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_119 
+ gnd vdd decode_b[7] decode[7] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_120 
+ gnd vdd predecode_1[0] predecode_55[8] decode_b[8] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_121 
+ gnd vdd decode_b[8] decode[8] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_122 
+ gnd vdd predecode_1[0] predecode_55[9] decode_b[9] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_123 
+ gnd vdd decode_b[9] decode[9] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_124 
+ gnd vdd predecode_1[0] predecode_55[10] decode_b[10] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_125 
+ gnd vdd decode_b[10] decode[10] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_126 
+ gnd vdd predecode_1[0] predecode_55[11] decode_b[11] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_127 
+ gnd vdd decode_b[11] decode[11] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_128 
+ gnd vdd predecode_1[0] predecode_55[12] decode_b[12] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_129 
+ gnd vdd decode_b[12] decode[12] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_130 
+ gnd vdd predecode_1[0] predecode_55[13] decode_b[13] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_131 
+ gnd vdd decode_b[13] decode[13] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_132 
+ gnd vdd predecode_1[0] predecode_55[14] decode_b[14] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_133 
+ gnd vdd decode_b[14] decode[14] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_134 
+ gnd vdd predecode_1[0] predecode_55[15] decode_b[15] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_135 
+ gnd vdd decode_b[15] decode[15] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_136 
+ gnd vdd predecode_1[1] predecode_55[0] decode_b[16] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_137 
+ gnd vdd decode_b[16] decode[16] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_138 
+ gnd vdd predecode_1[1] predecode_55[1] decode_b[17] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_139 
+ gnd vdd decode_b[17] decode[17] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_140 
+ gnd vdd predecode_1[1] predecode_55[2] decode_b[18] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_141 
+ gnd vdd decode_b[18] decode[18] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_142 
+ gnd vdd predecode_1[1] predecode_55[3] decode_b[19] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_143 
+ gnd vdd decode_b[19] decode[19] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_144 
+ gnd vdd predecode_1[1] predecode_55[4] decode_b[20] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_145 
+ gnd vdd decode_b[20] decode[20] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_146 
+ gnd vdd predecode_1[1] predecode_55[5] decode_b[21] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_147 
+ gnd vdd decode_b[21] decode[21] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_148 
+ gnd vdd predecode_1[1] predecode_55[6] decode_b[22] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_149 
+ gnd vdd decode_b[22] decode[22] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_150 
+ gnd vdd predecode_1[1] predecode_55[7] decode_b[23] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_151 
+ gnd vdd decode_b[23] decode[23] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_152 
+ gnd vdd predecode_1[1] predecode_55[8] decode_b[24] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_153 
+ gnd vdd decode_b[24] decode[24] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_154 
+ gnd vdd predecode_1[1] predecode_55[9] decode_b[25] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_155 
+ gnd vdd decode_b[25] decode[25] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_156 
+ gnd vdd predecode_1[1] predecode_55[10] decode_b[26] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_157 
+ gnd vdd decode_b[26] decode[26] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_158 
+ gnd vdd predecode_1[1] predecode_55[11] decode_b[27] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_159 
+ gnd vdd decode_b[27] decode[27] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_160 
+ gnd vdd predecode_1[1] predecode_55[12] decode_b[28] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_161 
+ gnd vdd decode_b[28] decode[28] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_162 
+ gnd vdd predecode_1[1] predecode_55[13] decode_b[29] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_163 
+ gnd vdd decode_b[29] decode[29] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_164 
+ gnd vdd predecode_1[1] predecode_55[14] decode_b[30] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_165 
+ gnd vdd decode_b[30] decode[30] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_166 
+ gnd vdd predecode_1[1] predecode_55[15] decode_b[31] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_167 
+ gnd vdd decode_b[31] decode[31] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_168 
+ gnd vdd predecode_1[2] predecode_55[0] decode_b[32] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_169 
+ gnd vdd decode_b[32] decode[32] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_170 
+ gnd vdd predecode_1[2] predecode_55[1] decode_b[33] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_171 
+ gnd vdd decode_b[33] decode[33] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_172 
+ gnd vdd predecode_1[2] predecode_55[2] decode_b[34] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_173 
+ gnd vdd decode_b[34] decode[34] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_174 
+ gnd vdd predecode_1[2] predecode_55[3] decode_b[35] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_175 
+ gnd vdd decode_b[35] decode[35] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_176 
+ gnd vdd predecode_1[2] predecode_55[4] decode_b[36] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_177 
+ gnd vdd decode_b[36] decode[36] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_178 
+ gnd vdd predecode_1[2] predecode_55[5] decode_b[37] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_179 
+ gnd vdd decode_b[37] decode[37] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_180 
+ gnd vdd predecode_1[2] predecode_55[6] decode_b[38] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_181 
+ gnd vdd decode_b[38] decode[38] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_182 
+ gnd vdd predecode_1[2] predecode_55[7] decode_b[39] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_183 
+ gnd vdd decode_b[39] decode[39] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_184 
+ gnd vdd predecode_1[2] predecode_55[8] decode_b[40] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_185 
+ gnd vdd decode_b[40] decode[40] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_186 
+ gnd vdd predecode_1[2] predecode_55[9] decode_b[41] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_187 
+ gnd vdd decode_b[41] decode[41] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_188 
+ gnd vdd predecode_1[2] predecode_55[10] decode_b[42] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_189 
+ gnd vdd decode_b[42] decode[42] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_190 
+ gnd vdd predecode_1[2] predecode_55[11] decode_b[43] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_191 
+ gnd vdd decode_b[43] decode[43] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_192 
+ gnd vdd predecode_1[2] predecode_55[12] decode_b[44] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_193 
+ gnd vdd decode_b[44] decode[44] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_194 
+ gnd vdd predecode_1[2] predecode_55[13] decode_b[45] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_195 
+ gnd vdd decode_b[45] decode[45] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_196 
+ gnd vdd predecode_1[2] predecode_55[14] decode_b[46] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_197 
+ gnd vdd decode_b[46] decode[46] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_198 
+ gnd vdd predecode_1[2] predecode_55[15] decode_b[47] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_199 
+ gnd vdd decode_b[47] decode[47] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_200 
+ gnd vdd predecode_1[3] predecode_55[0] decode_b[48] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_201 
+ gnd vdd decode_b[48] decode[48] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_202 
+ gnd vdd predecode_1[3] predecode_55[1] decode_b[49] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_203 
+ gnd vdd decode_b[49] decode[49] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_204 
+ gnd vdd predecode_1[3] predecode_55[2] decode_b[50] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_205 
+ gnd vdd decode_b[50] decode[50] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_206 
+ gnd vdd predecode_1[3] predecode_55[3] decode_b[51] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_207 
+ gnd vdd decode_b[51] decode[51] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_208 
+ gnd vdd predecode_1[3] predecode_55[4] decode_b[52] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_209 
+ gnd vdd decode_b[52] decode[52] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_210 
+ gnd vdd predecode_1[3] predecode_55[5] decode_b[53] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_211 
+ gnd vdd decode_b[53] decode[53] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_212 
+ gnd vdd predecode_1[3] predecode_55[6] decode_b[54] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_213 
+ gnd vdd decode_b[54] decode[54] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_214 
+ gnd vdd predecode_1[3] predecode_55[7] decode_b[55] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_215 
+ gnd vdd decode_b[55] decode[55] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_216 
+ gnd vdd predecode_1[3] predecode_55[8] decode_b[56] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_217 
+ gnd vdd decode_b[56] decode[56] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_218 
+ gnd vdd predecode_1[3] predecode_55[9] decode_b[57] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_219 
+ gnd vdd decode_b[57] decode[57] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_220 
+ gnd vdd predecode_1[3] predecode_55[10] decode_b[58] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_221 
+ gnd vdd decode_b[58] decode[58] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_222 
+ gnd vdd predecode_1[3] predecode_55[11] decode_b[59] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_223 
+ gnd vdd decode_b[59] decode[59] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_224 
+ gnd vdd predecode_1[3] predecode_55[12] decode_b[60] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_225 
+ gnd vdd decode_b[60] decode[60] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_226 
+ gnd vdd predecode_1[3] predecode_55[13] decode_b[61] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_227 
+ gnd vdd decode_b[61] decode[61] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_228 
+ gnd vdd predecode_1[3] predecode_55[14] decode_b[62] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_229 
+ gnd vdd decode_b[62] decode[62] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_230 
+ gnd vdd predecode_1[3] predecode_55[15] decode_b[63] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_231 
+ gnd vdd decode_b[63] decode[63] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_232 
+ gnd vdd predecode_1[4] predecode_55[0] decode_b[64] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_233 
+ gnd vdd decode_b[64] decode[64] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_234 
+ gnd vdd predecode_1[4] predecode_55[1] decode_b[65] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_235 
+ gnd vdd decode_b[65] decode[65] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_236 
+ gnd vdd predecode_1[4] predecode_55[2] decode_b[66] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_237 
+ gnd vdd decode_b[66] decode[66] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_238 
+ gnd vdd predecode_1[4] predecode_55[3] decode_b[67] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_239 
+ gnd vdd decode_b[67] decode[67] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_240 
+ gnd vdd predecode_1[4] predecode_55[4] decode_b[68] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_241 
+ gnd vdd decode_b[68] decode[68] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_242 
+ gnd vdd predecode_1[4] predecode_55[5] decode_b[69] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_243 
+ gnd vdd decode_b[69] decode[69] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_244 
+ gnd vdd predecode_1[4] predecode_55[6] decode_b[70] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_245 
+ gnd vdd decode_b[70] decode[70] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_246 
+ gnd vdd predecode_1[4] predecode_55[7] decode_b[71] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_247 
+ gnd vdd decode_b[71] decode[71] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_248 
+ gnd vdd predecode_1[4] predecode_55[8] decode_b[72] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_249 
+ gnd vdd decode_b[72] decode[72] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_250 
+ gnd vdd predecode_1[4] predecode_55[9] decode_b[73] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_251 
+ gnd vdd decode_b[73] decode[73] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_252 
+ gnd vdd predecode_1[4] predecode_55[10] decode_b[74] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_253 
+ gnd vdd decode_b[74] decode[74] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_254 
+ gnd vdd predecode_1[4] predecode_55[11] decode_b[75] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_255 
+ gnd vdd decode_b[75] decode[75] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_256 
+ gnd vdd predecode_1[4] predecode_55[12] decode_b[76] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_257 
+ gnd vdd decode_b[76] decode[76] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_258 
+ gnd vdd predecode_1[4] predecode_55[13] decode_b[77] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_259 
+ gnd vdd decode_b[77] decode[77] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_260 
+ gnd vdd predecode_1[4] predecode_55[14] decode_b[78] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_261 
+ gnd vdd decode_b[78] decode[78] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_262 
+ gnd vdd predecode_1[4] predecode_55[15] decode_b[79] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_263 
+ gnd vdd decode_b[79] decode[79] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_264 
+ gnd vdd predecode_1[5] predecode_55[0] decode_b[80] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_265 
+ gnd vdd decode_b[80] decode[80] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_266 
+ gnd vdd predecode_1[5] predecode_55[1] decode_b[81] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_267 
+ gnd vdd decode_b[81] decode[81] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_268 
+ gnd vdd predecode_1[5] predecode_55[2] decode_b[82] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_269 
+ gnd vdd decode_b[82] decode[82] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_270 
+ gnd vdd predecode_1[5] predecode_55[3] decode_b[83] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_271 
+ gnd vdd decode_b[83] decode[83] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_272 
+ gnd vdd predecode_1[5] predecode_55[4] decode_b[84] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_273 
+ gnd vdd decode_b[84] decode[84] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_274 
+ gnd vdd predecode_1[5] predecode_55[5] decode_b[85] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_275 
+ gnd vdd decode_b[85] decode[85] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_276 
+ gnd vdd predecode_1[5] predecode_55[6] decode_b[86] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_277 
+ gnd vdd decode_b[86] decode[86] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_278 
+ gnd vdd predecode_1[5] predecode_55[7] decode_b[87] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_279 
+ gnd vdd decode_b[87] decode[87] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_280 
+ gnd vdd predecode_1[5] predecode_55[8] decode_b[88] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_281 
+ gnd vdd decode_b[88] decode[88] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_282 
+ gnd vdd predecode_1[5] predecode_55[9] decode_b[89] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_283 
+ gnd vdd decode_b[89] decode[89] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_284 
+ gnd vdd predecode_1[5] predecode_55[10] decode_b[90] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_285 
+ gnd vdd decode_b[90] decode[90] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_286 
+ gnd vdd predecode_1[5] predecode_55[11] decode_b[91] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_287 
+ gnd vdd decode_b[91] decode[91] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_288 
+ gnd vdd predecode_1[5] predecode_55[12] decode_b[92] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_289 
+ gnd vdd decode_b[92] decode[92] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_290 
+ gnd vdd predecode_1[5] predecode_55[13] decode_b[93] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_291 
+ gnd vdd decode_b[93] decode[93] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_292 
+ gnd vdd predecode_1[5] predecode_55[14] decode_b[94] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_293 
+ gnd vdd decode_b[94] decode[94] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_294 
+ gnd vdd predecode_1[5] predecode_55[15] decode_b[95] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_295 
+ gnd vdd decode_b[95] decode[95] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_296 
+ gnd vdd predecode_1[6] predecode_55[0] decode_b[96] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_297 
+ gnd vdd decode_b[96] decode[96] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_298 
+ gnd vdd predecode_1[6] predecode_55[1] decode_b[97] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_299 
+ gnd vdd decode_b[97] decode[97] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_300 
+ gnd vdd predecode_1[6] predecode_55[2] decode_b[98] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_301 
+ gnd vdd decode_b[98] decode[98] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_302 
+ gnd vdd predecode_1[6] predecode_55[3] decode_b[99] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_303 
+ gnd vdd decode_b[99] decode[99] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_304 
+ gnd vdd predecode_1[6] predecode_55[4] decode_b[100] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_305 
+ gnd vdd decode_b[100] decode[100] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_306 
+ gnd vdd predecode_1[6] predecode_55[5] decode_b[101] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_307 
+ gnd vdd decode_b[101] decode[101] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_308 
+ gnd vdd predecode_1[6] predecode_55[6] decode_b[102] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_309 
+ gnd vdd decode_b[102] decode[102] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_310 
+ gnd vdd predecode_1[6] predecode_55[7] decode_b[103] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_311 
+ gnd vdd decode_b[103] decode[103] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_312 
+ gnd vdd predecode_1[6] predecode_55[8] decode_b[104] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_313 
+ gnd vdd decode_b[104] decode[104] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_314 
+ gnd vdd predecode_1[6] predecode_55[9] decode_b[105] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_315 
+ gnd vdd decode_b[105] decode[105] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_316 
+ gnd vdd predecode_1[6] predecode_55[10] decode_b[106] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_317 
+ gnd vdd decode_b[106] decode[106] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_318 
+ gnd vdd predecode_1[6] predecode_55[11] decode_b[107] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_319 
+ gnd vdd decode_b[107] decode[107] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_320 
+ gnd vdd predecode_1[6] predecode_55[12] decode_b[108] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_321 
+ gnd vdd decode_b[108] decode[108] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_322 
+ gnd vdd predecode_1[6] predecode_55[13] decode_b[109] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_323 
+ gnd vdd decode_b[109] decode[109] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_324 
+ gnd vdd predecode_1[6] predecode_55[14] decode_b[110] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_325 
+ gnd vdd decode_b[110] decode[110] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_326 
+ gnd vdd predecode_1[6] predecode_55[15] decode_b[111] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_327 
+ gnd vdd decode_b[111] decode[111] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_328 
+ gnd vdd predecode_1[7] predecode_55[0] decode_b[112] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_329 
+ gnd vdd decode_b[112] decode[112] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_330 
+ gnd vdd predecode_1[7] predecode_55[1] decode_b[113] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_331 
+ gnd vdd decode_b[113] decode[113] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_332 
+ gnd vdd predecode_1[7] predecode_55[2] decode_b[114] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_333 
+ gnd vdd decode_b[114] decode[114] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_334 
+ gnd vdd predecode_1[7] predecode_55[3] decode_b[115] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_335 
+ gnd vdd decode_b[115] decode[115] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_336 
+ gnd vdd predecode_1[7] predecode_55[4] decode_b[116] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_337 
+ gnd vdd decode_b[116] decode[116] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_338 
+ gnd vdd predecode_1[7] predecode_55[5] decode_b[117] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_339 
+ gnd vdd decode_b[117] decode[117] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_340 
+ gnd vdd predecode_1[7] predecode_55[6] decode_b[118] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_341 
+ gnd vdd decode_b[118] decode[118] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_342 
+ gnd vdd predecode_1[7] predecode_55[7] decode_b[119] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_343 
+ gnd vdd decode_b[119] decode[119] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_344 
+ gnd vdd predecode_1[7] predecode_55[8] decode_b[120] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_345 
+ gnd vdd decode_b[120] decode[120] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_346 
+ gnd vdd predecode_1[7] predecode_55[9] decode_b[121] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_347 
+ gnd vdd decode_b[121] decode[121] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_348 
+ gnd vdd predecode_1[7] predecode_55[10] decode_b[122] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_349 
+ gnd vdd decode_b[122] decode[122] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_350 
+ gnd vdd predecode_1[7] predecode_55[11] decode_b[123] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_351 
+ gnd vdd decode_b[123] decode[123] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_352 
+ gnd vdd predecode_1[7] predecode_55[12] decode_b[124] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_353 
+ gnd vdd decode_b[124] decode[124] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_354 
+ gnd vdd predecode_1[7] predecode_55[13] decode_b[125] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_355 
+ gnd vdd decode_b[125] decode[125] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_356 
+ gnd vdd predecode_1[7] predecode_55[14] decode_b[126] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_357 
+ gnd vdd decode_b[126] decode[126] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_358 
+ gnd vdd predecode_1[7] predecode_55[15] decode_b[127] 
+ hierarchical_decoder_nand_29 
* No parameters

xinv_359 
+ gnd vdd decode_b[127] decode[127] 
+ hierarchical_decoder_inv_3 
* No parameters

.ENDS

.SUBCKT column_decoder_nand_1 
+ gnd vdd a b c y 

xn1 
+ x1 a gnd gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='3.2' l='0.15' 

xn2 
+ x2 b x1 gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='3.2' l='0.15' 

xn3 
+ y c x2 gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='3.2' l='0.15' 

xp1 
+ y a vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.4' l='0.15' 

xp2 
+ y b vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.4' l='0.15' 

xp3 
+ y c vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.4' l='0.15' 

.ENDS

.SUBCKT column_decoder_inv_2 
+ gnd vdd din din_b 

xn 
+ din_b din gnd gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='1.6' l='0.15' 

xp 
+ din_b din vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.4' l='0.15' 

.ENDS

.SUBCKT column_decoder 
+ vdd gnd addr[2] addr[1] addr[0] addr_b[2] addr_b[1] addr_b[0] decode[7] decode[6] decode[5] decode[4] decode[3] decode[2] decode[1] decode[0] decode_b[7] decode_b[6] decode_b[5] decode_b[4] decode_b[3] decode_b[2] decode_b[1] decode_b[0] 

xnand_3 
+ gnd vdd addr_b[2] addr_b[1] addr_b[0] decode_b[0] 
+ column_decoder_nand_1 
* No parameters

xinv_4 
+ gnd vdd decode_b[0] decode[0] 
+ column_decoder_inv_2 
* No parameters

xnand_5 
+ gnd vdd addr_b[2] addr_b[1] addr[0] decode_b[1] 
+ column_decoder_nand_1 
* No parameters

xinv_6 
+ gnd vdd decode_b[1] decode[1] 
+ column_decoder_inv_2 
* No parameters

xnand_7 
+ gnd vdd addr_b[2] addr[1] addr_b[0] decode_b[2] 
+ column_decoder_nand_1 
* No parameters

xinv_8 
+ gnd vdd decode_b[2] decode[2] 
+ column_decoder_inv_2 
* No parameters

xnand_9 
+ gnd vdd addr_b[2] addr[1] addr[0] decode_b[3] 
+ column_decoder_nand_1 
* No parameters

xinv_10 
+ gnd vdd decode_b[3] decode[3] 
+ column_decoder_inv_2 
* No parameters

xnand_11 
+ gnd vdd addr[2] addr_b[1] addr_b[0] decode_b[4] 
+ column_decoder_nand_1 
* No parameters

xinv_12 
+ gnd vdd decode_b[4] decode[4] 
+ column_decoder_inv_2 
* No parameters

xnand_13 
+ gnd vdd addr[2] addr_b[1] addr[0] decode_b[5] 
+ column_decoder_nand_1 
* No parameters

xinv_14 
+ gnd vdd decode_b[5] decode[5] 
+ column_decoder_inv_2 
* No parameters

xnand_15 
+ gnd vdd addr[2] addr[1] addr_b[0] decode_b[6] 
+ column_decoder_nand_1 
* No parameters

xinv_16 
+ gnd vdd decode_b[6] decode[6] 
+ column_decoder_inv_2 
* No parameters

xnand_17 
+ gnd vdd addr[2] addr[1] addr[0] decode_b[7] 
+ column_decoder_nand_1 
* No parameters

xinv_18 
+ gnd vdd decode_b[7] decode[7] 
+ column_decoder_inv_2 
* No parameters

.ENDS

.SUBCKT wordline_driver_and2_nand 
+ gnd vdd a b y 

xn1 
+ x a gnd gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='3.2' l='0.15' 

xn2 
+ y b x gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='3.2' l='0.15' 

xp1 
+ y a vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.4' l='0.15' 

xp2 
+ y b vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.4' l='0.15' 

.ENDS

.SUBCKT wordline_driver_and2_inv 
+ gnd vdd din din_b 

xn 
+ din_b din gnd gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='1.6' l='0.15' 

xp 
+ din_b din vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.4' l='0.15' 

.ENDS

.SUBCKT wordline_driver_and2 
+ a b y vdd vss 

xnand 
+ vss vdd a b tmp 
+ wordline_driver_and2_nand 
* No parameters

xinv 
+ vss vdd tmp y 
+ wordline_driver_and2_inv 
* No parameters

.ENDS

.SUBCKT wordline_driver 
+ vdd vss din wl_en wl 

xand2 
+ din wl_en wl vdd vss 
+ wordline_driver_and2 
* No parameters

.ENDS

.SUBCKT wordline_driver_array 
+ vdd vss din[127] din[126] din[125] din[124] din[123] din[122] din[121] din[120] din[119] din[118] din[117] din[116] din[115] din[114] din[113] din[112] din[111] din[110] din[109] din[108] din[107] din[106] din[105] din[104] din[103] din[102] din[101] din[100] din[99] din[98] din[97] din[96] din[95] din[94] din[93] din[92] din[91] din[90] din[89] din[88] din[87] din[86] din[85] din[84] din[83] din[82] din[81] din[80] din[79] din[78] din[77] din[76] din[75] din[74] din[73] din[72] din[71] din[70] din[69] din[68] din[67] din[66] din[65] din[64] din[63] din[62] din[61] din[60] din[59] din[58] din[57] din[56] din[55] din[54] din[53] din[52] din[51] din[50] din[49] din[48] din[47] din[46] din[45] din[44] din[43] din[42] din[41] din[40] din[39] din[38] din[37] din[36] din[35] din[34] din[33] din[32] din[31] din[30] din[29] din[28] din[27] din[26] din[25] din[24] din[23] din[22] din[21] din[20] din[19] din[18] din[17] din[16] din[15] din[14] din[13] din[12] din[11] din[10] din[9] din[8] din[7] din[6] din[5] din[4] din[3] din[2] din[1] din[0] wl_en wl[127] wl[126] wl[125] wl[124] wl[123] wl[122] wl[121] wl[120] wl[119] wl[118] wl[117] wl[116] wl[115] wl[114] wl[113] wl[112] wl[111] wl[110] wl[109] wl[108] wl[107] wl[106] wl[105] wl[104] wl[103] wl[102] wl[101] wl[100] wl[99] wl[98] wl[97] wl[96] wl[95] wl[94] wl[93] wl[92] wl[91] wl[90] wl[89] wl[88] wl[87] wl[86] wl[85] wl[84] wl[83] wl[82] wl[81] wl[80] wl[79] wl[78] wl[77] wl[76] wl[75] wl[74] wl[73] wl[72] wl[71] wl[70] wl[69] wl[68] wl[67] wl[66] wl[65] wl[64] wl[63] wl[62] wl[61] wl[60] wl[59] wl[58] wl[57] wl[56] wl[55] wl[54] wl[53] wl[52] wl[51] wl[50] wl[49] wl[48] wl[47] wl[46] wl[45] wl[44] wl[43] wl[42] wl[41] wl[40] wl[39] wl[38] wl[37] wl[36] wl[35] wl[34] wl[33] wl[32] wl[31] wl[30] wl[29] wl[28] wl[27] wl[26] wl[25] wl[24] wl[23] wl[22] wl[21] wl[20] wl[19] wl[18] wl[17] wl[16] wl[15] wl[14] wl[13] wl[12] wl[11] wl[10] wl[9] wl[8] wl[7] wl[6] wl[5] wl[4] wl[3] wl[2] wl[1] wl[0] 

xwl_driver_0 
+ vdd vss din[0] wl_en wl[0] 
+ wordline_driver 
* No parameters

xwl_driver_1 
+ vdd vss din[1] wl_en wl[1] 
+ wordline_driver 
* No parameters

xwl_driver_2 
+ vdd vss din[2] wl_en wl[2] 
+ wordline_driver 
* No parameters

xwl_driver_3 
+ vdd vss din[3] wl_en wl[3] 
+ wordline_driver 
* No parameters

xwl_driver_4 
+ vdd vss din[4] wl_en wl[4] 
+ wordline_driver 
* No parameters

xwl_driver_5 
+ vdd vss din[5] wl_en wl[5] 
+ wordline_driver 
* No parameters

xwl_driver_6 
+ vdd vss din[6] wl_en wl[6] 
+ wordline_driver 
* No parameters

xwl_driver_7 
+ vdd vss din[7] wl_en wl[7] 
+ wordline_driver 
* No parameters

xwl_driver_8 
+ vdd vss din[8] wl_en wl[8] 
+ wordline_driver 
* No parameters

xwl_driver_9 
+ vdd vss din[9] wl_en wl[9] 
+ wordline_driver 
* No parameters

xwl_driver_10 
+ vdd vss din[10] wl_en wl[10] 
+ wordline_driver 
* No parameters

xwl_driver_11 
+ vdd vss din[11] wl_en wl[11] 
+ wordline_driver 
* No parameters

xwl_driver_12 
+ vdd vss din[12] wl_en wl[12] 
+ wordline_driver 
* No parameters

xwl_driver_13 
+ vdd vss din[13] wl_en wl[13] 
+ wordline_driver 
* No parameters

xwl_driver_14 
+ vdd vss din[14] wl_en wl[14] 
+ wordline_driver 
* No parameters

xwl_driver_15 
+ vdd vss din[15] wl_en wl[15] 
+ wordline_driver 
* No parameters

xwl_driver_16 
+ vdd vss din[16] wl_en wl[16] 
+ wordline_driver 
* No parameters

xwl_driver_17 
+ vdd vss din[17] wl_en wl[17] 
+ wordline_driver 
* No parameters

xwl_driver_18 
+ vdd vss din[18] wl_en wl[18] 
+ wordline_driver 
* No parameters

xwl_driver_19 
+ vdd vss din[19] wl_en wl[19] 
+ wordline_driver 
* No parameters

xwl_driver_20 
+ vdd vss din[20] wl_en wl[20] 
+ wordline_driver 
* No parameters

xwl_driver_21 
+ vdd vss din[21] wl_en wl[21] 
+ wordline_driver 
* No parameters

xwl_driver_22 
+ vdd vss din[22] wl_en wl[22] 
+ wordline_driver 
* No parameters

xwl_driver_23 
+ vdd vss din[23] wl_en wl[23] 
+ wordline_driver 
* No parameters

xwl_driver_24 
+ vdd vss din[24] wl_en wl[24] 
+ wordline_driver 
* No parameters

xwl_driver_25 
+ vdd vss din[25] wl_en wl[25] 
+ wordline_driver 
* No parameters

xwl_driver_26 
+ vdd vss din[26] wl_en wl[26] 
+ wordline_driver 
* No parameters

xwl_driver_27 
+ vdd vss din[27] wl_en wl[27] 
+ wordline_driver 
* No parameters

xwl_driver_28 
+ vdd vss din[28] wl_en wl[28] 
+ wordline_driver 
* No parameters

xwl_driver_29 
+ vdd vss din[29] wl_en wl[29] 
+ wordline_driver 
* No parameters

xwl_driver_30 
+ vdd vss din[30] wl_en wl[30] 
+ wordline_driver 
* No parameters

xwl_driver_31 
+ vdd vss din[31] wl_en wl[31] 
+ wordline_driver 
* No parameters

xwl_driver_32 
+ vdd vss din[32] wl_en wl[32] 
+ wordline_driver 
* No parameters

xwl_driver_33 
+ vdd vss din[33] wl_en wl[33] 
+ wordline_driver 
* No parameters

xwl_driver_34 
+ vdd vss din[34] wl_en wl[34] 
+ wordline_driver 
* No parameters

xwl_driver_35 
+ vdd vss din[35] wl_en wl[35] 
+ wordline_driver 
* No parameters

xwl_driver_36 
+ vdd vss din[36] wl_en wl[36] 
+ wordline_driver 
* No parameters

xwl_driver_37 
+ vdd vss din[37] wl_en wl[37] 
+ wordline_driver 
* No parameters

xwl_driver_38 
+ vdd vss din[38] wl_en wl[38] 
+ wordline_driver 
* No parameters

xwl_driver_39 
+ vdd vss din[39] wl_en wl[39] 
+ wordline_driver 
* No parameters

xwl_driver_40 
+ vdd vss din[40] wl_en wl[40] 
+ wordline_driver 
* No parameters

xwl_driver_41 
+ vdd vss din[41] wl_en wl[41] 
+ wordline_driver 
* No parameters

xwl_driver_42 
+ vdd vss din[42] wl_en wl[42] 
+ wordline_driver 
* No parameters

xwl_driver_43 
+ vdd vss din[43] wl_en wl[43] 
+ wordline_driver 
* No parameters

xwl_driver_44 
+ vdd vss din[44] wl_en wl[44] 
+ wordline_driver 
* No parameters

xwl_driver_45 
+ vdd vss din[45] wl_en wl[45] 
+ wordline_driver 
* No parameters

xwl_driver_46 
+ vdd vss din[46] wl_en wl[46] 
+ wordline_driver 
* No parameters

xwl_driver_47 
+ vdd vss din[47] wl_en wl[47] 
+ wordline_driver 
* No parameters

xwl_driver_48 
+ vdd vss din[48] wl_en wl[48] 
+ wordline_driver 
* No parameters

xwl_driver_49 
+ vdd vss din[49] wl_en wl[49] 
+ wordline_driver 
* No parameters

xwl_driver_50 
+ vdd vss din[50] wl_en wl[50] 
+ wordline_driver 
* No parameters

xwl_driver_51 
+ vdd vss din[51] wl_en wl[51] 
+ wordline_driver 
* No parameters

xwl_driver_52 
+ vdd vss din[52] wl_en wl[52] 
+ wordline_driver 
* No parameters

xwl_driver_53 
+ vdd vss din[53] wl_en wl[53] 
+ wordline_driver 
* No parameters

xwl_driver_54 
+ vdd vss din[54] wl_en wl[54] 
+ wordline_driver 
* No parameters

xwl_driver_55 
+ vdd vss din[55] wl_en wl[55] 
+ wordline_driver 
* No parameters

xwl_driver_56 
+ vdd vss din[56] wl_en wl[56] 
+ wordline_driver 
* No parameters

xwl_driver_57 
+ vdd vss din[57] wl_en wl[57] 
+ wordline_driver 
* No parameters

xwl_driver_58 
+ vdd vss din[58] wl_en wl[58] 
+ wordline_driver 
* No parameters

xwl_driver_59 
+ vdd vss din[59] wl_en wl[59] 
+ wordline_driver 
* No parameters

xwl_driver_60 
+ vdd vss din[60] wl_en wl[60] 
+ wordline_driver 
* No parameters

xwl_driver_61 
+ vdd vss din[61] wl_en wl[61] 
+ wordline_driver 
* No parameters

xwl_driver_62 
+ vdd vss din[62] wl_en wl[62] 
+ wordline_driver 
* No parameters

xwl_driver_63 
+ vdd vss din[63] wl_en wl[63] 
+ wordline_driver 
* No parameters

xwl_driver_64 
+ vdd vss din[64] wl_en wl[64] 
+ wordline_driver 
* No parameters

xwl_driver_65 
+ vdd vss din[65] wl_en wl[65] 
+ wordline_driver 
* No parameters

xwl_driver_66 
+ vdd vss din[66] wl_en wl[66] 
+ wordline_driver 
* No parameters

xwl_driver_67 
+ vdd vss din[67] wl_en wl[67] 
+ wordline_driver 
* No parameters

xwl_driver_68 
+ vdd vss din[68] wl_en wl[68] 
+ wordline_driver 
* No parameters

xwl_driver_69 
+ vdd vss din[69] wl_en wl[69] 
+ wordline_driver 
* No parameters

xwl_driver_70 
+ vdd vss din[70] wl_en wl[70] 
+ wordline_driver 
* No parameters

xwl_driver_71 
+ vdd vss din[71] wl_en wl[71] 
+ wordline_driver 
* No parameters

xwl_driver_72 
+ vdd vss din[72] wl_en wl[72] 
+ wordline_driver 
* No parameters

xwl_driver_73 
+ vdd vss din[73] wl_en wl[73] 
+ wordline_driver 
* No parameters

xwl_driver_74 
+ vdd vss din[74] wl_en wl[74] 
+ wordline_driver 
* No parameters

xwl_driver_75 
+ vdd vss din[75] wl_en wl[75] 
+ wordline_driver 
* No parameters

xwl_driver_76 
+ vdd vss din[76] wl_en wl[76] 
+ wordline_driver 
* No parameters

xwl_driver_77 
+ vdd vss din[77] wl_en wl[77] 
+ wordline_driver 
* No parameters

xwl_driver_78 
+ vdd vss din[78] wl_en wl[78] 
+ wordline_driver 
* No parameters

xwl_driver_79 
+ vdd vss din[79] wl_en wl[79] 
+ wordline_driver 
* No parameters

xwl_driver_80 
+ vdd vss din[80] wl_en wl[80] 
+ wordline_driver 
* No parameters

xwl_driver_81 
+ vdd vss din[81] wl_en wl[81] 
+ wordline_driver 
* No parameters

xwl_driver_82 
+ vdd vss din[82] wl_en wl[82] 
+ wordline_driver 
* No parameters

xwl_driver_83 
+ vdd vss din[83] wl_en wl[83] 
+ wordline_driver 
* No parameters

xwl_driver_84 
+ vdd vss din[84] wl_en wl[84] 
+ wordline_driver 
* No parameters

xwl_driver_85 
+ vdd vss din[85] wl_en wl[85] 
+ wordline_driver 
* No parameters

xwl_driver_86 
+ vdd vss din[86] wl_en wl[86] 
+ wordline_driver 
* No parameters

xwl_driver_87 
+ vdd vss din[87] wl_en wl[87] 
+ wordline_driver 
* No parameters

xwl_driver_88 
+ vdd vss din[88] wl_en wl[88] 
+ wordline_driver 
* No parameters

xwl_driver_89 
+ vdd vss din[89] wl_en wl[89] 
+ wordline_driver 
* No parameters

xwl_driver_90 
+ vdd vss din[90] wl_en wl[90] 
+ wordline_driver 
* No parameters

xwl_driver_91 
+ vdd vss din[91] wl_en wl[91] 
+ wordline_driver 
* No parameters

xwl_driver_92 
+ vdd vss din[92] wl_en wl[92] 
+ wordline_driver 
* No parameters

xwl_driver_93 
+ vdd vss din[93] wl_en wl[93] 
+ wordline_driver 
* No parameters

xwl_driver_94 
+ vdd vss din[94] wl_en wl[94] 
+ wordline_driver 
* No parameters

xwl_driver_95 
+ vdd vss din[95] wl_en wl[95] 
+ wordline_driver 
* No parameters

xwl_driver_96 
+ vdd vss din[96] wl_en wl[96] 
+ wordline_driver 
* No parameters

xwl_driver_97 
+ vdd vss din[97] wl_en wl[97] 
+ wordline_driver 
* No parameters

xwl_driver_98 
+ vdd vss din[98] wl_en wl[98] 
+ wordline_driver 
* No parameters

xwl_driver_99 
+ vdd vss din[99] wl_en wl[99] 
+ wordline_driver 
* No parameters

xwl_driver_100 
+ vdd vss din[100] wl_en wl[100] 
+ wordline_driver 
* No parameters

xwl_driver_101 
+ vdd vss din[101] wl_en wl[101] 
+ wordline_driver 
* No parameters

xwl_driver_102 
+ vdd vss din[102] wl_en wl[102] 
+ wordline_driver 
* No parameters

xwl_driver_103 
+ vdd vss din[103] wl_en wl[103] 
+ wordline_driver 
* No parameters

xwl_driver_104 
+ vdd vss din[104] wl_en wl[104] 
+ wordline_driver 
* No parameters

xwl_driver_105 
+ vdd vss din[105] wl_en wl[105] 
+ wordline_driver 
* No parameters

xwl_driver_106 
+ vdd vss din[106] wl_en wl[106] 
+ wordline_driver 
* No parameters

xwl_driver_107 
+ vdd vss din[107] wl_en wl[107] 
+ wordline_driver 
* No parameters

xwl_driver_108 
+ vdd vss din[108] wl_en wl[108] 
+ wordline_driver 
* No parameters

xwl_driver_109 
+ vdd vss din[109] wl_en wl[109] 
+ wordline_driver 
* No parameters

xwl_driver_110 
+ vdd vss din[110] wl_en wl[110] 
+ wordline_driver 
* No parameters

xwl_driver_111 
+ vdd vss din[111] wl_en wl[111] 
+ wordline_driver 
* No parameters

xwl_driver_112 
+ vdd vss din[112] wl_en wl[112] 
+ wordline_driver 
* No parameters

xwl_driver_113 
+ vdd vss din[113] wl_en wl[113] 
+ wordline_driver 
* No parameters

xwl_driver_114 
+ vdd vss din[114] wl_en wl[114] 
+ wordline_driver 
* No parameters

xwl_driver_115 
+ vdd vss din[115] wl_en wl[115] 
+ wordline_driver 
* No parameters

xwl_driver_116 
+ vdd vss din[116] wl_en wl[116] 
+ wordline_driver 
* No parameters

xwl_driver_117 
+ vdd vss din[117] wl_en wl[117] 
+ wordline_driver 
* No parameters

xwl_driver_118 
+ vdd vss din[118] wl_en wl[118] 
+ wordline_driver 
* No parameters

xwl_driver_119 
+ vdd vss din[119] wl_en wl[119] 
+ wordline_driver 
* No parameters

xwl_driver_120 
+ vdd vss din[120] wl_en wl[120] 
+ wordline_driver 
* No parameters

xwl_driver_121 
+ vdd vss din[121] wl_en wl[121] 
+ wordline_driver 
* No parameters

xwl_driver_122 
+ vdd vss din[122] wl_en wl[122] 
+ wordline_driver 
* No parameters

xwl_driver_123 
+ vdd vss din[123] wl_en wl[123] 
+ wordline_driver 
* No parameters

xwl_driver_124 
+ vdd vss din[124] wl_en wl[124] 
+ wordline_driver 
* No parameters

xwl_driver_125 
+ vdd vss din[125] wl_en wl[125] 
+ wordline_driver 
* No parameters

xwl_driver_126 
+ vdd vss din[126] wl_en wl[126] 
+ wordline_driver 
* No parameters

xwl_driver_127 
+ vdd vss din[127] wl_en wl[127] 
+ wordline_driver 
* No parameters

.ENDS

.SUBCKT bitcell_array 
+ vdd vss bl[255] bl[254] bl[253] bl[252] bl[251] bl[250] bl[249] bl[248] bl[247] bl[246] bl[245] bl[244] bl[243] bl[242] bl[241] bl[240] bl[239] bl[238] bl[237] bl[236] bl[235] bl[234] bl[233] bl[232] bl[231] bl[230] bl[229] bl[228] bl[227] bl[226] bl[225] bl[224] bl[223] bl[222] bl[221] bl[220] bl[219] bl[218] bl[217] bl[216] bl[215] bl[214] bl[213] bl[212] bl[211] bl[210] bl[209] bl[208] bl[207] bl[206] bl[205] bl[204] bl[203] bl[202] bl[201] bl[200] bl[199] bl[198] bl[197] bl[196] bl[195] bl[194] bl[193] bl[192] bl[191] bl[190] bl[189] bl[188] bl[187] bl[186] bl[185] bl[184] bl[183] bl[182] bl[181] bl[180] bl[179] bl[178] bl[177] bl[176] bl[175] bl[174] bl[173] bl[172] bl[171] bl[170] bl[169] bl[168] bl[167] bl[166] bl[165] bl[164] bl[163] bl[162] bl[161] bl[160] bl[159] bl[158] bl[157] bl[156] bl[155] bl[154] bl[153] bl[152] bl[151] bl[150] bl[149] bl[148] bl[147] bl[146] bl[145] bl[144] bl[143] bl[142] bl[141] bl[140] bl[139] bl[138] bl[137] bl[136] bl[135] bl[134] bl[133] bl[132] bl[131] bl[130] bl[129] bl[128] bl[127] bl[126] bl[125] bl[124] bl[123] bl[122] bl[121] bl[120] bl[119] bl[118] bl[117] bl[116] bl[115] bl[114] bl[113] bl[112] bl[111] bl[110] bl[109] bl[108] bl[107] bl[106] bl[105] bl[104] bl[103] bl[102] bl[101] bl[100] bl[99] bl[98] bl[97] bl[96] bl[95] bl[94] bl[93] bl[92] bl[91] bl[90] bl[89] bl[88] bl[87] bl[86] bl[85] bl[84] bl[83] bl[82] bl[81] bl[80] bl[79] bl[78] bl[77] bl[76] bl[75] bl[74] bl[73] bl[72] bl[71] bl[70] bl[69] bl[68] bl[67] bl[66] bl[65] bl[64] bl[63] bl[62] bl[61] bl[60] bl[59] bl[58] bl[57] bl[56] bl[55] bl[54] bl[53] bl[52] bl[51] bl[50] bl[49] bl[48] bl[47] bl[46] bl[45] bl[44] bl[43] bl[42] bl[41] bl[40] bl[39] bl[38] bl[37] bl[36] bl[35] bl[34] bl[33] bl[32] bl[31] bl[30] bl[29] bl[28] bl[27] bl[26] bl[25] bl[24] bl[23] bl[22] bl[21] bl[20] bl[19] bl[18] bl[17] bl[16] bl[15] bl[14] bl[13] bl[12] bl[11] bl[10] bl[9] bl[8] bl[7] bl[6] bl[5] bl[4] bl[3] bl[2] bl[1] bl[0] br[255] br[254] br[253] br[252] br[251] br[250] br[249] br[248] br[247] br[246] br[245] br[244] br[243] br[242] br[241] br[240] br[239] br[238] br[237] br[236] br[235] br[234] br[233] br[232] br[231] br[230] br[229] br[228] br[227] br[226] br[225] br[224] br[223] br[222] br[221] br[220] br[219] br[218] br[217] br[216] br[215] br[214] br[213] br[212] br[211] br[210] br[209] br[208] br[207] br[206] br[205] br[204] br[203] br[202] br[201] br[200] br[199] br[198] br[197] br[196] br[195] br[194] br[193] br[192] br[191] br[190] br[189] br[188] br[187] br[186] br[185] br[184] br[183] br[182] br[181] br[180] br[179] br[178] br[177] br[176] br[175] br[174] br[173] br[172] br[171] br[170] br[169] br[168] br[167] br[166] br[165] br[164] br[163] br[162] br[161] br[160] br[159] br[158] br[157] br[156] br[155] br[154] br[153] br[152] br[151] br[150] br[149] br[148] br[147] br[146] br[145] br[144] br[143] br[142] br[141] br[140] br[139] br[138] br[137] br[136] br[135] br[134] br[133] br[132] br[131] br[130] br[129] br[128] br[127] br[126] br[125] br[124] br[123] br[122] br[121] br[120] br[119] br[118] br[117] br[116] br[115] br[114] br[113] br[112] br[111] br[110] br[109] br[108] br[107] br[106] br[105] br[104] br[103] br[102] br[101] br[100] br[99] br[98] br[97] br[96] br[95] br[94] br[93] br[92] br[91] br[90] br[89] br[88] br[87] br[86] br[85] br[84] br[83] br[82] br[81] br[80] br[79] br[78] br[77] br[76] br[75] br[74] br[73] br[72] br[71] br[70] br[69] br[68] br[67] br[66] br[65] br[64] br[63] br[62] br[61] br[60] br[59] br[58] br[57] br[56] br[55] br[54] br[53] br[52] br[51] br[50] br[49] br[48] br[47] br[46] br[45] br[44] br[43] br[42] br[41] br[40] br[39] br[38] br[37] br[36] br[35] br[34] br[33] br[32] br[31] br[30] br[29] br[28] br[27] br[26] br[25] br[24] br[23] br[22] br[21] br[20] br[19] br[18] br[17] br[16] br[15] br[14] br[13] br[12] br[11] br[10] br[9] br[8] br[7] br[6] br[5] br[4] br[3] br[2] br[1] br[0] wl[127] wl[126] wl[125] wl[124] wl[123] wl[122] wl[121] wl[120] wl[119] wl[118] wl[117] wl[116] wl[115] wl[114] wl[113] wl[112] wl[111] wl[110] wl[109] wl[108] wl[107] wl[106] wl[105] wl[104] wl[103] wl[102] wl[101] wl[100] wl[99] wl[98] wl[97] wl[96] wl[95] wl[94] wl[93] wl[92] wl[91] wl[90] wl[89] wl[88] wl[87] wl[86] wl[85] wl[84] wl[83] wl[82] wl[81] wl[80] wl[79] wl[78] wl[77] wl[76] wl[75] wl[74] wl[73] wl[72] wl[71] wl[70] wl[69] wl[68] wl[67] wl[66] wl[65] wl[64] wl[63] wl[62] wl[61] wl[60] wl[59] wl[58] wl[57] wl[56] wl[55] wl[54] wl[53] wl[52] wl[51] wl[50] wl[49] wl[48] wl[47] wl[46] wl[45] wl[44] wl[43] wl[42] wl[41] wl[40] wl[39] wl[38] wl[37] wl[36] wl[35] wl[34] wl[33] wl[32] wl[31] wl[30] wl[29] wl[28] wl[27] wl[26] wl[25] wl[24] wl[23] wl[22] wl[21] wl[20] wl[19] wl[18] wl[17] wl[16] wl[15] wl[14] wl[13] wl[12] wl[11] wl[10] wl[9] wl[8] wl[7] wl[6] wl[5] wl[4] wl[3] wl[2] wl[1] wl[0] vnb vpb rbl rbr 

xbitcell_0_0 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_1 
+ rbl rbr vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_2 
+ bl[0] br[0] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_3 
+ bl[1] br[1] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_4 
+ bl[2] br[2] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_5 
+ bl[3] br[3] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_6 
+ bl[4] br[4] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_7 
+ bl[5] br[5] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_8 
+ bl[6] br[6] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_9 
+ bl[7] br[7] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_10 
+ bl[8] br[8] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_11 
+ bl[9] br[9] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_12 
+ bl[10] br[10] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_13 
+ bl[11] br[11] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_14 
+ bl[12] br[12] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_15 
+ bl[13] br[13] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_16 
+ bl[14] br[14] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_17 
+ bl[15] br[15] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_18 
+ bl[16] br[16] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_19 
+ bl[17] br[17] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_20 
+ bl[18] br[18] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_21 
+ bl[19] br[19] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_22 
+ bl[20] br[20] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_23 
+ bl[21] br[21] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_24 
+ bl[22] br[22] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_25 
+ bl[23] br[23] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_26 
+ bl[24] br[24] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_27 
+ bl[25] br[25] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_28 
+ bl[26] br[26] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_29 
+ bl[27] br[27] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_30 
+ bl[28] br[28] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_31 
+ bl[29] br[29] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_32 
+ bl[30] br[30] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_33 
+ bl[31] br[31] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_34 
+ bl[32] br[32] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_35 
+ bl[33] br[33] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_36 
+ bl[34] br[34] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_37 
+ bl[35] br[35] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_38 
+ bl[36] br[36] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_39 
+ bl[37] br[37] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_40 
+ bl[38] br[38] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_41 
+ bl[39] br[39] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_42 
+ bl[40] br[40] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_43 
+ bl[41] br[41] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_44 
+ bl[42] br[42] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_45 
+ bl[43] br[43] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_46 
+ bl[44] br[44] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_47 
+ bl[45] br[45] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_48 
+ bl[46] br[46] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_49 
+ bl[47] br[47] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_50 
+ bl[48] br[48] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_51 
+ bl[49] br[49] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_52 
+ bl[50] br[50] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_53 
+ bl[51] br[51] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_54 
+ bl[52] br[52] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_55 
+ bl[53] br[53] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_56 
+ bl[54] br[54] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_57 
+ bl[55] br[55] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_58 
+ bl[56] br[56] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_59 
+ bl[57] br[57] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_60 
+ bl[58] br[58] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_61 
+ bl[59] br[59] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_62 
+ bl[60] br[60] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_63 
+ bl[61] br[61] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_64 
+ bl[62] br[62] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_65 
+ bl[63] br[63] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_66 
+ bl[64] br[64] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_67 
+ bl[65] br[65] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_68 
+ bl[66] br[66] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_69 
+ bl[67] br[67] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_70 
+ bl[68] br[68] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_71 
+ bl[69] br[69] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_72 
+ bl[70] br[70] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_73 
+ bl[71] br[71] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_74 
+ bl[72] br[72] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_75 
+ bl[73] br[73] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_76 
+ bl[74] br[74] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_77 
+ bl[75] br[75] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_78 
+ bl[76] br[76] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_79 
+ bl[77] br[77] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_80 
+ bl[78] br[78] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_81 
+ bl[79] br[79] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_82 
+ bl[80] br[80] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_83 
+ bl[81] br[81] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_84 
+ bl[82] br[82] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_85 
+ bl[83] br[83] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_86 
+ bl[84] br[84] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_87 
+ bl[85] br[85] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_88 
+ bl[86] br[86] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_89 
+ bl[87] br[87] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_90 
+ bl[88] br[88] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_91 
+ bl[89] br[89] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_92 
+ bl[90] br[90] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_93 
+ bl[91] br[91] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_94 
+ bl[92] br[92] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_95 
+ bl[93] br[93] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_96 
+ bl[94] br[94] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_97 
+ bl[95] br[95] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_98 
+ bl[96] br[96] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_99 
+ bl[97] br[97] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_100 
+ bl[98] br[98] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_101 
+ bl[99] br[99] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_102 
+ bl[100] br[100] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_103 
+ bl[101] br[101] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_104 
+ bl[102] br[102] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_105 
+ bl[103] br[103] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_106 
+ bl[104] br[104] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_107 
+ bl[105] br[105] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_108 
+ bl[106] br[106] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_109 
+ bl[107] br[107] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_110 
+ bl[108] br[108] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_111 
+ bl[109] br[109] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_112 
+ bl[110] br[110] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_113 
+ bl[111] br[111] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_114 
+ bl[112] br[112] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_115 
+ bl[113] br[113] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_116 
+ bl[114] br[114] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_117 
+ bl[115] br[115] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_118 
+ bl[116] br[116] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_119 
+ bl[117] br[117] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_120 
+ bl[118] br[118] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_121 
+ bl[119] br[119] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_122 
+ bl[120] br[120] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_123 
+ bl[121] br[121] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_124 
+ bl[122] br[122] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_125 
+ bl[123] br[123] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_126 
+ bl[124] br[124] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_127 
+ bl[125] br[125] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_128 
+ bl[126] br[126] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_129 
+ bl[127] br[127] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_130 
+ bl[128] br[128] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_131 
+ bl[129] br[129] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_132 
+ bl[130] br[130] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_133 
+ bl[131] br[131] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_134 
+ bl[132] br[132] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_135 
+ bl[133] br[133] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_136 
+ bl[134] br[134] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_137 
+ bl[135] br[135] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_138 
+ bl[136] br[136] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_139 
+ bl[137] br[137] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_140 
+ bl[138] br[138] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_141 
+ bl[139] br[139] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_142 
+ bl[140] br[140] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_143 
+ bl[141] br[141] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_144 
+ bl[142] br[142] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_145 
+ bl[143] br[143] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_146 
+ bl[144] br[144] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_147 
+ bl[145] br[145] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_148 
+ bl[146] br[146] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_149 
+ bl[147] br[147] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_150 
+ bl[148] br[148] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_151 
+ bl[149] br[149] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_152 
+ bl[150] br[150] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_153 
+ bl[151] br[151] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_154 
+ bl[152] br[152] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_155 
+ bl[153] br[153] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_156 
+ bl[154] br[154] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_157 
+ bl[155] br[155] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_158 
+ bl[156] br[156] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_159 
+ bl[157] br[157] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_160 
+ bl[158] br[158] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_161 
+ bl[159] br[159] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_162 
+ bl[160] br[160] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_163 
+ bl[161] br[161] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_164 
+ bl[162] br[162] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_165 
+ bl[163] br[163] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_166 
+ bl[164] br[164] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_167 
+ bl[165] br[165] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_168 
+ bl[166] br[166] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_169 
+ bl[167] br[167] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_170 
+ bl[168] br[168] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_171 
+ bl[169] br[169] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_172 
+ bl[170] br[170] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_173 
+ bl[171] br[171] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_174 
+ bl[172] br[172] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_175 
+ bl[173] br[173] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_176 
+ bl[174] br[174] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_177 
+ bl[175] br[175] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_178 
+ bl[176] br[176] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_179 
+ bl[177] br[177] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_180 
+ bl[178] br[178] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_181 
+ bl[179] br[179] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_182 
+ bl[180] br[180] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_183 
+ bl[181] br[181] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_184 
+ bl[182] br[182] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_185 
+ bl[183] br[183] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_186 
+ bl[184] br[184] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_187 
+ bl[185] br[185] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_188 
+ bl[186] br[186] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_189 
+ bl[187] br[187] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_190 
+ bl[188] br[188] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_191 
+ bl[189] br[189] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_192 
+ bl[190] br[190] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_193 
+ bl[191] br[191] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_194 
+ bl[192] br[192] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_195 
+ bl[193] br[193] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_196 
+ bl[194] br[194] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_197 
+ bl[195] br[195] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_198 
+ bl[196] br[196] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_199 
+ bl[197] br[197] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_200 
+ bl[198] br[198] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_201 
+ bl[199] br[199] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_202 
+ bl[200] br[200] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_203 
+ bl[201] br[201] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_204 
+ bl[202] br[202] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_205 
+ bl[203] br[203] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_206 
+ bl[204] br[204] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_207 
+ bl[205] br[205] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_208 
+ bl[206] br[206] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_209 
+ bl[207] br[207] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_210 
+ bl[208] br[208] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_211 
+ bl[209] br[209] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_212 
+ bl[210] br[210] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_213 
+ bl[211] br[211] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_214 
+ bl[212] br[212] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_215 
+ bl[213] br[213] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_216 
+ bl[214] br[214] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_217 
+ bl[215] br[215] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_218 
+ bl[216] br[216] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_219 
+ bl[217] br[217] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_220 
+ bl[218] br[218] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_221 
+ bl[219] br[219] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_222 
+ bl[220] br[220] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_223 
+ bl[221] br[221] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_224 
+ bl[222] br[222] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_225 
+ bl[223] br[223] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_226 
+ bl[224] br[224] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_227 
+ bl[225] br[225] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_228 
+ bl[226] br[226] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_229 
+ bl[227] br[227] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_230 
+ bl[228] br[228] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_231 
+ bl[229] br[229] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_232 
+ bl[230] br[230] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_233 
+ bl[231] br[231] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_234 
+ bl[232] br[232] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_235 
+ bl[233] br[233] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_236 
+ bl[234] br[234] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_237 
+ bl[235] br[235] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_238 
+ bl[236] br[236] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_239 
+ bl[237] br[237] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_240 
+ bl[238] br[238] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_241 
+ bl[239] br[239] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_242 
+ bl[240] br[240] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_243 
+ bl[241] br[241] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_244 
+ bl[242] br[242] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_245 
+ bl[243] br[243] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_246 
+ bl[244] br[244] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_247 
+ bl[245] br[245] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_248 
+ bl[246] br[246] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_249 
+ bl[247] br[247] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_250 
+ bl[248] br[248] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_251 
+ bl[249] br[249] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_252 
+ bl[250] br[250] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_253 
+ bl[251] br[251] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_254 
+ bl[252] br[252] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_255 
+ bl[253] br[253] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_256 
+ bl[254] br[254] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_257 
+ bl[255] br[255] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_258 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_259 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_0 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_1 
+ rbl rbr vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_2 
+ bl[0] br[0] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_3 
+ bl[1] br[1] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_4 
+ bl[2] br[2] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_5 
+ bl[3] br[3] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_6 
+ bl[4] br[4] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_7 
+ bl[5] br[5] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_8 
+ bl[6] br[6] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_9 
+ bl[7] br[7] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_10 
+ bl[8] br[8] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_11 
+ bl[9] br[9] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_12 
+ bl[10] br[10] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_13 
+ bl[11] br[11] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_14 
+ bl[12] br[12] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_15 
+ bl[13] br[13] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_16 
+ bl[14] br[14] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_17 
+ bl[15] br[15] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_18 
+ bl[16] br[16] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_19 
+ bl[17] br[17] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_20 
+ bl[18] br[18] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_21 
+ bl[19] br[19] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_22 
+ bl[20] br[20] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_23 
+ bl[21] br[21] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_24 
+ bl[22] br[22] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_25 
+ bl[23] br[23] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_26 
+ bl[24] br[24] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_27 
+ bl[25] br[25] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_28 
+ bl[26] br[26] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_29 
+ bl[27] br[27] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_30 
+ bl[28] br[28] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_31 
+ bl[29] br[29] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_32 
+ bl[30] br[30] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_33 
+ bl[31] br[31] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_34 
+ bl[32] br[32] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_35 
+ bl[33] br[33] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_36 
+ bl[34] br[34] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_37 
+ bl[35] br[35] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_38 
+ bl[36] br[36] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_39 
+ bl[37] br[37] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_40 
+ bl[38] br[38] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_41 
+ bl[39] br[39] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_42 
+ bl[40] br[40] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_43 
+ bl[41] br[41] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_44 
+ bl[42] br[42] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_45 
+ bl[43] br[43] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_46 
+ bl[44] br[44] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_47 
+ bl[45] br[45] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_48 
+ bl[46] br[46] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_49 
+ bl[47] br[47] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_50 
+ bl[48] br[48] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_51 
+ bl[49] br[49] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_52 
+ bl[50] br[50] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_53 
+ bl[51] br[51] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_54 
+ bl[52] br[52] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_55 
+ bl[53] br[53] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_56 
+ bl[54] br[54] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_57 
+ bl[55] br[55] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_58 
+ bl[56] br[56] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_59 
+ bl[57] br[57] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_60 
+ bl[58] br[58] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_61 
+ bl[59] br[59] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_62 
+ bl[60] br[60] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_63 
+ bl[61] br[61] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_64 
+ bl[62] br[62] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_65 
+ bl[63] br[63] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_66 
+ bl[64] br[64] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_67 
+ bl[65] br[65] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_68 
+ bl[66] br[66] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_69 
+ bl[67] br[67] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_70 
+ bl[68] br[68] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_71 
+ bl[69] br[69] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_72 
+ bl[70] br[70] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_73 
+ bl[71] br[71] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_74 
+ bl[72] br[72] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_75 
+ bl[73] br[73] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_76 
+ bl[74] br[74] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_77 
+ bl[75] br[75] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_78 
+ bl[76] br[76] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_79 
+ bl[77] br[77] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_80 
+ bl[78] br[78] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_81 
+ bl[79] br[79] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_82 
+ bl[80] br[80] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_83 
+ bl[81] br[81] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_84 
+ bl[82] br[82] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_85 
+ bl[83] br[83] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_86 
+ bl[84] br[84] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_87 
+ bl[85] br[85] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_88 
+ bl[86] br[86] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_89 
+ bl[87] br[87] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_90 
+ bl[88] br[88] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_91 
+ bl[89] br[89] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_92 
+ bl[90] br[90] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_93 
+ bl[91] br[91] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_94 
+ bl[92] br[92] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_95 
+ bl[93] br[93] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_96 
+ bl[94] br[94] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_97 
+ bl[95] br[95] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_98 
+ bl[96] br[96] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_99 
+ bl[97] br[97] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_100 
+ bl[98] br[98] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_101 
+ bl[99] br[99] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_102 
+ bl[100] br[100] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_103 
+ bl[101] br[101] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_104 
+ bl[102] br[102] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_105 
+ bl[103] br[103] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_106 
+ bl[104] br[104] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_107 
+ bl[105] br[105] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_108 
+ bl[106] br[106] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_109 
+ bl[107] br[107] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_110 
+ bl[108] br[108] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_111 
+ bl[109] br[109] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_112 
+ bl[110] br[110] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_113 
+ bl[111] br[111] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_114 
+ bl[112] br[112] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_115 
+ bl[113] br[113] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_116 
+ bl[114] br[114] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_117 
+ bl[115] br[115] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_118 
+ bl[116] br[116] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_119 
+ bl[117] br[117] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_120 
+ bl[118] br[118] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_121 
+ bl[119] br[119] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_122 
+ bl[120] br[120] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_123 
+ bl[121] br[121] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_124 
+ bl[122] br[122] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_125 
+ bl[123] br[123] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_126 
+ bl[124] br[124] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_127 
+ bl[125] br[125] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_128 
+ bl[126] br[126] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_129 
+ bl[127] br[127] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_130 
+ bl[128] br[128] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_131 
+ bl[129] br[129] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_132 
+ bl[130] br[130] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_133 
+ bl[131] br[131] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_134 
+ bl[132] br[132] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_135 
+ bl[133] br[133] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_136 
+ bl[134] br[134] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_137 
+ bl[135] br[135] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_138 
+ bl[136] br[136] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_139 
+ bl[137] br[137] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_140 
+ bl[138] br[138] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_141 
+ bl[139] br[139] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_142 
+ bl[140] br[140] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_143 
+ bl[141] br[141] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_144 
+ bl[142] br[142] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_145 
+ bl[143] br[143] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_146 
+ bl[144] br[144] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_147 
+ bl[145] br[145] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_148 
+ bl[146] br[146] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_149 
+ bl[147] br[147] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_150 
+ bl[148] br[148] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_151 
+ bl[149] br[149] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_152 
+ bl[150] br[150] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_153 
+ bl[151] br[151] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_154 
+ bl[152] br[152] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_155 
+ bl[153] br[153] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_156 
+ bl[154] br[154] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_157 
+ bl[155] br[155] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_158 
+ bl[156] br[156] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_159 
+ bl[157] br[157] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_160 
+ bl[158] br[158] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_161 
+ bl[159] br[159] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_162 
+ bl[160] br[160] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_163 
+ bl[161] br[161] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_164 
+ bl[162] br[162] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_165 
+ bl[163] br[163] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_166 
+ bl[164] br[164] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_167 
+ bl[165] br[165] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_168 
+ bl[166] br[166] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_169 
+ bl[167] br[167] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_170 
+ bl[168] br[168] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_171 
+ bl[169] br[169] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_172 
+ bl[170] br[170] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_173 
+ bl[171] br[171] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_174 
+ bl[172] br[172] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_175 
+ bl[173] br[173] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_176 
+ bl[174] br[174] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_177 
+ bl[175] br[175] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_178 
+ bl[176] br[176] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_179 
+ bl[177] br[177] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_180 
+ bl[178] br[178] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_181 
+ bl[179] br[179] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_182 
+ bl[180] br[180] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_183 
+ bl[181] br[181] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_184 
+ bl[182] br[182] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_185 
+ bl[183] br[183] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_186 
+ bl[184] br[184] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_187 
+ bl[185] br[185] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_188 
+ bl[186] br[186] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_189 
+ bl[187] br[187] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_190 
+ bl[188] br[188] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_191 
+ bl[189] br[189] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_192 
+ bl[190] br[190] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_193 
+ bl[191] br[191] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_194 
+ bl[192] br[192] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_195 
+ bl[193] br[193] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_196 
+ bl[194] br[194] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_197 
+ bl[195] br[195] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_198 
+ bl[196] br[196] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_199 
+ bl[197] br[197] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_200 
+ bl[198] br[198] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_201 
+ bl[199] br[199] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_202 
+ bl[200] br[200] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_203 
+ bl[201] br[201] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_204 
+ bl[202] br[202] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_205 
+ bl[203] br[203] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_206 
+ bl[204] br[204] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_207 
+ bl[205] br[205] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_208 
+ bl[206] br[206] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_209 
+ bl[207] br[207] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_210 
+ bl[208] br[208] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_211 
+ bl[209] br[209] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_212 
+ bl[210] br[210] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_213 
+ bl[211] br[211] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_214 
+ bl[212] br[212] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_215 
+ bl[213] br[213] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_216 
+ bl[214] br[214] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_217 
+ bl[215] br[215] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_218 
+ bl[216] br[216] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_219 
+ bl[217] br[217] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_220 
+ bl[218] br[218] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_221 
+ bl[219] br[219] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_222 
+ bl[220] br[220] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_223 
+ bl[221] br[221] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_224 
+ bl[222] br[222] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_225 
+ bl[223] br[223] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_226 
+ bl[224] br[224] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_227 
+ bl[225] br[225] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_228 
+ bl[226] br[226] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_229 
+ bl[227] br[227] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_230 
+ bl[228] br[228] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_231 
+ bl[229] br[229] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_232 
+ bl[230] br[230] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_233 
+ bl[231] br[231] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_234 
+ bl[232] br[232] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_235 
+ bl[233] br[233] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_236 
+ bl[234] br[234] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_237 
+ bl[235] br[235] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_238 
+ bl[236] br[236] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_239 
+ bl[237] br[237] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_240 
+ bl[238] br[238] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_241 
+ bl[239] br[239] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_242 
+ bl[240] br[240] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_243 
+ bl[241] br[241] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_244 
+ bl[242] br[242] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_245 
+ bl[243] br[243] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_246 
+ bl[244] br[244] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_247 
+ bl[245] br[245] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_248 
+ bl[246] br[246] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_249 
+ bl[247] br[247] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_250 
+ bl[248] br[248] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_251 
+ bl[249] br[249] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_252 
+ bl[250] br[250] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_253 
+ bl[251] br[251] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_254 
+ bl[252] br[252] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_255 
+ bl[253] br[253] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_256 
+ bl[254] br[254] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_257 
+ bl[255] br[255] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_258 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_259 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_0 
+ vdd vdd vss vdd vpb vnb wl[0] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_2_1 
+ rbl rbr vss vdd vpb vnb wl[0] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_2_2 
+ bl[0] br[0] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_3 
+ bl[1] br[1] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_4 
+ bl[2] br[2] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_5 
+ bl[3] br[3] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_6 
+ bl[4] br[4] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_7 
+ bl[5] br[5] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_8 
+ bl[6] br[6] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_9 
+ bl[7] br[7] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_10 
+ bl[8] br[8] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_11 
+ bl[9] br[9] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_12 
+ bl[10] br[10] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_13 
+ bl[11] br[11] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_14 
+ bl[12] br[12] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_15 
+ bl[13] br[13] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_16 
+ bl[14] br[14] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_17 
+ bl[15] br[15] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_18 
+ bl[16] br[16] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_19 
+ bl[17] br[17] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_20 
+ bl[18] br[18] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_21 
+ bl[19] br[19] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_22 
+ bl[20] br[20] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_23 
+ bl[21] br[21] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_24 
+ bl[22] br[22] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_25 
+ bl[23] br[23] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_26 
+ bl[24] br[24] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_27 
+ bl[25] br[25] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_28 
+ bl[26] br[26] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_29 
+ bl[27] br[27] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_30 
+ bl[28] br[28] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_31 
+ bl[29] br[29] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_32 
+ bl[30] br[30] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_33 
+ bl[31] br[31] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_34 
+ bl[32] br[32] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_35 
+ bl[33] br[33] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_36 
+ bl[34] br[34] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_37 
+ bl[35] br[35] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_38 
+ bl[36] br[36] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_39 
+ bl[37] br[37] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_40 
+ bl[38] br[38] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_41 
+ bl[39] br[39] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_42 
+ bl[40] br[40] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_43 
+ bl[41] br[41] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_44 
+ bl[42] br[42] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_45 
+ bl[43] br[43] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_46 
+ bl[44] br[44] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_47 
+ bl[45] br[45] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_48 
+ bl[46] br[46] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_49 
+ bl[47] br[47] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_50 
+ bl[48] br[48] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_51 
+ bl[49] br[49] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_52 
+ bl[50] br[50] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_53 
+ bl[51] br[51] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_54 
+ bl[52] br[52] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_55 
+ bl[53] br[53] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_56 
+ bl[54] br[54] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_57 
+ bl[55] br[55] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_58 
+ bl[56] br[56] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_59 
+ bl[57] br[57] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_60 
+ bl[58] br[58] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_61 
+ bl[59] br[59] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_62 
+ bl[60] br[60] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_63 
+ bl[61] br[61] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_64 
+ bl[62] br[62] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_65 
+ bl[63] br[63] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_66 
+ bl[64] br[64] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_67 
+ bl[65] br[65] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_68 
+ bl[66] br[66] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_69 
+ bl[67] br[67] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_70 
+ bl[68] br[68] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_71 
+ bl[69] br[69] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_72 
+ bl[70] br[70] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_73 
+ bl[71] br[71] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_74 
+ bl[72] br[72] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_75 
+ bl[73] br[73] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_76 
+ bl[74] br[74] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_77 
+ bl[75] br[75] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_78 
+ bl[76] br[76] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_79 
+ bl[77] br[77] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_80 
+ bl[78] br[78] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_81 
+ bl[79] br[79] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_82 
+ bl[80] br[80] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_83 
+ bl[81] br[81] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_84 
+ bl[82] br[82] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_85 
+ bl[83] br[83] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_86 
+ bl[84] br[84] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_87 
+ bl[85] br[85] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_88 
+ bl[86] br[86] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_89 
+ bl[87] br[87] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_90 
+ bl[88] br[88] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_91 
+ bl[89] br[89] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_92 
+ bl[90] br[90] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_93 
+ bl[91] br[91] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_94 
+ bl[92] br[92] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_95 
+ bl[93] br[93] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_96 
+ bl[94] br[94] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_97 
+ bl[95] br[95] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_98 
+ bl[96] br[96] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_99 
+ bl[97] br[97] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_100 
+ bl[98] br[98] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_101 
+ bl[99] br[99] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_102 
+ bl[100] br[100] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_103 
+ bl[101] br[101] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_104 
+ bl[102] br[102] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_105 
+ bl[103] br[103] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_106 
+ bl[104] br[104] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_107 
+ bl[105] br[105] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_108 
+ bl[106] br[106] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_109 
+ bl[107] br[107] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_110 
+ bl[108] br[108] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_111 
+ bl[109] br[109] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_112 
+ bl[110] br[110] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_113 
+ bl[111] br[111] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_114 
+ bl[112] br[112] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_115 
+ bl[113] br[113] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_116 
+ bl[114] br[114] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_117 
+ bl[115] br[115] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_118 
+ bl[116] br[116] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_119 
+ bl[117] br[117] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_120 
+ bl[118] br[118] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_121 
+ bl[119] br[119] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_122 
+ bl[120] br[120] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_123 
+ bl[121] br[121] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_124 
+ bl[122] br[122] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_125 
+ bl[123] br[123] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_126 
+ bl[124] br[124] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_127 
+ bl[125] br[125] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_128 
+ bl[126] br[126] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_129 
+ bl[127] br[127] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_130 
+ bl[128] br[128] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_131 
+ bl[129] br[129] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_132 
+ bl[130] br[130] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_133 
+ bl[131] br[131] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_134 
+ bl[132] br[132] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_135 
+ bl[133] br[133] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_136 
+ bl[134] br[134] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_137 
+ bl[135] br[135] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_138 
+ bl[136] br[136] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_139 
+ bl[137] br[137] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_140 
+ bl[138] br[138] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_141 
+ bl[139] br[139] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_142 
+ bl[140] br[140] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_143 
+ bl[141] br[141] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_144 
+ bl[142] br[142] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_145 
+ bl[143] br[143] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_146 
+ bl[144] br[144] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_147 
+ bl[145] br[145] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_148 
+ bl[146] br[146] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_149 
+ bl[147] br[147] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_150 
+ bl[148] br[148] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_151 
+ bl[149] br[149] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_152 
+ bl[150] br[150] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_153 
+ bl[151] br[151] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_154 
+ bl[152] br[152] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_155 
+ bl[153] br[153] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_156 
+ bl[154] br[154] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_157 
+ bl[155] br[155] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_158 
+ bl[156] br[156] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_159 
+ bl[157] br[157] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_160 
+ bl[158] br[158] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_161 
+ bl[159] br[159] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_162 
+ bl[160] br[160] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_163 
+ bl[161] br[161] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_164 
+ bl[162] br[162] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_165 
+ bl[163] br[163] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_166 
+ bl[164] br[164] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_167 
+ bl[165] br[165] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_168 
+ bl[166] br[166] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_169 
+ bl[167] br[167] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_170 
+ bl[168] br[168] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_171 
+ bl[169] br[169] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_172 
+ bl[170] br[170] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_173 
+ bl[171] br[171] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_174 
+ bl[172] br[172] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_175 
+ bl[173] br[173] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_176 
+ bl[174] br[174] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_177 
+ bl[175] br[175] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_178 
+ bl[176] br[176] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_179 
+ bl[177] br[177] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_180 
+ bl[178] br[178] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_181 
+ bl[179] br[179] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_182 
+ bl[180] br[180] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_183 
+ bl[181] br[181] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_184 
+ bl[182] br[182] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_185 
+ bl[183] br[183] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_186 
+ bl[184] br[184] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_187 
+ bl[185] br[185] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_188 
+ bl[186] br[186] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_189 
+ bl[187] br[187] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_190 
+ bl[188] br[188] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_191 
+ bl[189] br[189] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_192 
+ bl[190] br[190] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_193 
+ bl[191] br[191] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_194 
+ bl[192] br[192] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_195 
+ bl[193] br[193] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_196 
+ bl[194] br[194] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_197 
+ bl[195] br[195] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_198 
+ bl[196] br[196] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_199 
+ bl[197] br[197] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_200 
+ bl[198] br[198] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_201 
+ bl[199] br[199] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_202 
+ bl[200] br[200] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_203 
+ bl[201] br[201] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_204 
+ bl[202] br[202] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_205 
+ bl[203] br[203] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_206 
+ bl[204] br[204] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_207 
+ bl[205] br[205] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_208 
+ bl[206] br[206] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_209 
+ bl[207] br[207] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_210 
+ bl[208] br[208] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_211 
+ bl[209] br[209] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_212 
+ bl[210] br[210] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_213 
+ bl[211] br[211] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_214 
+ bl[212] br[212] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_215 
+ bl[213] br[213] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_216 
+ bl[214] br[214] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_217 
+ bl[215] br[215] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_218 
+ bl[216] br[216] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_219 
+ bl[217] br[217] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_220 
+ bl[218] br[218] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_221 
+ bl[219] br[219] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_222 
+ bl[220] br[220] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_223 
+ bl[221] br[221] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_224 
+ bl[222] br[222] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_225 
+ bl[223] br[223] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_226 
+ bl[224] br[224] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_227 
+ bl[225] br[225] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_228 
+ bl[226] br[226] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_229 
+ bl[227] br[227] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_230 
+ bl[228] br[228] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_231 
+ bl[229] br[229] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_232 
+ bl[230] br[230] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_233 
+ bl[231] br[231] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_234 
+ bl[232] br[232] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_235 
+ bl[233] br[233] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_236 
+ bl[234] br[234] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_237 
+ bl[235] br[235] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_238 
+ bl[236] br[236] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_239 
+ bl[237] br[237] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_240 
+ bl[238] br[238] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_241 
+ bl[239] br[239] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_242 
+ bl[240] br[240] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_243 
+ bl[241] br[241] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_244 
+ bl[242] br[242] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_245 
+ bl[243] br[243] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_246 
+ bl[244] br[244] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_247 
+ bl[245] br[245] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_248 
+ bl[246] br[246] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_249 
+ bl[247] br[247] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_250 
+ bl[248] br[248] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_251 
+ bl[249] br[249] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_252 
+ bl[250] br[250] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_253 
+ bl[251] br[251] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_254 
+ bl[252] br[252] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_255 
+ bl[253] br[253] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_256 
+ bl[254] br[254] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_257 
+ bl[255] br[255] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_258 
+ vdd vdd vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_259 
+ vdd vdd vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_0 
+ vdd vdd vss vdd vpb vnb wl[1] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_3_1 
+ rbl rbr vss vdd vpb vnb wl[1] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_3_2 
+ bl[0] br[0] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_3 
+ bl[1] br[1] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_4 
+ bl[2] br[2] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_5 
+ bl[3] br[3] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_6 
+ bl[4] br[4] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_7 
+ bl[5] br[5] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_8 
+ bl[6] br[6] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_9 
+ bl[7] br[7] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_10 
+ bl[8] br[8] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_11 
+ bl[9] br[9] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_12 
+ bl[10] br[10] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_13 
+ bl[11] br[11] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_14 
+ bl[12] br[12] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_15 
+ bl[13] br[13] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_16 
+ bl[14] br[14] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_17 
+ bl[15] br[15] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_18 
+ bl[16] br[16] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_19 
+ bl[17] br[17] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_20 
+ bl[18] br[18] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_21 
+ bl[19] br[19] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_22 
+ bl[20] br[20] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_23 
+ bl[21] br[21] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_24 
+ bl[22] br[22] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_25 
+ bl[23] br[23] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_26 
+ bl[24] br[24] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_27 
+ bl[25] br[25] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_28 
+ bl[26] br[26] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_29 
+ bl[27] br[27] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_30 
+ bl[28] br[28] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_31 
+ bl[29] br[29] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_32 
+ bl[30] br[30] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_33 
+ bl[31] br[31] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_34 
+ bl[32] br[32] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_35 
+ bl[33] br[33] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_36 
+ bl[34] br[34] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_37 
+ bl[35] br[35] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_38 
+ bl[36] br[36] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_39 
+ bl[37] br[37] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_40 
+ bl[38] br[38] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_41 
+ bl[39] br[39] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_42 
+ bl[40] br[40] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_43 
+ bl[41] br[41] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_44 
+ bl[42] br[42] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_45 
+ bl[43] br[43] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_46 
+ bl[44] br[44] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_47 
+ bl[45] br[45] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_48 
+ bl[46] br[46] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_49 
+ bl[47] br[47] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_50 
+ bl[48] br[48] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_51 
+ bl[49] br[49] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_52 
+ bl[50] br[50] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_53 
+ bl[51] br[51] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_54 
+ bl[52] br[52] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_55 
+ bl[53] br[53] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_56 
+ bl[54] br[54] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_57 
+ bl[55] br[55] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_58 
+ bl[56] br[56] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_59 
+ bl[57] br[57] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_60 
+ bl[58] br[58] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_61 
+ bl[59] br[59] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_62 
+ bl[60] br[60] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_63 
+ bl[61] br[61] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_64 
+ bl[62] br[62] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_65 
+ bl[63] br[63] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_66 
+ bl[64] br[64] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_67 
+ bl[65] br[65] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_68 
+ bl[66] br[66] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_69 
+ bl[67] br[67] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_70 
+ bl[68] br[68] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_71 
+ bl[69] br[69] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_72 
+ bl[70] br[70] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_73 
+ bl[71] br[71] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_74 
+ bl[72] br[72] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_75 
+ bl[73] br[73] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_76 
+ bl[74] br[74] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_77 
+ bl[75] br[75] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_78 
+ bl[76] br[76] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_79 
+ bl[77] br[77] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_80 
+ bl[78] br[78] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_81 
+ bl[79] br[79] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_82 
+ bl[80] br[80] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_83 
+ bl[81] br[81] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_84 
+ bl[82] br[82] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_85 
+ bl[83] br[83] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_86 
+ bl[84] br[84] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_87 
+ bl[85] br[85] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_88 
+ bl[86] br[86] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_89 
+ bl[87] br[87] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_90 
+ bl[88] br[88] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_91 
+ bl[89] br[89] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_92 
+ bl[90] br[90] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_93 
+ bl[91] br[91] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_94 
+ bl[92] br[92] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_95 
+ bl[93] br[93] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_96 
+ bl[94] br[94] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_97 
+ bl[95] br[95] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_98 
+ bl[96] br[96] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_99 
+ bl[97] br[97] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_100 
+ bl[98] br[98] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_101 
+ bl[99] br[99] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_102 
+ bl[100] br[100] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_103 
+ bl[101] br[101] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_104 
+ bl[102] br[102] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_105 
+ bl[103] br[103] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_106 
+ bl[104] br[104] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_107 
+ bl[105] br[105] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_108 
+ bl[106] br[106] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_109 
+ bl[107] br[107] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_110 
+ bl[108] br[108] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_111 
+ bl[109] br[109] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_112 
+ bl[110] br[110] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_113 
+ bl[111] br[111] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_114 
+ bl[112] br[112] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_115 
+ bl[113] br[113] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_116 
+ bl[114] br[114] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_117 
+ bl[115] br[115] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_118 
+ bl[116] br[116] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_119 
+ bl[117] br[117] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_120 
+ bl[118] br[118] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_121 
+ bl[119] br[119] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_122 
+ bl[120] br[120] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_123 
+ bl[121] br[121] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_124 
+ bl[122] br[122] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_125 
+ bl[123] br[123] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_126 
+ bl[124] br[124] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_127 
+ bl[125] br[125] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_128 
+ bl[126] br[126] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_129 
+ bl[127] br[127] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_130 
+ bl[128] br[128] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_131 
+ bl[129] br[129] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_132 
+ bl[130] br[130] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_133 
+ bl[131] br[131] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_134 
+ bl[132] br[132] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_135 
+ bl[133] br[133] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_136 
+ bl[134] br[134] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_137 
+ bl[135] br[135] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_138 
+ bl[136] br[136] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_139 
+ bl[137] br[137] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_140 
+ bl[138] br[138] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_141 
+ bl[139] br[139] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_142 
+ bl[140] br[140] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_143 
+ bl[141] br[141] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_144 
+ bl[142] br[142] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_145 
+ bl[143] br[143] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_146 
+ bl[144] br[144] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_147 
+ bl[145] br[145] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_148 
+ bl[146] br[146] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_149 
+ bl[147] br[147] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_150 
+ bl[148] br[148] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_151 
+ bl[149] br[149] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_152 
+ bl[150] br[150] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_153 
+ bl[151] br[151] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_154 
+ bl[152] br[152] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_155 
+ bl[153] br[153] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_156 
+ bl[154] br[154] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_157 
+ bl[155] br[155] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_158 
+ bl[156] br[156] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_159 
+ bl[157] br[157] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_160 
+ bl[158] br[158] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_161 
+ bl[159] br[159] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_162 
+ bl[160] br[160] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_163 
+ bl[161] br[161] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_164 
+ bl[162] br[162] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_165 
+ bl[163] br[163] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_166 
+ bl[164] br[164] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_167 
+ bl[165] br[165] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_168 
+ bl[166] br[166] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_169 
+ bl[167] br[167] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_170 
+ bl[168] br[168] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_171 
+ bl[169] br[169] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_172 
+ bl[170] br[170] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_173 
+ bl[171] br[171] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_174 
+ bl[172] br[172] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_175 
+ bl[173] br[173] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_176 
+ bl[174] br[174] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_177 
+ bl[175] br[175] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_178 
+ bl[176] br[176] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_179 
+ bl[177] br[177] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_180 
+ bl[178] br[178] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_181 
+ bl[179] br[179] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_182 
+ bl[180] br[180] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_183 
+ bl[181] br[181] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_184 
+ bl[182] br[182] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_185 
+ bl[183] br[183] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_186 
+ bl[184] br[184] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_187 
+ bl[185] br[185] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_188 
+ bl[186] br[186] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_189 
+ bl[187] br[187] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_190 
+ bl[188] br[188] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_191 
+ bl[189] br[189] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_192 
+ bl[190] br[190] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_193 
+ bl[191] br[191] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_194 
+ bl[192] br[192] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_195 
+ bl[193] br[193] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_196 
+ bl[194] br[194] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_197 
+ bl[195] br[195] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_198 
+ bl[196] br[196] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_199 
+ bl[197] br[197] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_200 
+ bl[198] br[198] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_201 
+ bl[199] br[199] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_202 
+ bl[200] br[200] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_203 
+ bl[201] br[201] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_204 
+ bl[202] br[202] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_205 
+ bl[203] br[203] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_206 
+ bl[204] br[204] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_207 
+ bl[205] br[205] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_208 
+ bl[206] br[206] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_209 
+ bl[207] br[207] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_210 
+ bl[208] br[208] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_211 
+ bl[209] br[209] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_212 
+ bl[210] br[210] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_213 
+ bl[211] br[211] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_214 
+ bl[212] br[212] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_215 
+ bl[213] br[213] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_216 
+ bl[214] br[214] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_217 
+ bl[215] br[215] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_218 
+ bl[216] br[216] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_219 
+ bl[217] br[217] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_220 
+ bl[218] br[218] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_221 
+ bl[219] br[219] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_222 
+ bl[220] br[220] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_223 
+ bl[221] br[221] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_224 
+ bl[222] br[222] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_225 
+ bl[223] br[223] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_226 
+ bl[224] br[224] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_227 
+ bl[225] br[225] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_228 
+ bl[226] br[226] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_229 
+ bl[227] br[227] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_230 
+ bl[228] br[228] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_231 
+ bl[229] br[229] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_232 
+ bl[230] br[230] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_233 
+ bl[231] br[231] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_234 
+ bl[232] br[232] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_235 
+ bl[233] br[233] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_236 
+ bl[234] br[234] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_237 
+ bl[235] br[235] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_238 
+ bl[236] br[236] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_239 
+ bl[237] br[237] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_240 
+ bl[238] br[238] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_241 
+ bl[239] br[239] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_242 
+ bl[240] br[240] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_243 
+ bl[241] br[241] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_244 
+ bl[242] br[242] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_245 
+ bl[243] br[243] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_246 
+ bl[244] br[244] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_247 
+ bl[245] br[245] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_248 
+ bl[246] br[246] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_249 
+ bl[247] br[247] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_250 
+ bl[248] br[248] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_251 
+ bl[249] br[249] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_252 
+ bl[250] br[250] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_253 
+ bl[251] br[251] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_254 
+ bl[252] br[252] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_255 
+ bl[253] br[253] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_256 
+ bl[254] br[254] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_257 
+ bl[255] br[255] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_258 
+ vdd vdd vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_259 
+ vdd vdd vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_0 
+ vdd vdd vss vdd vpb vnb wl[2] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_4_1 
+ rbl rbr vss vdd vpb vnb wl[2] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_4_2 
+ bl[0] br[0] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_3 
+ bl[1] br[1] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_4 
+ bl[2] br[2] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_5 
+ bl[3] br[3] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_6 
+ bl[4] br[4] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_7 
+ bl[5] br[5] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_8 
+ bl[6] br[6] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_9 
+ bl[7] br[7] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_10 
+ bl[8] br[8] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_11 
+ bl[9] br[9] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_12 
+ bl[10] br[10] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_13 
+ bl[11] br[11] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_14 
+ bl[12] br[12] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_15 
+ bl[13] br[13] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_16 
+ bl[14] br[14] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_17 
+ bl[15] br[15] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_18 
+ bl[16] br[16] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_19 
+ bl[17] br[17] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_20 
+ bl[18] br[18] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_21 
+ bl[19] br[19] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_22 
+ bl[20] br[20] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_23 
+ bl[21] br[21] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_24 
+ bl[22] br[22] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_25 
+ bl[23] br[23] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_26 
+ bl[24] br[24] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_27 
+ bl[25] br[25] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_28 
+ bl[26] br[26] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_29 
+ bl[27] br[27] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_30 
+ bl[28] br[28] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_31 
+ bl[29] br[29] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_32 
+ bl[30] br[30] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_33 
+ bl[31] br[31] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_34 
+ bl[32] br[32] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_35 
+ bl[33] br[33] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_36 
+ bl[34] br[34] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_37 
+ bl[35] br[35] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_38 
+ bl[36] br[36] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_39 
+ bl[37] br[37] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_40 
+ bl[38] br[38] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_41 
+ bl[39] br[39] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_42 
+ bl[40] br[40] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_43 
+ bl[41] br[41] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_44 
+ bl[42] br[42] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_45 
+ bl[43] br[43] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_46 
+ bl[44] br[44] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_47 
+ bl[45] br[45] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_48 
+ bl[46] br[46] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_49 
+ bl[47] br[47] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_50 
+ bl[48] br[48] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_51 
+ bl[49] br[49] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_52 
+ bl[50] br[50] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_53 
+ bl[51] br[51] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_54 
+ bl[52] br[52] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_55 
+ bl[53] br[53] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_56 
+ bl[54] br[54] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_57 
+ bl[55] br[55] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_58 
+ bl[56] br[56] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_59 
+ bl[57] br[57] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_60 
+ bl[58] br[58] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_61 
+ bl[59] br[59] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_62 
+ bl[60] br[60] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_63 
+ bl[61] br[61] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_64 
+ bl[62] br[62] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_65 
+ bl[63] br[63] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_66 
+ bl[64] br[64] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_67 
+ bl[65] br[65] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_68 
+ bl[66] br[66] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_69 
+ bl[67] br[67] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_70 
+ bl[68] br[68] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_71 
+ bl[69] br[69] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_72 
+ bl[70] br[70] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_73 
+ bl[71] br[71] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_74 
+ bl[72] br[72] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_75 
+ bl[73] br[73] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_76 
+ bl[74] br[74] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_77 
+ bl[75] br[75] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_78 
+ bl[76] br[76] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_79 
+ bl[77] br[77] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_80 
+ bl[78] br[78] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_81 
+ bl[79] br[79] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_82 
+ bl[80] br[80] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_83 
+ bl[81] br[81] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_84 
+ bl[82] br[82] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_85 
+ bl[83] br[83] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_86 
+ bl[84] br[84] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_87 
+ bl[85] br[85] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_88 
+ bl[86] br[86] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_89 
+ bl[87] br[87] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_90 
+ bl[88] br[88] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_91 
+ bl[89] br[89] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_92 
+ bl[90] br[90] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_93 
+ bl[91] br[91] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_94 
+ bl[92] br[92] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_95 
+ bl[93] br[93] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_96 
+ bl[94] br[94] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_97 
+ bl[95] br[95] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_98 
+ bl[96] br[96] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_99 
+ bl[97] br[97] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_100 
+ bl[98] br[98] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_101 
+ bl[99] br[99] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_102 
+ bl[100] br[100] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_103 
+ bl[101] br[101] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_104 
+ bl[102] br[102] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_105 
+ bl[103] br[103] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_106 
+ bl[104] br[104] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_107 
+ bl[105] br[105] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_108 
+ bl[106] br[106] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_109 
+ bl[107] br[107] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_110 
+ bl[108] br[108] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_111 
+ bl[109] br[109] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_112 
+ bl[110] br[110] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_113 
+ bl[111] br[111] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_114 
+ bl[112] br[112] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_115 
+ bl[113] br[113] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_116 
+ bl[114] br[114] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_117 
+ bl[115] br[115] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_118 
+ bl[116] br[116] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_119 
+ bl[117] br[117] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_120 
+ bl[118] br[118] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_121 
+ bl[119] br[119] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_122 
+ bl[120] br[120] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_123 
+ bl[121] br[121] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_124 
+ bl[122] br[122] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_125 
+ bl[123] br[123] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_126 
+ bl[124] br[124] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_127 
+ bl[125] br[125] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_128 
+ bl[126] br[126] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_129 
+ bl[127] br[127] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_130 
+ bl[128] br[128] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_131 
+ bl[129] br[129] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_132 
+ bl[130] br[130] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_133 
+ bl[131] br[131] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_134 
+ bl[132] br[132] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_135 
+ bl[133] br[133] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_136 
+ bl[134] br[134] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_137 
+ bl[135] br[135] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_138 
+ bl[136] br[136] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_139 
+ bl[137] br[137] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_140 
+ bl[138] br[138] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_141 
+ bl[139] br[139] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_142 
+ bl[140] br[140] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_143 
+ bl[141] br[141] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_144 
+ bl[142] br[142] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_145 
+ bl[143] br[143] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_146 
+ bl[144] br[144] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_147 
+ bl[145] br[145] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_148 
+ bl[146] br[146] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_149 
+ bl[147] br[147] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_150 
+ bl[148] br[148] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_151 
+ bl[149] br[149] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_152 
+ bl[150] br[150] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_153 
+ bl[151] br[151] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_154 
+ bl[152] br[152] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_155 
+ bl[153] br[153] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_156 
+ bl[154] br[154] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_157 
+ bl[155] br[155] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_158 
+ bl[156] br[156] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_159 
+ bl[157] br[157] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_160 
+ bl[158] br[158] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_161 
+ bl[159] br[159] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_162 
+ bl[160] br[160] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_163 
+ bl[161] br[161] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_164 
+ bl[162] br[162] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_165 
+ bl[163] br[163] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_166 
+ bl[164] br[164] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_167 
+ bl[165] br[165] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_168 
+ bl[166] br[166] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_169 
+ bl[167] br[167] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_170 
+ bl[168] br[168] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_171 
+ bl[169] br[169] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_172 
+ bl[170] br[170] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_173 
+ bl[171] br[171] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_174 
+ bl[172] br[172] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_175 
+ bl[173] br[173] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_176 
+ bl[174] br[174] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_177 
+ bl[175] br[175] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_178 
+ bl[176] br[176] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_179 
+ bl[177] br[177] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_180 
+ bl[178] br[178] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_181 
+ bl[179] br[179] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_182 
+ bl[180] br[180] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_183 
+ bl[181] br[181] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_184 
+ bl[182] br[182] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_185 
+ bl[183] br[183] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_186 
+ bl[184] br[184] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_187 
+ bl[185] br[185] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_188 
+ bl[186] br[186] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_189 
+ bl[187] br[187] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_190 
+ bl[188] br[188] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_191 
+ bl[189] br[189] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_192 
+ bl[190] br[190] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_193 
+ bl[191] br[191] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_194 
+ bl[192] br[192] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_195 
+ bl[193] br[193] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_196 
+ bl[194] br[194] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_197 
+ bl[195] br[195] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_198 
+ bl[196] br[196] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_199 
+ bl[197] br[197] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_200 
+ bl[198] br[198] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_201 
+ bl[199] br[199] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_202 
+ bl[200] br[200] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_203 
+ bl[201] br[201] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_204 
+ bl[202] br[202] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_205 
+ bl[203] br[203] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_206 
+ bl[204] br[204] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_207 
+ bl[205] br[205] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_208 
+ bl[206] br[206] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_209 
+ bl[207] br[207] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_210 
+ bl[208] br[208] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_211 
+ bl[209] br[209] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_212 
+ bl[210] br[210] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_213 
+ bl[211] br[211] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_214 
+ bl[212] br[212] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_215 
+ bl[213] br[213] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_216 
+ bl[214] br[214] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_217 
+ bl[215] br[215] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_218 
+ bl[216] br[216] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_219 
+ bl[217] br[217] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_220 
+ bl[218] br[218] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_221 
+ bl[219] br[219] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_222 
+ bl[220] br[220] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_223 
+ bl[221] br[221] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_224 
+ bl[222] br[222] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_225 
+ bl[223] br[223] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_226 
+ bl[224] br[224] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_227 
+ bl[225] br[225] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_228 
+ bl[226] br[226] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_229 
+ bl[227] br[227] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_230 
+ bl[228] br[228] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_231 
+ bl[229] br[229] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_232 
+ bl[230] br[230] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_233 
+ bl[231] br[231] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_234 
+ bl[232] br[232] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_235 
+ bl[233] br[233] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_236 
+ bl[234] br[234] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_237 
+ bl[235] br[235] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_238 
+ bl[236] br[236] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_239 
+ bl[237] br[237] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_240 
+ bl[238] br[238] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_241 
+ bl[239] br[239] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_242 
+ bl[240] br[240] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_243 
+ bl[241] br[241] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_244 
+ bl[242] br[242] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_245 
+ bl[243] br[243] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_246 
+ bl[244] br[244] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_247 
+ bl[245] br[245] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_248 
+ bl[246] br[246] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_249 
+ bl[247] br[247] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_250 
+ bl[248] br[248] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_251 
+ bl[249] br[249] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_252 
+ bl[250] br[250] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_253 
+ bl[251] br[251] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_254 
+ bl[252] br[252] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_255 
+ bl[253] br[253] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_256 
+ bl[254] br[254] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_257 
+ bl[255] br[255] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_258 
+ vdd vdd vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_259 
+ vdd vdd vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_0 
+ vdd vdd vss vdd vpb vnb wl[3] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_5_1 
+ rbl rbr vss vdd vpb vnb wl[3] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_5_2 
+ bl[0] br[0] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_3 
+ bl[1] br[1] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_4 
+ bl[2] br[2] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_5 
+ bl[3] br[3] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_6 
+ bl[4] br[4] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_7 
+ bl[5] br[5] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_8 
+ bl[6] br[6] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_9 
+ bl[7] br[7] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_10 
+ bl[8] br[8] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_11 
+ bl[9] br[9] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_12 
+ bl[10] br[10] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_13 
+ bl[11] br[11] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_14 
+ bl[12] br[12] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_15 
+ bl[13] br[13] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_16 
+ bl[14] br[14] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_17 
+ bl[15] br[15] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_18 
+ bl[16] br[16] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_19 
+ bl[17] br[17] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_20 
+ bl[18] br[18] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_21 
+ bl[19] br[19] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_22 
+ bl[20] br[20] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_23 
+ bl[21] br[21] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_24 
+ bl[22] br[22] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_25 
+ bl[23] br[23] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_26 
+ bl[24] br[24] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_27 
+ bl[25] br[25] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_28 
+ bl[26] br[26] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_29 
+ bl[27] br[27] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_30 
+ bl[28] br[28] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_31 
+ bl[29] br[29] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_32 
+ bl[30] br[30] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_33 
+ bl[31] br[31] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_34 
+ bl[32] br[32] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_35 
+ bl[33] br[33] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_36 
+ bl[34] br[34] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_37 
+ bl[35] br[35] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_38 
+ bl[36] br[36] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_39 
+ bl[37] br[37] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_40 
+ bl[38] br[38] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_41 
+ bl[39] br[39] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_42 
+ bl[40] br[40] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_43 
+ bl[41] br[41] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_44 
+ bl[42] br[42] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_45 
+ bl[43] br[43] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_46 
+ bl[44] br[44] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_47 
+ bl[45] br[45] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_48 
+ bl[46] br[46] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_49 
+ bl[47] br[47] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_50 
+ bl[48] br[48] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_51 
+ bl[49] br[49] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_52 
+ bl[50] br[50] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_53 
+ bl[51] br[51] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_54 
+ bl[52] br[52] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_55 
+ bl[53] br[53] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_56 
+ bl[54] br[54] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_57 
+ bl[55] br[55] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_58 
+ bl[56] br[56] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_59 
+ bl[57] br[57] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_60 
+ bl[58] br[58] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_61 
+ bl[59] br[59] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_62 
+ bl[60] br[60] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_63 
+ bl[61] br[61] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_64 
+ bl[62] br[62] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_65 
+ bl[63] br[63] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_66 
+ bl[64] br[64] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_67 
+ bl[65] br[65] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_68 
+ bl[66] br[66] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_69 
+ bl[67] br[67] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_70 
+ bl[68] br[68] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_71 
+ bl[69] br[69] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_72 
+ bl[70] br[70] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_73 
+ bl[71] br[71] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_74 
+ bl[72] br[72] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_75 
+ bl[73] br[73] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_76 
+ bl[74] br[74] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_77 
+ bl[75] br[75] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_78 
+ bl[76] br[76] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_79 
+ bl[77] br[77] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_80 
+ bl[78] br[78] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_81 
+ bl[79] br[79] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_82 
+ bl[80] br[80] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_83 
+ bl[81] br[81] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_84 
+ bl[82] br[82] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_85 
+ bl[83] br[83] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_86 
+ bl[84] br[84] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_87 
+ bl[85] br[85] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_88 
+ bl[86] br[86] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_89 
+ bl[87] br[87] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_90 
+ bl[88] br[88] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_91 
+ bl[89] br[89] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_92 
+ bl[90] br[90] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_93 
+ bl[91] br[91] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_94 
+ bl[92] br[92] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_95 
+ bl[93] br[93] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_96 
+ bl[94] br[94] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_97 
+ bl[95] br[95] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_98 
+ bl[96] br[96] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_99 
+ bl[97] br[97] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_100 
+ bl[98] br[98] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_101 
+ bl[99] br[99] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_102 
+ bl[100] br[100] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_103 
+ bl[101] br[101] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_104 
+ bl[102] br[102] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_105 
+ bl[103] br[103] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_106 
+ bl[104] br[104] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_107 
+ bl[105] br[105] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_108 
+ bl[106] br[106] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_109 
+ bl[107] br[107] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_110 
+ bl[108] br[108] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_111 
+ bl[109] br[109] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_112 
+ bl[110] br[110] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_113 
+ bl[111] br[111] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_114 
+ bl[112] br[112] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_115 
+ bl[113] br[113] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_116 
+ bl[114] br[114] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_117 
+ bl[115] br[115] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_118 
+ bl[116] br[116] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_119 
+ bl[117] br[117] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_120 
+ bl[118] br[118] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_121 
+ bl[119] br[119] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_122 
+ bl[120] br[120] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_123 
+ bl[121] br[121] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_124 
+ bl[122] br[122] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_125 
+ bl[123] br[123] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_126 
+ bl[124] br[124] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_127 
+ bl[125] br[125] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_128 
+ bl[126] br[126] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_129 
+ bl[127] br[127] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_130 
+ bl[128] br[128] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_131 
+ bl[129] br[129] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_132 
+ bl[130] br[130] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_133 
+ bl[131] br[131] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_134 
+ bl[132] br[132] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_135 
+ bl[133] br[133] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_136 
+ bl[134] br[134] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_137 
+ bl[135] br[135] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_138 
+ bl[136] br[136] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_139 
+ bl[137] br[137] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_140 
+ bl[138] br[138] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_141 
+ bl[139] br[139] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_142 
+ bl[140] br[140] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_143 
+ bl[141] br[141] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_144 
+ bl[142] br[142] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_145 
+ bl[143] br[143] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_146 
+ bl[144] br[144] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_147 
+ bl[145] br[145] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_148 
+ bl[146] br[146] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_149 
+ bl[147] br[147] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_150 
+ bl[148] br[148] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_151 
+ bl[149] br[149] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_152 
+ bl[150] br[150] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_153 
+ bl[151] br[151] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_154 
+ bl[152] br[152] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_155 
+ bl[153] br[153] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_156 
+ bl[154] br[154] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_157 
+ bl[155] br[155] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_158 
+ bl[156] br[156] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_159 
+ bl[157] br[157] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_160 
+ bl[158] br[158] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_161 
+ bl[159] br[159] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_162 
+ bl[160] br[160] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_163 
+ bl[161] br[161] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_164 
+ bl[162] br[162] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_165 
+ bl[163] br[163] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_166 
+ bl[164] br[164] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_167 
+ bl[165] br[165] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_168 
+ bl[166] br[166] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_169 
+ bl[167] br[167] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_170 
+ bl[168] br[168] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_171 
+ bl[169] br[169] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_172 
+ bl[170] br[170] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_173 
+ bl[171] br[171] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_174 
+ bl[172] br[172] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_175 
+ bl[173] br[173] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_176 
+ bl[174] br[174] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_177 
+ bl[175] br[175] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_178 
+ bl[176] br[176] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_179 
+ bl[177] br[177] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_180 
+ bl[178] br[178] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_181 
+ bl[179] br[179] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_182 
+ bl[180] br[180] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_183 
+ bl[181] br[181] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_184 
+ bl[182] br[182] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_185 
+ bl[183] br[183] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_186 
+ bl[184] br[184] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_187 
+ bl[185] br[185] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_188 
+ bl[186] br[186] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_189 
+ bl[187] br[187] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_190 
+ bl[188] br[188] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_191 
+ bl[189] br[189] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_192 
+ bl[190] br[190] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_193 
+ bl[191] br[191] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_194 
+ bl[192] br[192] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_195 
+ bl[193] br[193] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_196 
+ bl[194] br[194] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_197 
+ bl[195] br[195] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_198 
+ bl[196] br[196] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_199 
+ bl[197] br[197] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_200 
+ bl[198] br[198] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_201 
+ bl[199] br[199] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_202 
+ bl[200] br[200] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_203 
+ bl[201] br[201] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_204 
+ bl[202] br[202] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_205 
+ bl[203] br[203] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_206 
+ bl[204] br[204] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_207 
+ bl[205] br[205] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_208 
+ bl[206] br[206] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_209 
+ bl[207] br[207] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_210 
+ bl[208] br[208] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_211 
+ bl[209] br[209] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_212 
+ bl[210] br[210] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_213 
+ bl[211] br[211] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_214 
+ bl[212] br[212] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_215 
+ bl[213] br[213] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_216 
+ bl[214] br[214] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_217 
+ bl[215] br[215] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_218 
+ bl[216] br[216] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_219 
+ bl[217] br[217] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_220 
+ bl[218] br[218] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_221 
+ bl[219] br[219] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_222 
+ bl[220] br[220] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_223 
+ bl[221] br[221] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_224 
+ bl[222] br[222] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_225 
+ bl[223] br[223] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_226 
+ bl[224] br[224] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_227 
+ bl[225] br[225] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_228 
+ bl[226] br[226] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_229 
+ bl[227] br[227] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_230 
+ bl[228] br[228] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_231 
+ bl[229] br[229] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_232 
+ bl[230] br[230] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_233 
+ bl[231] br[231] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_234 
+ bl[232] br[232] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_235 
+ bl[233] br[233] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_236 
+ bl[234] br[234] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_237 
+ bl[235] br[235] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_238 
+ bl[236] br[236] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_239 
+ bl[237] br[237] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_240 
+ bl[238] br[238] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_241 
+ bl[239] br[239] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_242 
+ bl[240] br[240] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_243 
+ bl[241] br[241] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_244 
+ bl[242] br[242] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_245 
+ bl[243] br[243] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_246 
+ bl[244] br[244] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_247 
+ bl[245] br[245] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_248 
+ bl[246] br[246] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_249 
+ bl[247] br[247] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_250 
+ bl[248] br[248] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_251 
+ bl[249] br[249] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_252 
+ bl[250] br[250] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_253 
+ bl[251] br[251] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_254 
+ bl[252] br[252] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_255 
+ bl[253] br[253] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_256 
+ bl[254] br[254] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_257 
+ bl[255] br[255] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_258 
+ vdd vdd vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_259 
+ vdd vdd vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_0 
+ vdd vdd vss vdd vpb vnb wl[4] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_6_1 
+ rbl rbr vss vdd vpb vnb wl[4] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_6_2 
+ bl[0] br[0] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_3 
+ bl[1] br[1] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_4 
+ bl[2] br[2] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_5 
+ bl[3] br[3] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_6 
+ bl[4] br[4] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_7 
+ bl[5] br[5] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_8 
+ bl[6] br[6] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_9 
+ bl[7] br[7] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_10 
+ bl[8] br[8] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_11 
+ bl[9] br[9] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_12 
+ bl[10] br[10] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_13 
+ bl[11] br[11] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_14 
+ bl[12] br[12] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_15 
+ bl[13] br[13] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_16 
+ bl[14] br[14] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_17 
+ bl[15] br[15] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_18 
+ bl[16] br[16] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_19 
+ bl[17] br[17] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_20 
+ bl[18] br[18] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_21 
+ bl[19] br[19] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_22 
+ bl[20] br[20] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_23 
+ bl[21] br[21] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_24 
+ bl[22] br[22] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_25 
+ bl[23] br[23] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_26 
+ bl[24] br[24] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_27 
+ bl[25] br[25] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_28 
+ bl[26] br[26] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_29 
+ bl[27] br[27] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_30 
+ bl[28] br[28] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_31 
+ bl[29] br[29] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_32 
+ bl[30] br[30] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_33 
+ bl[31] br[31] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_34 
+ bl[32] br[32] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_35 
+ bl[33] br[33] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_36 
+ bl[34] br[34] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_37 
+ bl[35] br[35] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_38 
+ bl[36] br[36] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_39 
+ bl[37] br[37] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_40 
+ bl[38] br[38] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_41 
+ bl[39] br[39] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_42 
+ bl[40] br[40] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_43 
+ bl[41] br[41] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_44 
+ bl[42] br[42] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_45 
+ bl[43] br[43] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_46 
+ bl[44] br[44] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_47 
+ bl[45] br[45] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_48 
+ bl[46] br[46] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_49 
+ bl[47] br[47] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_50 
+ bl[48] br[48] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_51 
+ bl[49] br[49] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_52 
+ bl[50] br[50] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_53 
+ bl[51] br[51] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_54 
+ bl[52] br[52] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_55 
+ bl[53] br[53] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_56 
+ bl[54] br[54] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_57 
+ bl[55] br[55] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_58 
+ bl[56] br[56] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_59 
+ bl[57] br[57] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_60 
+ bl[58] br[58] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_61 
+ bl[59] br[59] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_62 
+ bl[60] br[60] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_63 
+ bl[61] br[61] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_64 
+ bl[62] br[62] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_65 
+ bl[63] br[63] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_66 
+ bl[64] br[64] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_67 
+ bl[65] br[65] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_68 
+ bl[66] br[66] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_69 
+ bl[67] br[67] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_70 
+ bl[68] br[68] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_71 
+ bl[69] br[69] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_72 
+ bl[70] br[70] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_73 
+ bl[71] br[71] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_74 
+ bl[72] br[72] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_75 
+ bl[73] br[73] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_76 
+ bl[74] br[74] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_77 
+ bl[75] br[75] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_78 
+ bl[76] br[76] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_79 
+ bl[77] br[77] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_80 
+ bl[78] br[78] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_81 
+ bl[79] br[79] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_82 
+ bl[80] br[80] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_83 
+ bl[81] br[81] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_84 
+ bl[82] br[82] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_85 
+ bl[83] br[83] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_86 
+ bl[84] br[84] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_87 
+ bl[85] br[85] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_88 
+ bl[86] br[86] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_89 
+ bl[87] br[87] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_90 
+ bl[88] br[88] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_91 
+ bl[89] br[89] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_92 
+ bl[90] br[90] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_93 
+ bl[91] br[91] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_94 
+ bl[92] br[92] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_95 
+ bl[93] br[93] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_96 
+ bl[94] br[94] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_97 
+ bl[95] br[95] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_98 
+ bl[96] br[96] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_99 
+ bl[97] br[97] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_100 
+ bl[98] br[98] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_101 
+ bl[99] br[99] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_102 
+ bl[100] br[100] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_103 
+ bl[101] br[101] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_104 
+ bl[102] br[102] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_105 
+ bl[103] br[103] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_106 
+ bl[104] br[104] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_107 
+ bl[105] br[105] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_108 
+ bl[106] br[106] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_109 
+ bl[107] br[107] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_110 
+ bl[108] br[108] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_111 
+ bl[109] br[109] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_112 
+ bl[110] br[110] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_113 
+ bl[111] br[111] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_114 
+ bl[112] br[112] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_115 
+ bl[113] br[113] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_116 
+ bl[114] br[114] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_117 
+ bl[115] br[115] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_118 
+ bl[116] br[116] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_119 
+ bl[117] br[117] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_120 
+ bl[118] br[118] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_121 
+ bl[119] br[119] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_122 
+ bl[120] br[120] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_123 
+ bl[121] br[121] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_124 
+ bl[122] br[122] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_125 
+ bl[123] br[123] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_126 
+ bl[124] br[124] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_127 
+ bl[125] br[125] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_128 
+ bl[126] br[126] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_129 
+ bl[127] br[127] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_130 
+ bl[128] br[128] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_131 
+ bl[129] br[129] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_132 
+ bl[130] br[130] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_133 
+ bl[131] br[131] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_134 
+ bl[132] br[132] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_135 
+ bl[133] br[133] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_136 
+ bl[134] br[134] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_137 
+ bl[135] br[135] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_138 
+ bl[136] br[136] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_139 
+ bl[137] br[137] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_140 
+ bl[138] br[138] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_141 
+ bl[139] br[139] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_142 
+ bl[140] br[140] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_143 
+ bl[141] br[141] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_144 
+ bl[142] br[142] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_145 
+ bl[143] br[143] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_146 
+ bl[144] br[144] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_147 
+ bl[145] br[145] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_148 
+ bl[146] br[146] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_149 
+ bl[147] br[147] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_150 
+ bl[148] br[148] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_151 
+ bl[149] br[149] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_152 
+ bl[150] br[150] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_153 
+ bl[151] br[151] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_154 
+ bl[152] br[152] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_155 
+ bl[153] br[153] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_156 
+ bl[154] br[154] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_157 
+ bl[155] br[155] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_158 
+ bl[156] br[156] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_159 
+ bl[157] br[157] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_160 
+ bl[158] br[158] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_161 
+ bl[159] br[159] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_162 
+ bl[160] br[160] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_163 
+ bl[161] br[161] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_164 
+ bl[162] br[162] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_165 
+ bl[163] br[163] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_166 
+ bl[164] br[164] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_167 
+ bl[165] br[165] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_168 
+ bl[166] br[166] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_169 
+ bl[167] br[167] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_170 
+ bl[168] br[168] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_171 
+ bl[169] br[169] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_172 
+ bl[170] br[170] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_173 
+ bl[171] br[171] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_174 
+ bl[172] br[172] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_175 
+ bl[173] br[173] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_176 
+ bl[174] br[174] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_177 
+ bl[175] br[175] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_178 
+ bl[176] br[176] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_179 
+ bl[177] br[177] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_180 
+ bl[178] br[178] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_181 
+ bl[179] br[179] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_182 
+ bl[180] br[180] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_183 
+ bl[181] br[181] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_184 
+ bl[182] br[182] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_185 
+ bl[183] br[183] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_186 
+ bl[184] br[184] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_187 
+ bl[185] br[185] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_188 
+ bl[186] br[186] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_189 
+ bl[187] br[187] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_190 
+ bl[188] br[188] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_191 
+ bl[189] br[189] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_192 
+ bl[190] br[190] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_193 
+ bl[191] br[191] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_194 
+ bl[192] br[192] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_195 
+ bl[193] br[193] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_196 
+ bl[194] br[194] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_197 
+ bl[195] br[195] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_198 
+ bl[196] br[196] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_199 
+ bl[197] br[197] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_200 
+ bl[198] br[198] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_201 
+ bl[199] br[199] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_202 
+ bl[200] br[200] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_203 
+ bl[201] br[201] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_204 
+ bl[202] br[202] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_205 
+ bl[203] br[203] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_206 
+ bl[204] br[204] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_207 
+ bl[205] br[205] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_208 
+ bl[206] br[206] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_209 
+ bl[207] br[207] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_210 
+ bl[208] br[208] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_211 
+ bl[209] br[209] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_212 
+ bl[210] br[210] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_213 
+ bl[211] br[211] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_214 
+ bl[212] br[212] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_215 
+ bl[213] br[213] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_216 
+ bl[214] br[214] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_217 
+ bl[215] br[215] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_218 
+ bl[216] br[216] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_219 
+ bl[217] br[217] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_220 
+ bl[218] br[218] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_221 
+ bl[219] br[219] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_222 
+ bl[220] br[220] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_223 
+ bl[221] br[221] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_224 
+ bl[222] br[222] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_225 
+ bl[223] br[223] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_226 
+ bl[224] br[224] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_227 
+ bl[225] br[225] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_228 
+ bl[226] br[226] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_229 
+ bl[227] br[227] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_230 
+ bl[228] br[228] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_231 
+ bl[229] br[229] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_232 
+ bl[230] br[230] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_233 
+ bl[231] br[231] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_234 
+ bl[232] br[232] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_235 
+ bl[233] br[233] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_236 
+ bl[234] br[234] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_237 
+ bl[235] br[235] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_238 
+ bl[236] br[236] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_239 
+ bl[237] br[237] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_240 
+ bl[238] br[238] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_241 
+ bl[239] br[239] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_242 
+ bl[240] br[240] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_243 
+ bl[241] br[241] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_244 
+ bl[242] br[242] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_245 
+ bl[243] br[243] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_246 
+ bl[244] br[244] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_247 
+ bl[245] br[245] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_248 
+ bl[246] br[246] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_249 
+ bl[247] br[247] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_250 
+ bl[248] br[248] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_251 
+ bl[249] br[249] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_252 
+ bl[250] br[250] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_253 
+ bl[251] br[251] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_254 
+ bl[252] br[252] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_255 
+ bl[253] br[253] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_256 
+ bl[254] br[254] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_257 
+ bl[255] br[255] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_258 
+ vdd vdd vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_259 
+ vdd vdd vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_0 
+ vdd vdd vss vdd vpb vnb wl[5] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_7_1 
+ rbl rbr vss vdd vpb vnb wl[5] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_7_2 
+ bl[0] br[0] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_3 
+ bl[1] br[1] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_4 
+ bl[2] br[2] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_5 
+ bl[3] br[3] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_6 
+ bl[4] br[4] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_7 
+ bl[5] br[5] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_8 
+ bl[6] br[6] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_9 
+ bl[7] br[7] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_10 
+ bl[8] br[8] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_11 
+ bl[9] br[9] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_12 
+ bl[10] br[10] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_13 
+ bl[11] br[11] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_14 
+ bl[12] br[12] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_15 
+ bl[13] br[13] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_16 
+ bl[14] br[14] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_17 
+ bl[15] br[15] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_18 
+ bl[16] br[16] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_19 
+ bl[17] br[17] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_20 
+ bl[18] br[18] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_21 
+ bl[19] br[19] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_22 
+ bl[20] br[20] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_23 
+ bl[21] br[21] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_24 
+ bl[22] br[22] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_25 
+ bl[23] br[23] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_26 
+ bl[24] br[24] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_27 
+ bl[25] br[25] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_28 
+ bl[26] br[26] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_29 
+ bl[27] br[27] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_30 
+ bl[28] br[28] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_31 
+ bl[29] br[29] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_32 
+ bl[30] br[30] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_33 
+ bl[31] br[31] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_34 
+ bl[32] br[32] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_35 
+ bl[33] br[33] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_36 
+ bl[34] br[34] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_37 
+ bl[35] br[35] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_38 
+ bl[36] br[36] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_39 
+ bl[37] br[37] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_40 
+ bl[38] br[38] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_41 
+ bl[39] br[39] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_42 
+ bl[40] br[40] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_43 
+ bl[41] br[41] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_44 
+ bl[42] br[42] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_45 
+ bl[43] br[43] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_46 
+ bl[44] br[44] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_47 
+ bl[45] br[45] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_48 
+ bl[46] br[46] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_49 
+ bl[47] br[47] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_50 
+ bl[48] br[48] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_51 
+ bl[49] br[49] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_52 
+ bl[50] br[50] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_53 
+ bl[51] br[51] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_54 
+ bl[52] br[52] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_55 
+ bl[53] br[53] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_56 
+ bl[54] br[54] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_57 
+ bl[55] br[55] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_58 
+ bl[56] br[56] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_59 
+ bl[57] br[57] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_60 
+ bl[58] br[58] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_61 
+ bl[59] br[59] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_62 
+ bl[60] br[60] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_63 
+ bl[61] br[61] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_64 
+ bl[62] br[62] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_65 
+ bl[63] br[63] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_66 
+ bl[64] br[64] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_67 
+ bl[65] br[65] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_68 
+ bl[66] br[66] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_69 
+ bl[67] br[67] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_70 
+ bl[68] br[68] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_71 
+ bl[69] br[69] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_72 
+ bl[70] br[70] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_73 
+ bl[71] br[71] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_74 
+ bl[72] br[72] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_75 
+ bl[73] br[73] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_76 
+ bl[74] br[74] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_77 
+ bl[75] br[75] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_78 
+ bl[76] br[76] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_79 
+ bl[77] br[77] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_80 
+ bl[78] br[78] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_81 
+ bl[79] br[79] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_82 
+ bl[80] br[80] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_83 
+ bl[81] br[81] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_84 
+ bl[82] br[82] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_85 
+ bl[83] br[83] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_86 
+ bl[84] br[84] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_87 
+ bl[85] br[85] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_88 
+ bl[86] br[86] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_89 
+ bl[87] br[87] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_90 
+ bl[88] br[88] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_91 
+ bl[89] br[89] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_92 
+ bl[90] br[90] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_93 
+ bl[91] br[91] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_94 
+ bl[92] br[92] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_95 
+ bl[93] br[93] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_96 
+ bl[94] br[94] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_97 
+ bl[95] br[95] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_98 
+ bl[96] br[96] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_99 
+ bl[97] br[97] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_100 
+ bl[98] br[98] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_101 
+ bl[99] br[99] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_102 
+ bl[100] br[100] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_103 
+ bl[101] br[101] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_104 
+ bl[102] br[102] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_105 
+ bl[103] br[103] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_106 
+ bl[104] br[104] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_107 
+ bl[105] br[105] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_108 
+ bl[106] br[106] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_109 
+ bl[107] br[107] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_110 
+ bl[108] br[108] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_111 
+ bl[109] br[109] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_112 
+ bl[110] br[110] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_113 
+ bl[111] br[111] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_114 
+ bl[112] br[112] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_115 
+ bl[113] br[113] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_116 
+ bl[114] br[114] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_117 
+ bl[115] br[115] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_118 
+ bl[116] br[116] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_119 
+ bl[117] br[117] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_120 
+ bl[118] br[118] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_121 
+ bl[119] br[119] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_122 
+ bl[120] br[120] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_123 
+ bl[121] br[121] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_124 
+ bl[122] br[122] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_125 
+ bl[123] br[123] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_126 
+ bl[124] br[124] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_127 
+ bl[125] br[125] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_128 
+ bl[126] br[126] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_129 
+ bl[127] br[127] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_130 
+ bl[128] br[128] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_131 
+ bl[129] br[129] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_132 
+ bl[130] br[130] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_133 
+ bl[131] br[131] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_134 
+ bl[132] br[132] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_135 
+ bl[133] br[133] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_136 
+ bl[134] br[134] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_137 
+ bl[135] br[135] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_138 
+ bl[136] br[136] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_139 
+ bl[137] br[137] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_140 
+ bl[138] br[138] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_141 
+ bl[139] br[139] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_142 
+ bl[140] br[140] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_143 
+ bl[141] br[141] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_144 
+ bl[142] br[142] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_145 
+ bl[143] br[143] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_146 
+ bl[144] br[144] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_147 
+ bl[145] br[145] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_148 
+ bl[146] br[146] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_149 
+ bl[147] br[147] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_150 
+ bl[148] br[148] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_151 
+ bl[149] br[149] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_152 
+ bl[150] br[150] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_153 
+ bl[151] br[151] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_154 
+ bl[152] br[152] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_155 
+ bl[153] br[153] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_156 
+ bl[154] br[154] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_157 
+ bl[155] br[155] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_158 
+ bl[156] br[156] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_159 
+ bl[157] br[157] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_160 
+ bl[158] br[158] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_161 
+ bl[159] br[159] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_162 
+ bl[160] br[160] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_163 
+ bl[161] br[161] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_164 
+ bl[162] br[162] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_165 
+ bl[163] br[163] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_166 
+ bl[164] br[164] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_167 
+ bl[165] br[165] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_168 
+ bl[166] br[166] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_169 
+ bl[167] br[167] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_170 
+ bl[168] br[168] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_171 
+ bl[169] br[169] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_172 
+ bl[170] br[170] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_173 
+ bl[171] br[171] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_174 
+ bl[172] br[172] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_175 
+ bl[173] br[173] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_176 
+ bl[174] br[174] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_177 
+ bl[175] br[175] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_178 
+ bl[176] br[176] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_179 
+ bl[177] br[177] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_180 
+ bl[178] br[178] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_181 
+ bl[179] br[179] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_182 
+ bl[180] br[180] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_183 
+ bl[181] br[181] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_184 
+ bl[182] br[182] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_185 
+ bl[183] br[183] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_186 
+ bl[184] br[184] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_187 
+ bl[185] br[185] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_188 
+ bl[186] br[186] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_189 
+ bl[187] br[187] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_190 
+ bl[188] br[188] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_191 
+ bl[189] br[189] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_192 
+ bl[190] br[190] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_193 
+ bl[191] br[191] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_194 
+ bl[192] br[192] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_195 
+ bl[193] br[193] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_196 
+ bl[194] br[194] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_197 
+ bl[195] br[195] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_198 
+ bl[196] br[196] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_199 
+ bl[197] br[197] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_200 
+ bl[198] br[198] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_201 
+ bl[199] br[199] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_202 
+ bl[200] br[200] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_203 
+ bl[201] br[201] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_204 
+ bl[202] br[202] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_205 
+ bl[203] br[203] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_206 
+ bl[204] br[204] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_207 
+ bl[205] br[205] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_208 
+ bl[206] br[206] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_209 
+ bl[207] br[207] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_210 
+ bl[208] br[208] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_211 
+ bl[209] br[209] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_212 
+ bl[210] br[210] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_213 
+ bl[211] br[211] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_214 
+ bl[212] br[212] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_215 
+ bl[213] br[213] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_216 
+ bl[214] br[214] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_217 
+ bl[215] br[215] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_218 
+ bl[216] br[216] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_219 
+ bl[217] br[217] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_220 
+ bl[218] br[218] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_221 
+ bl[219] br[219] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_222 
+ bl[220] br[220] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_223 
+ bl[221] br[221] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_224 
+ bl[222] br[222] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_225 
+ bl[223] br[223] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_226 
+ bl[224] br[224] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_227 
+ bl[225] br[225] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_228 
+ bl[226] br[226] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_229 
+ bl[227] br[227] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_230 
+ bl[228] br[228] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_231 
+ bl[229] br[229] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_232 
+ bl[230] br[230] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_233 
+ bl[231] br[231] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_234 
+ bl[232] br[232] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_235 
+ bl[233] br[233] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_236 
+ bl[234] br[234] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_237 
+ bl[235] br[235] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_238 
+ bl[236] br[236] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_239 
+ bl[237] br[237] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_240 
+ bl[238] br[238] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_241 
+ bl[239] br[239] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_242 
+ bl[240] br[240] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_243 
+ bl[241] br[241] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_244 
+ bl[242] br[242] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_245 
+ bl[243] br[243] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_246 
+ bl[244] br[244] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_247 
+ bl[245] br[245] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_248 
+ bl[246] br[246] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_249 
+ bl[247] br[247] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_250 
+ bl[248] br[248] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_251 
+ bl[249] br[249] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_252 
+ bl[250] br[250] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_253 
+ bl[251] br[251] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_254 
+ bl[252] br[252] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_255 
+ bl[253] br[253] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_256 
+ bl[254] br[254] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_257 
+ bl[255] br[255] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_258 
+ vdd vdd vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_259 
+ vdd vdd vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_0 
+ vdd vdd vss vdd vpb vnb wl[6] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_8_1 
+ rbl rbr vss vdd vpb vnb wl[6] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_8_2 
+ bl[0] br[0] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_3 
+ bl[1] br[1] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_4 
+ bl[2] br[2] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_5 
+ bl[3] br[3] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_6 
+ bl[4] br[4] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_7 
+ bl[5] br[5] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_8 
+ bl[6] br[6] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_9 
+ bl[7] br[7] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_10 
+ bl[8] br[8] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_11 
+ bl[9] br[9] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_12 
+ bl[10] br[10] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_13 
+ bl[11] br[11] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_14 
+ bl[12] br[12] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_15 
+ bl[13] br[13] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_16 
+ bl[14] br[14] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_17 
+ bl[15] br[15] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_18 
+ bl[16] br[16] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_19 
+ bl[17] br[17] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_20 
+ bl[18] br[18] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_21 
+ bl[19] br[19] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_22 
+ bl[20] br[20] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_23 
+ bl[21] br[21] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_24 
+ bl[22] br[22] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_25 
+ bl[23] br[23] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_26 
+ bl[24] br[24] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_27 
+ bl[25] br[25] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_28 
+ bl[26] br[26] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_29 
+ bl[27] br[27] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_30 
+ bl[28] br[28] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_31 
+ bl[29] br[29] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_32 
+ bl[30] br[30] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_33 
+ bl[31] br[31] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_34 
+ bl[32] br[32] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_35 
+ bl[33] br[33] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_36 
+ bl[34] br[34] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_37 
+ bl[35] br[35] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_38 
+ bl[36] br[36] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_39 
+ bl[37] br[37] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_40 
+ bl[38] br[38] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_41 
+ bl[39] br[39] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_42 
+ bl[40] br[40] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_43 
+ bl[41] br[41] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_44 
+ bl[42] br[42] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_45 
+ bl[43] br[43] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_46 
+ bl[44] br[44] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_47 
+ bl[45] br[45] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_48 
+ bl[46] br[46] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_49 
+ bl[47] br[47] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_50 
+ bl[48] br[48] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_51 
+ bl[49] br[49] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_52 
+ bl[50] br[50] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_53 
+ bl[51] br[51] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_54 
+ bl[52] br[52] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_55 
+ bl[53] br[53] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_56 
+ bl[54] br[54] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_57 
+ bl[55] br[55] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_58 
+ bl[56] br[56] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_59 
+ bl[57] br[57] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_60 
+ bl[58] br[58] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_61 
+ bl[59] br[59] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_62 
+ bl[60] br[60] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_63 
+ bl[61] br[61] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_64 
+ bl[62] br[62] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_65 
+ bl[63] br[63] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_66 
+ bl[64] br[64] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_67 
+ bl[65] br[65] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_68 
+ bl[66] br[66] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_69 
+ bl[67] br[67] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_70 
+ bl[68] br[68] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_71 
+ bl[69] br[69] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_72 
+ bl[70] br[70] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_73 
+ bl[71] br[71] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_74 
+ bl[72] br[72] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_75 
+ bl[73] br[73] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_76 
+ bl[74] br[74] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_77 
+ bl[75] br[75] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_78 
+ bl[76] br[76] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_79 
+ bl[77] br[77] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_80 
+ bl[78] br[78] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_81 
+ bl[79] br[79] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_82 
+ bl[80] br[80] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_83 
+ bl[81] br[81] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_84 
+ bl[82] br[82] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_85 
+ bl[83] br[83] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_86 
+ bl[84] br[84] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_87 
+ bl[85] br[85] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_88 
+ bl[86] br[86] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_89 
+ bl[87] br[87] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_90 
+ bl[88] br[88] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_91 
+ bl[89] br[89] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_92 
+ bl[90] br[90] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_93 
+ bl[91] br[91] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_94 
+ bl[92] br[92] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_95 
+ bl[93] br[93] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_96 
+ bl[94] br[94] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_97 
+ bl[95] br[95] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_98 
+ bl[96] br[96] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_99 
+ bl[97] br[97] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_100 
+ bl[98] br[98] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_101 
+ bl[99] br[99] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_102 
+ bl[100] br[100] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_103 
+ bl[101] br[101] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_104 
+ bl[102] br[102] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_105 
+ bl[103] br[103] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_106 
+ bl[104] br[104] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_107 
+ bl[105] br[105] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_108 
+ bl[106] br[106] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_109 
+ bl[107] br[107] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_110 
+ bl[108] br[108] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_111 
+ bl[109] br[109] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_112 
+ bl[110] br[110] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_113 
+ bl[111] br[111] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_114 
+ bl[112] br[112] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_115 
+ bl[113] br[113] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_116 
+ bl[114] br[114] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_117 
+ bl[115] br[115] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_118 
+ bl[116] br[116] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_119 
+ bl[117] br[117] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_120 
+ bl[118] br[118] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_121 
+ bl[119] br[119] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_122 
+ bl[120] br[120] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_123 
+ bl[121] br[121] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_124 
+ bl[122] br[122] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_125 
+ bl[123] br[123] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_126 
+ bl[124] br[124] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_127 
+ bl[125] br[125] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_128 
+ bl[126] br[126] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_129 
+ bl[127] br[127] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_130 
+ bl[128] br[128] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_131 
+ bl[129] br[129] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_132 
+ bl[130] br[130] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_133 
+ bl[131] br[131] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_134 
+ bl[132] br[132] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_135 
+ bl[133] br[133] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_136 
+ bl[134] br[134] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_137 
+ bl[135] br[135] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_138 
+ bl[136] br[136] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_139 
+ bl[137] br[137] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_140 
+ bl[138] br[138] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_141 
+ bl[139] br[139] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_142 
+ bl[140] br[140] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_143 
+ bl[141] br[141] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_144 
+ bl[142] br[142] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_145 
+ bl[143] br[143] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_146 
+ bl[144] br[144] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_147 
+ bl[145] br[145] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_148 
+ bl[146] br[146] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_149 
+ bl[147] br[147] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_150 
+ bl[148] br[148] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_151 
+ bl[149] br[149] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_152 
+ bl[150] br[150] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_153 
+ bl[151] br[151] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_154 
+ bl[152] br[152] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_155 
+ bl[153] br[153] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_156 
+ bl[154] br[154] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_157 
+ bl[155] br[155] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_158 
+ bl[156] br[156] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_159 
+ bl[157] br[157] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_160 
+ bl[158] br[158] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_161 
+ bl[159] br[159] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_162 
+ bl[160] br[160] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_163 
+ bl[161] br[161] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_164 
+ bl[162] br[162] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_165 
+ bl[163] br[163] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_166 
+ bl[164] br[164] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_167 
+ bl[165] br[165] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_168 
+ bl[166] br[166] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_169 
+ bl[167] br[167] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_170 
+ bl[168] br[168] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_171 
+ bl[169] br[169] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_172 
+ bl[170] br[170] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_173 
+ bl[171] br[171] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_174 
+ bl[172] br[172] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_175 
+ bl[173] br[173] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_176 
+ bl[174] br[174] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_177 
+ bl[175] br[175] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_178 
+ bl[176] br[176] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_179 
+ bl[177] br[177] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_180 
+ bl[178] br[178] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_181 
+ bl[179] br[179] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_182 
+ bl[180] br[180] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_183 
+ bl[181] br[181] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_184 
+ bl[182] br[182] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_185 
+ bl[183] br[183] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_186 
+ bl[184] br[184] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_187 
+ bl[185] br[185] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_188 
+ bl[186] br[186] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_189 
+ bl[187] br[187] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_190 
+ bl[188] br[188] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_191 
+ bl[189] br[189] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_192 
+ bl[190] br[190] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_193 
+ bl[191] br[191] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_194 
+ bl[192] br[192] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_195 
+ bl[193] br[193] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_196 
+ bl[194] br[194] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_197 
+ bl[195] br[195] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_198 
+ bl[196] br[196] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_199 
+ bl[197] br[197] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_200 
+ bl[198] br[198] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_201 
+ bl[199] br[199] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_202 
+ bl[200] br[200] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_203 
+ bl[201] br[201] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_204 
+ bl[202] br[202] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_205 
+ bl[203] br[203] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_206 
+ bl[204] br[204] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_207 
+ bl[205] br[205] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_208 
+ bl[206] br[206] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_209 
+ bl[207] br[207] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_210 
+ bl[208] br[208] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_211 
+ bl[209] br[209] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_212 
+ bl[210] br[210] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_213 
+ bl[211] br[211] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_214 
+ bl[212] br[212] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_215 
+ bl[213] br[213] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_216 
+ bl[214] br[214] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_217 
+ bl[215] br[215] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_218 
+ bl[216] br[216] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_219 
+ bl[217] br[217] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_220 
+ bl[218] br[218] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_221 
+ bl[219] br[219] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_222 
+ bl[220] br[220] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_223 
+ bl[221] br[221] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_224 
+ bl[222] br[222] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_225 
+ bl[223] br[223] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_226 
+ bl[224] br[224] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_227 
+ bl[225] br[225] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_228 
+ bl[226] br[226] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_229 
+ bl[227] br[227] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_230 
+ bl[228] br[228] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_231 
+ bl[229] br[229] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_232 
+ bl[230] br[230] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_233 
+ bl[231] br[231] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_234 
+ bl[232] br[232] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_235 
+ bl[233] br[233] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_236 
+ bl[234] br[234] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_237 
+ bl[235] br[235] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_238 
+ bl[236] br[236] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_239 
+ bl[237] br[237] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_240 
+ bl[238] br[238] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_241 
+ bl[239] br[239] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_242 
+ bl[240] br[240] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_243 
+ bl[241] br[241] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_244 
+ bl[242] br[242] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_245 
+ bl[243] br[243] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_246 
+ bl[244] br[244] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_247 
+ bl[245] br[245] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_248 
+ bl[246] br[246] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_249 
+ bl[247] br[247] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_250 
+ bl[248] br[248] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_251 
+ bl[249] br[249] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_252 
+ bl[250] br[250] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_253 
+ bl[251] br[251] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_254 
+ bl[252] br[252] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_255 
+ bl[253] br[253] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_256 
+ bl[254] br[254] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_257 
+ bl[255] br[255] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_258 
+ vdd vdd vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_259 
+ vdd vdd vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_0 
+ vdd vdd vss vdd vpb vnb wl[7] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_9_1 
+ rbl rbr vss vdd vpb vnb wl[7] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_9_2 
+ bl[0] br[0] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_3 
+ bl[1] br[1] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_4 
+ bl[2] br[2] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_5 
+ bl[3] br[3] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_6 
+ bl[4] br[4] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_7 
+ bl[5] br[5] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_8 
+ bl[6] br[6] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_9 
+ bl[7] br[7] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_10 
+ bl[8] br[8] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_11 
+ bl[9] br[9] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_12 
+ bl[10] br[10] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_13 
+ bl[11] br[11] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_14 
+ bl[12] br[12] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_15 
+ bl[13] br[13] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_16 
+ bl[14] br[14] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_17 
+ bl[15] br[15] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_18 
+ bl[16] br[16] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_19 
+ bl[17] br[17] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_20 
+ bl[18] br[18] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_21 
+ bl[19] br[19] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_22 
+ bl[20] br[20] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_23 
+ bl[21] br[21] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_24 
+ bl[22] br[22] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_25 
+ bl[23] br[23] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_26 
+ bl[24] br[24] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_27 
+ bl[25] br[25] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_28 
+ bl[26] br[26] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_29 
+ bl[27] br[27] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_30 
+ bl[28] br[28] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_31 
+ bl[29] br[29] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_32 
+ bl[30] br[30] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_33 
+ bl[31] br[31] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_34 
+ bl[32] br[32] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_35 
+ bl[33] br[33] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_36 
+ bl[34] br[34] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_37 
+ bl[35] br[35] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_38 
+ bl[36] br[36] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_39 
+ bl[37] br[37] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_40 
+ bl[38] br[38] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_41 
+ bl[39] br[39] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_42 
+ bl[40] br[40] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_43 
+ bl[41] br[41] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_44 
+ bl[42] br[42] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_45 
+ bl[43] br[43] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_46 
+ bl[44] br[44] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_47 
+ bl[45] br[45] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_48 
+ bl[46] br[46] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_49 
+ bl[47] br[47] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_50 
+ bl[48] br[48] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_51 
+ bl[49] br[49] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_52 
+ bl[50] br[50] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_53 
+ bl[51] br[51] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_54 
+ bl[52] br[52] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_55 
+ bl[53] br[53] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_56 
+ bl[54] br[54] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_57 
+ bl[55] br[55] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_58 
+ bl[56] br[56] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_59 
+ bl[57] br[57] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_60 
+ bl[58] br[58] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_61 
+ bl[59] br[59] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_62 
+ bl[60] br[60] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_63 
+ bl[61] br[61] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_64 
+ bl[62] br[62] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_65 
+ bl[63] br[63] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_66 
+ bl[64] br[64] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_67 
+ bl[65] br[65] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_68 
+ bl[66] br[66] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_69 
+ bl[67] br[67] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_70 
+ bl[68] br[68] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_71 
+ bl[69] br[69] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_72 
+ bl[70] br[70] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_73 
+ bl[71] br[71] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_74 
+ bl[72] br[72] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_75 
+ bl[73] br[73] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_76 
+ bl[74] br[74] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_77 
+ bl[75] br[75] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_78 
+ bl[76] br[76] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_79 
+ bl[77] br[77] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_80 
+ bl[78] br[78] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_81 
+ bl[79] br[79] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_82 
+ bl[80] br[80] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_83 
+ bl[81] br[81] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_84 
+ bl[82] br[82] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_85 
+ bl[83] br[83] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_86 
+ bl[84] br[84] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_87 
+ bl[85] br[85] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_88 
+ bl[86] br[86] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_89 
+ bl[87] br[87] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_90 
+ bl[88] br[88] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_91 
+ bl[89] br[89] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_92 
+ bl[90] br[90] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_93 
+ bl[91] br[91] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_94 
+ bl[92] br[92] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_95 
+ bl[93] br[93] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_96 
+ bl[94] br[94] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_97 
+ bl[95] br[95] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_98 
+ bl[96] br[96] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_99 
+ bl[97] br[97] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_100 
+ bl[98] br[98] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_101 
+ bl[99] br[99] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_102 
+ bl[100] br[100] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_103 
+ bl[101] br[101] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_104 
+ bl[102] br[102] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_105 
+ bl[103] br[103] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_106 
+ bl[104] br[104] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_107 
+ bl[105] br[105] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_108 
+ bl[106] br[106] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_109 
+ bl[107] br[107] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_110 
+ bl[108] br[108] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_111 
+ bl[109] br[109] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_112 
+ bl[110] br[110] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_113 
+ bl[111] br[111] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_114 
+ bl[112] br[112] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_115 
+ bl[113] br[113] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_116 
+ bl[114] br[114] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_117 
+ bl[115] br[115] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_118 
+ bl[116] br[116] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_119 
+ bl[117] br[117] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_120 
+ bl[118] br[118] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_121 
+ bl[119] br[119] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_122 
+ bl[120] br[120] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_123 
+ bl[121] br[121] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_124 
+ bl[122] br[122] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_125 
+ bl[123] br[123] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_126 
+ bl[124] br[124] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_127 
+ bl[125] br[125] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_128 
+ bl[126] br[126] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_129 
+ bl[127] br[127] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_130 
+ bl[128] br[128] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_131 
+ bl[129] br[129] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_132 
+ bl[130] br[130] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_133 
+ bl[131] br[131] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_134 
+ bl[132] br[132] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_135 
+ bl[133] br[133] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_136 
+ bl[134] br[134] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_137 
+ bl[135] br[135] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_138 
+ bl[136] br[136] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_139 
+ bl[137] br[137] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_140 
+ bl[138] br[138] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_141 
+ bl[139] br[139] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_142 
+ bl[140] br[140] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_143 
+ bl[141] br[141] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_144 
+ bl[142] br[142] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_145 
+ bl[143] br[143] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_146 
+ bl[144] br[144] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_147 
+ bl[145] br[145] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_148 
+ bl[146] br[146] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_149 
+ bl[147] br[147] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_150 
+ bl[148] br[148] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_151 
+ bl[149] br[149] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_152 
+ bl[150] br[150] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_153 
+ bl[151] br[151] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_154 
+ bl[152] br[152] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_155 
+ bl[153] br[153] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_156 
+ bl[154] br[154] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_157 
+ bl[155] br[155] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_158 
+ bl[156] br[156] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_159 
+ bl[157] br[157] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_160 
+ bl[158] br[158] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_161 
+ bl[159] br[159] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_162 
+ bl[160] br[160] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_163 
+ bl[161] br[161] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_164 
+ bl[162] br[162] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_165 
+ bl[163] br[163] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_166 
+ bl[164] br[164] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_167 
+ bl[165] br[165] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_168 
+ bl[166] br[166] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_169 
+ bl[167] br[167] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_170 
+ bl[168] br[168] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_171 
+ bl[169] br[169] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_172 
+ bl[170] br[170] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_173 
+ bl[171] br[171] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_174 
+ bl[172] br[172] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_175 
+ bl[173] br[173] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_176 
+ bl[174] br[174] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_177 
+ bl[175] br[175] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_178 
+ bl[176] br[176] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_179 
+ bl[177] br[177] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_180 
+ bl[178] br[178] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_181 
+ bl[179] br[179] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_182 
+ bl[180] br[180] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_183 
+ bl[181] br[181] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_184 
+ bl[182] br[182] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_185 
+ bl[183] br[183] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_186 
+ bl[184] br[184] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_187 
+ bl[185] br[185] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_188 
+ bl[186] br[186] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_189 
+ bl[187] br[187] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_190 
+ bl[188] br[188] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_191 
+ bl[189] br[189] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_192 
+ bl[190] br[190] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_193 
+ bl[191] br[191] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_194 
+ bl[192] br[192] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_195 
+ bl[193] br[193] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_196 
+ bl[194] br[194] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_197 
+ bl[195] br[195] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_198 
+ bl[196] br[196] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_199 
+ bl[197] br[197] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_200 
+ bl[198] br[198] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_201 
+ bl[199] br[199] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_202 
+ bl[200] br[200] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_203 
+ bl[201] br[201] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_204 
+ bl[202] br[202] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_205 
+ bl[203] br[203] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_206 
+ bl[204] br[204] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_207 
+ bl[205] br[205] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_208 
+ bl[206] br[206] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_209 
+ bl[207] br[207] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_210 
+ bl[208] br[208] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_211 
+ bl[209] br[209] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_212 
+ bl[210] br[210] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_213 
+ bl[211] br[211] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_214 
+ bl[212] br[212] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_215 
+ bl[213] br[213] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_216 
+ bl[214] br[214] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_217 
+ bl[215] br[215] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_218 
+ bl[216] br[216] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_219 
+ bl[217] br[217] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_220 
+ bl[218] br[218] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_221 
+ bl[219] br[219] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_222 
+ bl[220] br[220] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_223 
+ bl[221] br[221] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_224 
+ bl[222] br[222] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_225 
+ bl[223] br[223] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_226 
+ bl[224] br[224] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_227 
+ bl[225] br[225] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_228 
+ bl[226] br[226] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_229 
+ bl[227] br[227] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_230 
+ bl[228] br[228] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_231 
+ bl[229] br[229] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_232 
+ bl[230] br[230] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_233 
+ bl[231] br[231] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_234 
+ bl[232] br[232] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_235 
+ bl[233] br[233] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_236 
+ bl[234] br[234] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_237 
+ bl[235] br[235] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_238 
+ bl[236] br[236] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_239 
+ bl[237] br[237] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_240 
+ bl[238] br[238] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_241 
+ bl[239] br[239] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_242 
+ bl[240] br[240] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_243 
+ bl[241] br[241] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_244 
+ bl[242] br[242] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_245 
+ bl[243] br[243] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_246 
+ bl[244] br[244] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_247 
+ bl[245] br[245] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_248 
+ bl[246] br[246] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_249 
+ bl[247] br[247] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_250 
+ bl[248] br[248] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_251 
+ bl[249] br[249] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_252 
+ bl[250] br[250] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_253 
+ bl[251] br[251] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_254 
+ bl[252] br[252] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_255 
+ bl[253] br[253] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_256 
+ bl[254] br[254] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_257 
+ bl[255] br[255] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_258 
+ vdd vdd vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_259 
+ vdd vdd vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_0 
+ vdd vdd vss vdd vpb vnb wl[8] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_10_1 
+ rbl rbr vss vdd vpb vnb wl[8] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_10_2 
+ bl[0] br[0] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_3 
+ bl[1] br[1] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_4 
+ bl[2] br[2] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_5 
+ bl[3] br[3] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_6 
+ bl[4] br[4] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_7 
+ bl[5] br[5] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_8 
+ bl[6] br[6] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_9 
+ bl[7] br[7] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_10 
+ bl[8] br[8] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_11 
+ bl[9] br[9] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_12 
+ bl[10] br[10] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_13 
+ bl[11] br[11] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_14 
+ bl[12] br[12] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_15 
+ bl[13] br[13] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_16 
+ bl[14] br[14] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_17 
+ bl[15] br[15] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_18 
+ bl[16] br[16] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_19 
+ bl[17] br[17] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_20 
+ bl[18] br[18] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_21 
+ bl[19] br[19] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_22 
+ bl[20] br[20] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_23 
+ bl[21] br[21] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_24 
+ bl[22] br[22] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_25 
+ bl[23] br[23] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_26 
+ bl[24] br[24] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_27 
+ bl[25] br[25] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_28 
+ bl[26] br[26] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_29 
+ bl[27] br[27] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_30 
+ bl[28] br[28] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_31 
+ bl[29] br[29] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_32 
+ bl[30] br[30] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_33 
+ bl[31] br[31] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_34 
+ bl[32] br[32] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_35 
+ bl[33] br[33] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_36 
+ bl[34] br[34] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_37 
+ bl[35] br[35] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_38 
+ bl[36] br[36] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_39 
+ bl[37] br[37] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_40 
+ bl[38] br[38] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_41 
+ bl[39] br[39] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_42 
+ bl[40] br[40] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_43 
+ bl[41] br[41] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_44 
+ bl[42] br[42] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_45 
+ bl[43] br[43] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_46 
+ bl[44] br[44] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_47 
+ bl[45] br[45] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_48 
+ bl[46] br[46] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_49 
+ bl[47] br[47] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_50 
+ bl[48] br[48] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_51 
+ bl[49] br[49] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_52 
+ bl[50] br[50] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_53 
+ bl[51] br[51] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_54 
+ bl[52] br[52] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_55 
+ bl[53] br[53] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_56 
+ bl[54] br[54] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_57 
+ bl[55] br[55] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_58 
+ bl[56] br[56] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_59 
+ bl[57] br[57] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_60 
+ bl[58] br[58] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_61 
+ bl[59] br[59] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_62 
+ bl[60] br[60] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_63 
+ bl[61] br[61] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_64 
+ bl[62] br[62] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_65 
+ bl[63] br[63] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_66 
+ bl[64] br[64] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_67 
+ bl[65] br[65] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_68 
+ bl[66] br[66] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_69 
+ bl[67] br[67] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_70 
+ bl[68] br[68] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_71 
+ bl[69] br[69] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_72 
+ bl[70] br[70] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_73 
+ bl[71] br[71] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_74 
+ bl[72] br[72] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_75 
+ bl[73] br[73] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_76 
+ bl[74] br[74] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_77 
+ bl[75] br[75] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_78 
+ bl[76] br[76] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_79 
+ bl[77] br[77] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_80 
+ bl[78] br[78] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_81 
+ bl[79] br[79] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_82 
+ bl[80] br[80] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_83 
+ bl[81] br[81] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_84 
+ bl[82] br[82] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_85 
+ bl[83] br[83] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_86 
+ bl[84] br[84] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_87 
+ bl[85] br[85] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_88 
+ bl[86] br[86] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_89 
+ bl[87] br[87] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_90 
+ bl[88] br[88] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_91 
+ bl[89] br[89] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_92 
+ bl[90] br[90] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_93 
+ bl[91] br[91] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_94 
+ bl[92] br[92] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_95 
+ bl[93] br[93] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_96 
+ bl[94] br[94] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_97 
+ bl[95] br[95] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_98 
+ bl[96] br[96] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_99 
+ bl[97] br[97] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_100 
+ bl[98] br[98] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_101 
+ bl[99] br[99] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_102 
+ bl[100] br[100] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_103 
+ bl[101] br[101] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_104 
+ bl[102] br[102] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_105 
+ bl[103] br[103] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_106 
+ bl[104] br[104] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_107 
+ bl[105] br[105] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_108 
+ bl[106] br[106] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_109 
+ bl[107] br[107] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_110 
+ bl[108] br[108] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_111 
+ bl[109] br[109] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_112 
+ bl[110] br[110] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_113 
+ bl[111] br[111] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_114 
+ bl[112] br[112] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_115 
+ bl[113] br[113] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_116 
+ bl[114] br[114] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_117 
+ bl[115] br[115] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_118 
+ bl[116] br[116] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_119 
+ bl[117] br[117] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_120 
+ bl[118] br[118] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_121 
+ bl[119] br[119] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_122 
+ bl[120] br[120] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_123 
+ bl[121] br[121] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_124 
+ bl[122] br[122] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_125 
+ bl[123] br[123] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_126 
+ bl[124] br[124] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_127 
+ bl[125] br[125] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_128 
+ bl[126] br[126] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_129 
+ bl[127] br[127] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_130 
+ bl[128] br[128] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_131 
+ bl[129] br[129] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_132 
+ bl[130] br[130] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_133 
+ bl[131] br[131] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_134 
+ bl[132] br[132] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_135 
+ bl[133] br[133] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_136 
+ bl[134] br[134] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_137 
+ bl[135] br[135] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_138 
+ bl[136] br[136] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_139 
+ bl[137] br[137] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_140 
+ bl[138] br[138] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_141 
+ bl[139] br[139] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_142 
+ bl[140] br[140] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_143 
+ bl[141] br[141] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_144 
+ bl[142] br[142] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_145 
+ bl[143] br[143] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_146 
+ bl[144] br[144] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_147 
+ bl[145] br[145] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_148 
+ bl[146] br[146] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_149 
+ bl[147] br[147] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_150 
+ bl[148] br[148] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_151 
+ bl[149] br[149] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_152 
+ bl[150] br[150] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_153 
+ bl[151] br[151] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_154 
+ bl[152] br[152] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_155 
+ bl[153] br[153] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_156 
+ bl[154] br[154] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_157 
+ bl[155] br[155] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_158 
+ bl[156] br[156] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_159 
+ bl[157] br[157] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_160 
+ bl[158] br[158] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_161 
+ bl[159] br[159] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_162 
+ bl[160] br[160] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_163 
+ bl[161] br[161] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_164 
+ bl[162] br[162] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_165 
+ bl[163] br[163] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_166 
+ bl[164] br[164] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_167 
+ bl[165] br[165] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_168 
+ bl[166] br[166] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_169 
+ bl[167] br[167] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_170 
+ bl[168] br[168] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_171 
+ bl[169] br[169] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_172 
+ bl[170] br[170] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_173 
+ bl[171] br[171] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_174 
+ bl[172] br[172] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_175 
+ bl[173] br[173] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_176 
+ bl[174] br[174] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_177 
+ bl[175] br[175] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_178 
+ bl[176] br[176] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_179 
+ bl[177] br[177] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_180 
+ bl[178] br[178] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_181 
+ bl[179] br[179] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_182 
+ bl[180] br[180] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_183 
+ bl[181] br[181] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_184 
+ bl[182] br[182] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_185 
+ bl[183] br[183] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_186 
+ bl[184] br[184] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_187 
+ bl[185] br[185] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_188 
+ bl[186] br[186] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_189 
+ bl[187] br[187] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_190 
+ bl[188] br[188] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_191 
+ bl[189] br[189] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_192 
+ bl[190] br[190] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_193 
+ bl[191] br[191] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_194 
+ bl[192] br[192] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_195 
+ bl[193] br[193] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_196 
+ bl[194] br[194] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_197 
+ bl[195] br[195] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_198 
+ bl[196] br[196] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_199 
+ bl[197] br[197] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_200 
+ bl[198] br[198] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_201 
+ bl[199] br[199] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_202 
+ bl[200] br[200] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_203 
+ bl[201] br[201] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_204 
+ bl[202] br[202] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_205 
+ bl[203] br[203] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_206 
+ bl[204] br[204] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_207 
+ bl[205] br[205] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_208 
+ bl[206] br[206] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_209 
+ bl[207] br[207] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_210 
+ bl[208] br[208] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_211 
+ bl[209] br[209] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_212 
+ bl[210] br[210] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_213 
+ bl[211] br[211] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_214 
+ bl[212] br[212] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_215 
+ bl[213] br[213] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_216 
+ bl[214] br[214] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_217 
+ bl[215] br[215] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_218 
+ bl[216] br[216] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_219 
+ bl[217] br[217] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_220 
+ bl[218] br[218] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_221 
+ bl[219] br[219] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_222 
+ bl[220] br[220] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_223 
+ bl[221] br[221] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_224 
+ bl[222] br[222] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_225 
+ bl[223] br[223] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_226 
+ bl[224] br[224] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_227 
+ bl[225] br[225] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_228 
+ bl[226] br[226] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_229 
+ bl[227] br[227] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_230 
+ bl[228] br[228] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_231 
+ bl[229] br[229] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_232 
+ bl[230] br[230] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_233 
+ bl[231] br[231] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_234 
+ bl[232] br[232] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_235 
+ bl[233] br[233] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_236 
+ bl[234] br[234] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_237 
+ bl[235] br[235] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_238 
+ bl[236] br[236] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_239 
+ bl[237] br[237] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_240 
+ bl[238] br[238] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_241 
+ bl[239] br[239] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_242 
+ bl[240] br[240] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_243 
+ bl[241] br[241] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_244 
+ bl[242] br[242] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_245 
+ bl[243] br[243] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_246 
+ bl[244] br[244] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_247 
+ bl[245] br[245] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_248 
+ bl[246] br[246] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_249 
+ bl[247] br[247] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_250 
+ bl[248] br[248] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_251 
+ bl[249] br[249] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_252 
+ bl[250] br[250] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_253 
+ bl[251] br[251] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_254 
+ bl[252] br[252] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_255 
+ bl[253] br[253] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_256 
+ bl[254] br[254] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_257 
+ bl[255] br[255] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_258 
+ vdd vdd vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_259 
+ vdd vdd vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_0 
+ vdd vdd vss vdd vpb vnb wl[9] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_11_1 
+ rbl rbr vss vdd vpb vnb wl[9] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_11_2 
+ bl[0] br[0] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_3 
+ bl[1] br[1] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_4 
+ bl[2] br[2] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_5 
+ bl[3] br[3] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_6 
+ bl[4] br[4] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_7 
+ bl[5] br[5] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_8 
+ bl[6] br[6] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_9 
+ bl[7] br[7] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_10 
+ bl[8] br[8] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_11 
+ bl[9] br[9] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_12 
+ bl[10] br[10] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_13 
+ bl[11] br[11] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_14 
+ bl[12] br[12] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_15 
+ bl[13] br[13] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_16 
+ bl[14] br[14] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_17 
+ bl[15] br[15] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_18 
+ bl[16] br[16] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_19 
+ bl[17] br[17] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_20 
+ bl[18] br[18] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_21 
+ bl[19] br[19] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_22 
+ bl[20] br[20] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_23 
+ bl[21] br[21] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_24 
+ bl[22] br[22] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_25 
+ bl[23] br[23] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_26 
+ bl[24] br[24] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_27 
+ bl[25] br[25] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_28 
+ bl[26] br[26] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_29 
+ bl[27] br[27] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_30 
+ bl[28] br[28] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_31 
+ bl[29] br[29] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_32 
+ bl[30] br[30] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_33 
+ bl[31] br[31] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_34 
+ bl[32] br[32] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_35 
+ bl[33] br[33] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_36 
+ bl[34] br[34] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_37 
+ bl[35] br[35] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_38 
+ bl[36] br[36] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_39 
+ bl[37] br[37] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_40 
+ bl[38] br[38] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_41 
+ bl[39] br[39] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_42 
+ bl[40] br[40] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_43 
+ bl[41] br[41] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_44 
+ bl[42] br[42] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_45 
+ bl[43] br[43] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_46 
+ bl[44] br[44] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_47 
+ bl[45] br[45] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_48 
+ bl[46] br[46] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_49 
+ bl[47] br[47] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_50 
+ bl[48] br[48] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_51 
+ bl[49] br[49] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_52 
+ bl[50] br[50] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_53 
+ bl[51] br[51] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_54 
+ bl[52] br[52] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_55 
+ bl[53] br[53] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_56 
+ bl[54] br[54] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_57 
+ bl[55] br[55] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_58 
+ bl[56] br[56] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_59 
+ bl[57] br[57] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_60 
+ bl[58] br[58] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_61 
+ bl[59] br[59] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_62 
+ bl[60] br[60] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_63 
+ bl[61] br[61] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_64 
+ bl[62] br[62] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_65 
+ bl[63] br[63] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_66 
+ bl[64] br[64] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_67 
+ bl[65] br[65] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_68 
+ bl[66] br[66] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_69 
+ bl[67] br[67] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_70 
+ bl[68] br[68] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_71 
+ bl[69] br[69] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_72 
+ bl[70] br[70] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_73 
+ bl[71] br[71] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_74 
+ bl[72] br[72] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_75 
+ bl[73] br[73] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_76 
+ bl[74] br[74] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_77 
+ bl[75] br[75] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_78 
+ bl[76] br[76] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_79 
+ bl[77] br[77] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_80 
+ bl[78] br[78] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_81 
+ bl[79] br[79] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_82 
+ bl[80] br[80] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_83 
+ bl[81] br[81] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_84 
+ bl[82] br[82] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_85 
+ bl[83] br[83] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_86 
+ bl[84] br[84] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_87 
+ bl[85] br[85] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_88 
+ bl[86] br[86] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_89 
+ bl[87] br[87] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_90 
+ bl[88] br[88] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_91 
+ bl[89] br[89] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_92 
+ bl[90] br[90] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_93 
+ bl[91] br[91] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_94 
+ bl[92] br[92] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_95 
+ bl[93] br[93] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_96 
+ bl[94] br[94] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_97 
+ bl[95] br[95] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_98 
+ bl[96] br[96] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_99 
+ bl[97] br[97] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_100 
+ bl[98] br[98] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_101 
+ bl[99] br[99] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_102 
+ bl[100] br[100] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_103 
+ bl[101] br[101] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_104 
+ bl[102] br[102] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_105 
+ bl[103] br[103] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_106 
+ bl[104] br[104] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_107 
+ bl[105] br[105] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_108 
+ bl[106] br[106] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_109 
+ bl[107] br[107] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_110 
+ bl[108] br[108] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_111 
+ bl[109] br[109] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_112 
+ bl[110] br[110] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_113 
+ bl[111] br[111] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_114 
+ bl[112] br[112] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_115 
+ bl[113] br[113] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_116 
+ bl[114] br[114] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_117 
+ bl[115] br[115] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_118 
+ bl[116] br[116] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_119 
+ bl[117] br[117] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_120 
+ bl[118] br[118] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_121 
+ bl[119] br[119] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_122 
+ bl[120] br[120] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_123 
+ bl[121] br[121] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_124 
+ bl[122] br[122] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_125 
+ bl[123] br[123] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_126 
+ bl[124] br[124] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_127 
+ bl[125] br[125] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_128 
+ bl[126] br[126] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_129 
+ bl[127] br[127] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_130 
+ bl[128] br[128] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_131 
+ bl[129] br[129] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_132 
+ bl[130] br[130] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_133 
+ bl[131] br[131] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_134 
+ bl[132] br[132] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_135 
+ bl[133] br[133] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_136 
+ bl[134] br[134] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_137 
+ bl[135] br[135] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_138 
+ bl[136] br[136] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_139 
+ bl[137] br[137] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_140 
+ bl[138] br[138] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_141 
+ bl[139] br[139] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_142 
+ bl[140] br[140] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_143 
+ bl[141] br[141] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_144 
+ bl[142] br[142] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_145 
+ bl[143] br[143] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_146 
+ bl[144] br[144] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_147 
+ bl[145] br[145] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_148 
+ bl[146] br[146] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_149 
+ bl[147] br[147] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_150 
+ bl[148] br[148] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_151 
+ bl[149] br[149] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_152 
+ bl[150] br[150] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_153 
+ bl[151] br[151] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_154 
+ bl[152] br[152] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_155 
+ bl[153] br[153] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_156 
+ bl[154] br[154] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_157 
+ bl[155] br[155] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_158 
+ bl[156] br[156] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_159 
+ bl[157] br[157] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_160 
+ bl[158] br[158] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_161 
+ bl[159] br[159] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_162 
+ bl[160] br[160] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_163 
+ bl[161] br[161] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_164 
+ bl[162] br[162] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_165 
+ bl[163] br[163] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_166 
+ bl[164] br[164] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_167 
+ bl[165] br[165] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_168 
+ bl[166] br[166] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_169 
+ bl[167] br[167] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_170 
+ bl[168] br[168] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_171 
+ bl[169] br[169] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_172 
+ bl[170] br[170] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_173 
+ bl[171] br[171] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_174 
+ bl[172] br[172] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_175 
+ bl[173] br[173] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_176 
+ bl[174] br[174] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_177 
+ bl[175] br[175] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_178 
+ bl[176] br[176] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_179 
+ bl[177] br[177] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_180 
+ bl[178] br[178] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_181 
+ bl[179] br[179] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_182 
+ bl[180] br[180] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_183 
+ bl[181] br[181] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_184 
+ bl[182] br[182] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_185 
+ bl[183] br[183] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_186 
+ bl[184] br[184] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_187 
+ bl[185] br[185] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_188 
+ bl[186] br[186] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_189 
+ bl[187] br[187] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_190 
+ bl[188] br[188] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_191 
+ bl[189] br[189] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_192 
+ bl[190] br[190] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_193 
+ bl[191] br[191] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_194 
+ bl[192] br[192] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_195 
+ bl[193] br[193] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_196 
+ bl[194] br[194] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_197 
+ bl[195] br[195] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_198 
+ bl[196] br[196] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_199 
+ bl[197] br[197] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_200 
+ bl[198] br[198] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_201 
+ bl[199] br[199] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_202 
+ bl[200] br[200] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_203 
+ bl[201] br[201] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_204 
+ bl[202] br[202] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_205 
+ bl[203] br[203] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_206 
+ bl[204] br[204] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_207 
+ bl[205] br[205] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_208 
+ bl[206] br[206] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_209 
+ bl[207] br[207] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_210 
+ bl[208] br[208] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_211 
+ bl[209] br[209] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_212 
+ bl[210] br[210] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_213 
+ bl[211] br[211] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_214 
+ bl[212] br[212] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_215 
+ bl[213] br[213] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_216 
+ bl[214] br[214] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_217 
+ bl[215] br[215] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_218 
+ bl[216] br[216] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_219 
+ bl[217] br[217] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_220 
+ bl[218] br[218] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_221 
+ bl[219] br[219] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_222 
+ bl[220] br[220] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_223 
+ bl[221] br[221] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_224 
+ bl[222] br[222] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_225 
+ bl[223] br[223] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_226 
+ bl[224] br[224] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_227 
+ bl[225] br[225] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_228 
+ bl[226] br[226] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_229 
+ bl[227] br[227] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_230 
+ bl[228] br[228] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_231 
+ bl[229] br[229] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_232 
+ bl[230] br[230] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_233 
+ bl[231] br[231] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_234 
+ bl[232] br[232] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_235 
+ bl[233] br[233] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_236 
+ bl[234] br[234] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_237 
+ bl[235] br[235] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_238 
+ bl[236] br[236] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_239 
+ bl[237] br[237] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_240 
+ bl[238] br[238] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_241 
+ bl[239] br[239] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_242 
+ bl[240] br[240] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_243 
+ bl[241] br[241] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_244 
+ bl[242] br[242] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_245 
+ bl[243] br[243] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_246 
+ bl[244] br[244] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_247 
+ bl[245] br[245] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_248 
+ bl[246] br[246] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_249 
+ bl[247] br[247] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_250 
+ bl[248] br[248] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_251 
+ bl[249] br[249] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_252 
+ bl[250] br[250] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_253 
+ bl[251] br[251] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_254 
+ bl[252] br[252] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_255 
+ bl[253] br[253] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_256 
+ bl[254] br[254] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_257 
+ bl[255] br[255] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_258 
+ vdd vdd vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_259 
+ vdd vdd vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_0 
+ vdd vdd vss vdd vpb vnb wl[10] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_12_1 
+ rbl rbr vss vdd vpb vnb wl[10] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_12_2 
+ bl[0] br[0] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_3 
+ bl[1] br[1] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_4 
+ bl[2] br[2] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_5 
+ bl[3] br[3] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_6 
+ bl[4] br[4] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_7 
+ bl[5] br[5] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_8 
+ bl[6] br[6] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_9 
+ bl[7] br[7] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_10 
+ bl[8] br[8] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_11 
+ bl[9] br[9] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_12 
+ bl[10] br[10] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_13 
+ bl[11] br[11] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_14 
+ bl[12] br[12] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_15 
+ bl[13] br[13] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_16 
+ bl[14] br[14] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_17 
+ bl[15] br[15] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_18 
+ bl[16] br[16] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_19 
+ bl[17] br[17] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_20 
+ bl[18] br[18] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_21 
+ bl[19] br[19] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_22 
+ bl[20] br[20] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_23 
+ bl[21] br[21] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_24 
+ bl[22] br[22] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_25 
+ bl[23] br[23] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_26 
+ bl[24] br[24] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_27 
+ bl[25] br[25] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_28 
+ bl[26] br[26] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_29 
+ bl[27] br[27] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_30 
+ bl[28] br[28] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_31 
+ bl[29] br[29] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_32 
+ bl[30] br[30] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_33 
+ bl[31] br[31] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_34 
+ bl[32] br[32] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_35 
+ bl[33] br[33] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_36 
+ bl[34] br[34] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_37 
+ bl[35] br[35] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_38 
+ bl[36] br[36] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_39 
+ bl[37] br[37] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_40 
+ bl[38] br[38] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_41 
+ bl[39] br[39] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_42 
+ bl[40] br[40] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_43 
+ bl[41] br[41] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_44 
+ bl[42] br[42] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_45 
+ bl[43] br[43] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_46 
+ bl[44] br[44] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_47 
+ bl[45] br[45] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_48 
+ bl[46] br[46] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_49 
+ bl[47] br[47] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_50 
+ bl[48] br[48] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_51 
+ bl[49] br[49] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_52 
+ bl[50] br[50] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_53 
+ bl[51] br[51] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_54 
+ bl[52] br[52] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_55 
+ bl[53] br[53] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_56 
+ bl[54] br[54] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_57 
+ bl[55] br[55] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_58 
+ bl[56] br[56] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_59 
+ bl[57] br[57] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_60 
+ bl[58] br[58] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_61 
+ bl[59] br[59] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_62 
+ bl[60] br[60] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_63 
+ bl[61] br[61] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_64 
+ bl[62] br[62] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_65 
+ bl[63] br[63] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_66 
+ bl[64] br[64] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_67 
+ bl[65] br[65] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_68 
+ bl[66] br[66] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_69 
+ bl[67] br[67] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_70 
+ bl[68] br[68] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_71 
+ bl[69] br[69] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_72 
+ bl[70] br[70] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_73 
+ bl[71] br[71] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_74 
+ bl[72] br[72] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_75 
+ bl[73] br[73] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_76 
+ bl[74] br[74] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_77 
+ bl[75] br[75] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_78 
+ bl[76] br[76] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_79 
+ bl[77] br[77] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_80 
+ bl[78] br[78] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_81 
+ bl[79] br[79] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_82 
+ bl[80] br[80] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_83 
+ bl[81] br[81] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_84 
+ bl[82] br[82] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_85 
+ bl[83] br[83] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_86 
+ bl[84] br[84] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_87 
+ bl[85] br[85] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_88 
+ bl[86] br[86] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_89 
+ bl[87] br[87] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_90 
+ bl[88] br[88] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_91 
+ bl[89] br[89] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_92 
+ bl[90] br[90] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_93 
+ bl[91] br[91] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_94 
+ bl[92] br[92] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_95 
+ bl[93] br[93] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_96 
+ bl[94] br[94] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_97 
+ bl[95] br[95] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_98 
+ bl[96] br[96] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_99 
+ bl[97] br[97] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_100 
+ bl[98] br[98] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_101 
+ bl[99] br[99] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_102 
+ bl[100] br[100] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_103 
+ bl[101] br[101] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_104 
+ bl[102] br[102] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_105 
+ bl[103] br[103] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_106 
+ bl[104] br[104] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_107 
+ bl[105] br[105] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_108 
+ bl[106] br[106] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_109 
+ bl[107] br[107] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_110 
+ bl[108] br[108] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_111 
+ bl[109] br[109] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_112 
+ bl[110] br[110] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_113 
+ bl[111] br[111] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_114 
+ bl[112] br[112] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_115 
+ bl[113] br[113] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_116 
+ bl[114] br[114] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_117 
+ bl[115] br[115] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_118 
+ bl[116] br[116] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_119 
+ bl[117] br[117] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_120 
+ bl[118] br[118] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_121 
+ bl[119] br[119] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_122 
+ bl[120] br[120] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_123 
+ bl[121] br[121] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_124 
+ bl[122] br[122] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_125 
+ bl[123] br[123] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_126 
+ bl[124] br[124] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_127 
+ bl[125] br[125] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_128 
+ bl[126] br[126] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_129 
+ bl[127] br[127] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_130 
+ bl[128] br[128] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_131 
+ bl[129] br[129] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_132 
+ bl[130] br[130] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_133 
+ bl[131] br[131] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_134 
+ bl[132] br[132] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_135 
+ bl[133] br[133] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_136 
+ bl[134] br[134] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_137 
+ bl[135] br[135] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_138 
+ bl[136] br[136] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_139 
+ bl[137] br[137] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_140 
+ bl[138] br[138] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_141 
+ bl[139] br[139] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_142 
+ bl[140] br[140] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_143 
+ bl[141] br[141] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_144 
+ bl[142] br[142] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_145 
+ bl[143] br[143] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_146 
+ bl[144] br[144] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_147 
+ bl[145] br[145] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_148 
+ bl[146] br[146] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_149 
+ bl[147] br[147] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_150 
+ bl[148] br[148] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_151 
+ bl[149] br[149] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_152 
+ bl[150] br[150] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_153 
+ bl[151] br[151] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_154 
+ bl[152] br[152] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_155 
+ bl[153] br[153] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_156 
+ bl[154] br[154] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_157 
+ bl[155] br[155] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_158 
+ bl[156] br[156] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_159 
+ bl[157] br[157] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_160 
+ bl[158] br[158] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_161 
+ bl[159] br[159] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_162 
+ bl[160] br[160] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_163 
+ bl[161] br[161] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_164 
+ bl[162] br[162] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_165 
+ bl[163] br[163] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_166 
+ bl[164] br[164] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_167 
+ bl[165] br[165] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_168 
+ bl[166] br[166] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_169 
+ bl[167] br[167] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_170 
+ bl[168] br[168] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_171 
+ bl[169] br[169] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_172 
+ bl[170] br[170] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_173 
+ bl[171] br[171] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_174 
+ bl[172] br[172] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_175 
+ bl[173] br[173] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_176 
+ bl[174] br[174] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_177 
+ bl[175] br[175] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_178 
+ bl[176] br[176] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_179 
+ bl[177] br[177] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_180 
+ bl[178] br[178] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_181 
+ bl[179] br[179] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_182 
+ bl[180] br[180] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_183 
+ bl[181] br[181] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_184 
+ bl[182] br[182] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_185 
+ bl[183] br[183] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_186 
+ bl[184] br[184] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_187 
+ bl[185] br[185] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_188 
+ bl[186] br[186] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_189 
+ bl[187] br[187] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_190 
+ bl[188] br[188] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_191 
+ bl[189] br[189] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_192 
+ bl[190] br[190] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_193 
+ bl[191] br[191] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_194 
+ bl[192] br[192] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_195 
+ bl[193] br[193] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_196 
+ bl[194] br[194] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_197 
+ bl[195] br[195] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_198 
+ bl[196] br[196] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_199 
+ bl[197] br[197] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_200 
+ bl[198] br[198] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_201 
+ bl[199] br[199] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_202 
+ bl[200] br[200] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_203 
+ bl[201] br[201] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_204 
+ bl[202] br[202] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_205 
+ bl[203] br[203] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_206 
+ bl[204] br[204] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_207 
+ bl[205] br[205] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_208 
+ bl[206] br[206] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_209 
+ bl[207] br[207] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_210 
+ bl[208] br[208] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_211 
+ bl[209] br[209] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_212 
+ bl[210] br[210] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_213 
+ bl[211] br[211] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_214 
+ bl[212] br[212] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_215 
+ bl[213] br[213] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_216 
+ bl[214] br[214] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_217 
+ bl[215] br[215] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_218 
+ bl[216] br[216] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_219 
+ bl[217] br[217] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_220 
+ bl[218] br[218] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_221 
+ bl[219] br[219] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_222 
+ bl[220] br[220] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_223 
+ bl[221] br[221] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_224 
+ bl[222] br[222] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_225 
+ bl[223] br[223] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_226 
+ bl[224] br[224] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_227 
+ bl[225] br[225] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_228 
+ bl[226] br[226] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_229 
+ bl[227] br[227] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_230 
+ bl[228] br[228] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_231 
+ bl[229] br[229] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_232 
+ bl[230] br[230] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_233 
+ bl[231] br[231] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_234 
+ bl[232] br[232] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_235 
+ bl[233] br[233] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_236 
+ bl[234] br[234] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_237 
+ bl[235] br[235] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_238 
+ bl[236] br[236] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_239 
+ bl[237] br[237] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_240 
+ bl[238] br[238] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_241 
+ bl[239] br[239] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_242 
+ bl[240] br[240] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_243 
+ bl[241] br[241] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_244 
+ bl[242] br[242] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_245 
+ bl[243] br[243] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_246 
+ bl[244] br[244] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_247 
+ bl[245] br[245] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_248 
+ bl[246] br[246] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_249 
+ bl[247] br[247] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_250 
+ bl[248] br[248] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_251 
+ bl[249] br[249] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_252 
+ bl[250] br[250] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_253 
+ bl[251] br[251] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_254 
+ bl[252] br[252] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_255 
+ bl[253] br[253] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_256 
+ bl[254] br[254] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_257 
+ bl[255] br[255] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_258 
+ vdd vdd vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_259 
+ vdd vdd vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_0 
+ vdd vdd vss vdd vpb vnb wl[11] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_13_1 
+ rbl rbr vss vdd vpb vnb wl[11] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_13_2 
+ bl[0] br[0] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_3 
+ bl[1] br[1] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_4 
+ bl[2] br[2] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_5 
+ bl[3] br[3] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_6 
+ bl[4] br[4] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_7 
+ bl[5] br[5] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_8 
+ bl[6] br[6] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_9 
+ bl[7] br[7] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_10 
+ bl[8] br[8] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_11 
+ bl[9] br[9] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_12 
+ bl[10] br[10] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_13 
+ bl[11] br[11] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_14 
+ bl[12] br[12] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_15 
+ bl[13] br[13] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_16 
+ bl[14] br[14] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_17 
+ bl[15] br[15] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_18 
+ bl[16] br[16] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_19 
+ bl[17] br[17] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_20 
+ bl[18] br[18] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_21 
+ bl[19] br[19] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_22 
+ bl[20] br[20] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_23 
+ bl[21] br[21] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_24 
+ bl[22] br[22] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_25 
+ bl[23] br[23] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_26 
+ bl[24] br[24] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_27 
+ bl[25] br[25] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_28 
+ bl[26] br[26] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_29 
+ bl[27] br[27] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_30 
+ bl[28] br[28] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_31 
+ bl[29] br[29] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_32 
+ bl[30] br[30] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_33 
+ bl[31] br[31] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_34 
+ bl[32] br[32] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_35 
+ bl[33] br[33] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_36 
+ bl[34] br[34] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_37 
+ bl[35] br[35] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_38 
+ bl[36] br[36] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_39 
+ bl[37] br[37] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_40 
+ bl[38] br[38] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_41 
+ bl[39] br[39] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_42 
+ bl[40] br[40] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_43 
+ bl[41] br[41] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_44 
+ bl[42] br[42] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_45 
+ bl[43] br[43] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_46 
+ bl[44] br[44] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_47 
+ bl[45] br[45] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_48 
+ bl[46] br[46] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_49 
+ bl[47] br[47] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_50 
+ bl[48] br[48] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_51 
+ bl[49] br[49] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_52 
+ bl[50] br[50] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_53 
+ bl[51] br[51] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_54 
+ bl[52] br[52] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_55 
+ bl[53] br[53] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_56 
+ bl[54] br[54] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_57 
+ bl[55] br[55] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_58 
+ bl[56] br[56] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_59 
+ bl[57] br[57] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_60 
+ bl[58] br[58] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_61 
+ bl[59] br[59] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_62 
+ bl[60] br[60] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_63 
+ bl[61] br[61] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_64 
+ bl[62] br[62] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_65 
+ bl[63] br[63] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_66 
+ bl[64] br[64] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_67 
+ bl[65] br[65] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_68 
+ bl[66] br[66] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_69 
+ bl[67] br[67] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_70 
+ bl[68] br[68] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_71 
+ bl[69] br[69] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_72 
+ bl[70] br[70] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_73 
+ bl[71] br[71] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_74 
+ bl[72] br[72] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_75 
+ bl[73] br[73] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_76 
+ bl[74] br[74] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_77 
+ bl[75] br[75] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_78 
+ bl[76] br[76] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_79 
+ bl[77] br[77] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_80 
+ bl[78] br[78] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_81 
+ bl[79] br[79] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_82 
+ bl[80] br[80] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_83 
+ bl[81] br[81] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_84 
+ bl[82] br[82] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_85 
+ bl[83] br[83] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_86 
+ bl[84] br[84] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_87 
+ bl[85] br[85] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_88 
+ bl[86] br[86] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_89 
+ bl[87] br[87] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_90 
+ bl[88] br[88] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_91 
+ bl[89] br[89] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_92 
+ bl[90] br[90] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_93 
+ bl[91] br[91] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_94 
+ bl[92] br[92] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_95 
+ bl[93] br[93] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_96 
+ bl[94] br[94] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_97 
+ bl[95] br[95] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_98 
+ bl[96] br[96] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_99 
+ bl[97] br[97] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_100 
+ bl[98] br[98] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_101 
+ bl[99] br[99] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_102 
+ bl[100] br[100] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_103 
+ bl[101] br[101] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_104 
+ bl[102] br[102] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_105 
+ bl[103] br[103] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_106 
+ bl[104] br[104] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_107 
+ bl[105] br[105] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_108 
+ bl[106] br[106] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_109 
+ bl[107] br[107] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_110 
+ bl[108] br[108] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_111 
+ bl[109] br[109] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_112 
+ bl[110] br[110] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_113 
+ bl[111] br[111] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_114 
+ bl[112] br[112] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_115 
+ bl[113] br[113] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_116 
+ bl[114] br[114] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_117 
+ bl[115] br[115] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_118 
+ bl[116] br[116] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_119 
+ bl[117] br[117] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_120 
+ bl[118] br[118] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_121 
+ bl[119] br[119] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_122 
+ bl[120] br[120] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_123 
+ bl[121] br[121] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_124 
+ bl[122] br[122] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_125 
+ bl[123] br[123] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_126 
+ bl[124] br[124] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_127 
+ bl[125] br[125] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_128 
+ bl[126] br[126] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_129 
+ bl[127] br[127] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_130 
+ bl[128] br[128] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_131 
+ bl[129] br[129] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_132 
+ bl[130] br[130] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_133 
+ bl[131] br[131] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_134 
+ bl[132] br[132] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_135 
+ bl[133] br[133] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_136 
+ bl[134] br[134] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_137 
+ bl[135] br[135] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_138 
+ bl[136] br[136] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_139 
+ bl[137] br[137] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_140 
+ bl[138] br[138] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_141 
+ bl[139] br[139] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_142 
+ bl[140] br[140] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_143 
+ bl[141] br[141] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_144 
+ bl[142] br[142] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_145 
+ bl[143] br[143] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_146 
+ bl[144] br[144] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_147 
+ bl[145] br[145] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_148 
+ bl[146] br[146] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_149 
+ bl[147] br[147] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_150 
+ bl[148] br[148] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_151 
+ bl[149] br[149] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_152 
+ bl[150] br[150] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_153 
+ bl[151] br[151] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_154 
+ bl[152] br[152] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_155 
+ bl[153] br[153] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_156 
+ bl[154] br[154] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_157 
+ bl[155] br[155] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_158 
+ bl[156] br[156] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_159 
+ bl[157] br[157] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_160 
+ bl[158] br[158] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_161 
+ bl[159] br[159] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_162 
+ bl[160] br[160] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_163 
+ bl[161] br[161] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_164 
+ bl[162] br[162] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_165 
+ bl[163] br[163] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_166 
+ bl[164] br[164] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_167 
+ bl[165] br[165] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_168 
+ bl[166] br[166] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_169 
+ bl[167] br[167] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_170 
+ bl[168] br[168] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_171 
+ bl[169] br[169] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_172 
+ bl[170] br[170] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_173 
+ bl[171] br[171] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_174 
+ bl[172] br[172] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_175 
+ bl[173] br[173] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_176 
+ bl[174] br[174] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_177 
+ bl[175] br[175] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_178 
+ bl[176] br[176] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_179 
+ bl[177] br[177] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_180 
+ bl[178] br[178] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_181 
+ bl[179] br[179] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_182 
+ bl[180] br[180] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_183 
+ bl[181] br[181] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_184 
+ bl[182] br[182] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_185 
+ bl[183] br[183] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_186 
+ bl[184] br[184] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_187 
+ bl[185] br[185] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_188 
+ bl[186] br[186] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_189 
+ bl[187] br[187] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_190 
+ bl[188] br[188] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_191 
+ bl[189] br[189] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_192 
+ bl[190] br[190] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_193 
+ bl[191] br[191] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_194 
+ bl[192] br[192] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_195 
+ bl[193] br[193] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_196 
+ bl[194] br[194] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_197 
+ bl[195] br[195] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_198 
+ bl[196] br[196] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_199 
+ bl[197] br[197] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_200 
+ bl[198] br[198] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_201 
+ bl[199] br[199] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_202 
+ bl[200] br[200] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_203 
+ bl[201] br[201] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_204 
+ bl[202] br[202] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_205 
+ bl[203] br[203] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_206 
+ bl[204] br[204] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_207 
+ bl[205] br[205] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_208 
+ bl[206] br[206] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_209 
+ bl[207] br[207] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_210 
+ bl[208] br[208] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_211 
+ bl[209] br[209] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_212 
+ bl[210] br[210] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_213 
+ bl[211] br[211] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_214 
+ bl[212] br[212] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_215 
+ bl[213] br[213] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_216 
+ bl[214] br[214] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_217 
+ bl[215] br[215] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_218 
+ bl[216] br[216] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_219 
+ bl[217] br[217] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_220 
+ bl[218] br[218] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_221 
+ bl[219] br[219] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_222 
+ bl[220] br[220] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_223 
+ bl[221] br[221] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_224 
+ bl[222] br[222] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_225 
+ bl[223] br[223] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_226 
+ bl[224] br[224] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_227 
+ bl[225] br[225] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_228 
+ bl[226] br[226] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_229 
+ bl[227] br[227] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_230 
+ bl[228] br[228] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_231 
+ bl[229] br[229] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_232 
+ bl[230] br[230] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_233 
+ bl[231] br[231] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_234 
+ bl[232] br[232] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_235 
+ bl[233] br[233] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_236 
+ bl[234] br[234] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_237 
+ bl[235] br[235] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_238 
+ bl[236] br[236] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_239 
+ bl[237] br[237] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_240 
+ bl[238] br[238] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_241 
+ bl[239] br[239] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_242 
+ bl[240] br[240] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_243 
+ bl[241] br[241] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_244 
+ bl[242] br[242] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_245 
+ bl[243] br[243] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_246 
+ bl[244] br[244] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_247 
+ bl[245] br[245] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_248 
+ bl[246] br[246] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_249 
+ bl[247] br[247] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_250 
+ bl[248] br[248] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_251 
+ bl[249] br[249] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_252 
+ bl[250] br[250] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_253 
+ bl[251] br[251] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_254 
+ bl[252] br[252] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_255 
+ bl[253] br[253] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_256 
+ bl[254] br[254] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_257 
+ bl[255] br[255] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_258 
+ vdd vdd vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_259 
+ vdd vdd vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_0 
+ vdd vdd vss vdd vpb vnb wl[12] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_14_1 
+ rbl rbr vss vdd vpb vnb wl[12] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_14_2 
+ bl[0] br[0] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_3 
+ bl[1] br[1] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_4 
+ bl[2] br[2] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_5 
+ bl[3] br[3] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_6 
+ bl[4] br[4] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_7 
+ bl[5] br[5] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_8 
+ bl[6] br[6] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_9 
+ bl[7] br[7] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_10 
+ bl[8] br[8] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_11 
+ bl[9] br[9] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_12 
+ bl[10] br[10] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_13 
+ bl[11] br[11] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_14 
+ bl[12] br[12] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_15 
+ bl[13] br[13] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_16 
+ bl[14] br[14] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_17 
+ bl[15] br[15] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_18 
+ bl[16] br[16] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_19 
+ bl[17] br[17] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_20 
+ bl[18] br[18] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_21 
+ bl[19] br[19] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_22 
+ bl[20] br[20] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_23 
+ bl[21] br[21] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_24 
+ bl[22] br[22] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_25 
+ bl[23] br[23] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_26 
+ bl[24] br[24] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_27 
+ bl[25] br[25] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_28 
+ bl[26] br[26] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_29 
+ bl[27] br[27] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_30 
+ bl[28] br[28] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_31 
+ bl[29] br[29] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_32 
+ bl[30] br[30] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_33 
+ bl[31] br[31] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_34 
+ bl[32] br[32] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_35 
+ bl[33] br[33] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_36 
+ bl[34] br[34] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_37 
+ bl[35] br[35] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_38 
+ bl[36] br[36] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_39 
+ bl[37] br[37] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_40 
+ bl[38] br[38] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_41 
+ bl[39] br[39] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_42 
+ bl[40] br[40] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_43 
+ bl[41] br[41] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_44 
+ bl[42] br[42] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_45 
+ bl[43] br[43] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_46 
+ bl[44] br[44] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_47 
+ bl[45] br[45] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_48 
+ bl[46] br[46] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_49 
+ bl[47] br[47] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_50 
+ bl[48] br[48] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_51 
+ bl[49] br[49] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_52 
+ bl[50] br[50] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_53 
+ bl[51] br[51] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_54 
+ bl[52] br[52] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_55 
+ bl[53] br[53] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_56 
+ bl[54] br[54] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_57 
+ bl[55] br[55] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_58 
+ bl[56] br[56] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_59 
+ bl[57] br[57] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_60 
+ bl[58] br[58] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_61 
+ bl[59] br[59] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_62 
+ bl[60] br[60] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_63 
+ bl[61] br[61] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_64 
+ bl[62] br[62] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_65 
+ bl[63] br[63] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_66 
+ bl[64] br[64] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_67 
+ bl[65] br[65] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_68 
+ bl[66] br[66] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_69 
+ bl[67] br[67] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_70 
+ bl[68] br[68] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_71 
+ bl[69] br[69] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_72 
+ bl[70] br[70] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_73 
+ bl[71] br[71] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_74 
+ bl[72] br[72] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_75 
+ bl[73] br[73] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_76 
+ bl[74] br[74] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_77 
+ bl[75] br[75] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_78 
+ bl[76] br[76] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_79 
+ bl[77] br[77] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_80 
+ bl[78] br[78] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_81 
+ bl[79] br[79] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_82 
+ bl[80] br[80] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_83 
+ bl[81] br[81] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_84 
+ bl[82] br[82] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_85 
+ bl[83] br[83] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_86 
+ bl[84] br[84] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_87 
+ bl[85] br[85] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_88 
+ bl[86] br[86] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_89 
+ bl[87] br[87] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_90 
+ bl[88] br[88] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_91 
+ bl[89] br[89] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_92 
+ bl[90] br[90] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_93 
+ bl[91] br[91] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_94 
+ bl[92] br[92] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_95 
+ bl[93] br[93] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_96 
+ bl[94] br[94] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_97 
+ bl[95] br[95] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_98 
+ bl[96] br[96] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_99 
+ bl[97] br[97] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_100 
+ bl[98] br[98] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_101 
+ bl[99] br[99] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_102 
+ bl[100] br[100] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_103 
+ bl[101] br[101] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_104 
+ bl[102] br[102] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_105 
+ bl[103] br[103] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_106 
+ bl[104] br[104] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_107 
+ bl[105] br[105] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_108 
+ bl[106] br[106] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_109 
+ bl[107] br[107] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_110 
+ bl[108] br[108] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_111 
+ bl[109] br[109] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_112 
+ bl[110] br[110] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_113 
+ bl[111] br[111] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_114 
+ bl[112] br[112] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_115 
+ bl[113] br[113] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_116 
+ bl[114] br[114] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_117 
+ bl[115] br[115] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_118 
+ bl[116] br[116] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_119 
+ bl[117] br[117] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_120 
+ bl[118] br[118] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_121 
+ bl[119] br[119] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_122 
+ bl[120] br[120] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_123 
+ bl[121] br[121] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_124 
+ bl[122] br[122] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_125 
+ bl[123] br[123] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_126 
+ bl[124] br[124] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_127 
+ bl[125] br[125] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_128 
+ bl[126] br[126] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_129 
+ bl[127] br[127] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_130 
+ bl[128] br[128] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_131 
+ bl[129] br[129] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_132 
+ bl[130] br[130] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_133 
+ bl[131] br[131] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_134 
+ bl[132] br[132] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_135 
+ bl[133] br[133] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_136 
+ bl[134] br[134] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_137 
+ bl[135] br[135] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_138 
+ bl[136] br[136] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_139 
+ bl[137] br[137] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_140 
+ bl[138] br[138] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_141 
+ bl[139] br[139] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_142 
+ bl[140] br[140] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_143 
+ bl[141] br[141] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_144 
+ bl[142] br[142] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_145 
+ bl[143] br[143] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_146 
+ bl[144] br[144] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_147 
+ bl[145] br[145] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_148 
+ bl[146] br[146] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_149 
+ bl[147] br[147] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_150 
+ bl[148] br[148] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_151 
+ bl[149] br[149] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_152 
+ bl[150] br[150] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_153 
+ bl[151] br[151] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_154 
+ bl[152] br[152] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_155 
+ bl[153] br[153] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_156 
+ bl[154] br[154] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_157 
+ bl[155] br[155] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_158 
+ bl[156] br[156] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_159 
+ bl[157] br[157] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_160 
+ bl[158] br[158] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_161 
+ bl[159] br[159] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_162 
+ bl[160] br[160] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_163 
+ bl[161] br[161] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_164 
+ bl[162] br[162] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_165 
+ bl[163] br[163] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_166 
+ bl[164] br[164] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_167 
+ bl[165] br[165] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_168 
+ bl[166] br[166] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_169 
+ bl[167] br[167] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_170 
+ bl[168] br[168] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_171 
+ bl[169] br[169] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_172 
+ bl[170] br[170] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_173 
+ bl[171] br[171] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_174 
+ bl[172] br[172] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_175 
+ bl[173] br[173] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_176 
+ bl[174] br[174] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_177 
+ bl[175] br[175] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_178 
+ bl[176] br[176] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_179 
+ bl[177] br[177] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_180 
+ bl[178] br[178] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_181 
+ bl[179] br[179] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_182 
+ bl[180] br[180] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_183 
+ bl[181] br[181] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_184 
+ bl[182] br[182] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_185 
+ bl[183] br[183] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_186 
+ bl[184] br[184] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_187 
+ bl[185] br[185] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_188 
+ bl[186] br[186] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_189 
+ bl[187] br[187] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_190 
+ bl[188] br[188] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_191 
+ bl[189] br[189] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_192 
+ bl[190] br[190] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_193 
+ bl[191] br[191] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_194 
+ bl[192] br[192] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_195 
+ bl[193] br[193] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_196 
+ bl[194] br[194] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_197 
+ bl[195] br[195] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_198 
+ bl[196] br[196] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_199 
+ bl[197] br[197] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_200 
+ bl[198] br[198] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_201 
+ bl[199] br[199] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_202 
+ bl[200] br[200] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_203 
+ bl[201] br[201] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_204 
+ bl[202] br[202] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_205 
+ bl[203] br[203] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_206 
+ bl[204] br[204] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_207 
+ bl[205] br[205] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_208 
+ bl[206] br[206] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_209 
+ bl[207] br[207] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_210 
+ bl[208] br[208] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_211 
+ bl[209] br[209] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_212 
+ bl[210] br[210] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_213 
+ bl[211] br[211] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_214 
+ bl[212] br[212] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_215 
+ bl[213] br[213] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_216 
+ bl[214] br[214] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_217 
+ bl[215] br[215] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_218 
+ bl[216] br[216] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_219 
+ bl[217] br[217] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_220 
+ bl[218] br[218] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_221 
+ bl[219] br[219] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_222 
+ bl[220] br[220] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_223 
+ bl[221] br[221] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_224 
+ bl[222] br[222] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_225 
+ bl[223] br[223] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_226 
+ bl[224] br[224] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_227 
+ bl[225] br[225] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_228 
+ bl[226] br[226] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_229 
+ bl[227] br[227] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_230 
+ bl[228] br[228] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_231 
+ bl[229] br[229] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_232 
+ bl[230] br[230] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_233 
+ bl[231] br[231] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_234 
+ bl[232] br[232] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_235 
+ bl[233] br[233] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_236 
+ bl[234] br[234] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_237 
+ bl[235] br[235] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_238 
+ bl[236] br[236] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_239 
+ bl[237] br[237] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_240 
+ bl[238] br[238] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_241 
+ bl[239] br[239] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_242 
+ bl[240] br[240] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_243 
+ bl[241] br[241] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_244 
+ bl[242] br[242] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_245 
+ bl[243] br[243] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_246 
+ bl[244] br[244] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_247 
+ bl[245] br[245] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_248 
+ bl[246] br[246] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_249 
+ bl[247] br[247] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_250 
+ bl[248] br[248] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_251 
+ bl[249] br[249] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_252 
+ bl[250] br[250] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_253 
+ bl[251] br[251] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_254 
+ bl[252] br[252] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_255 
+ bl[253] br[253] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_256 
+ bl[254] br[254] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_257 
+ bl[255] br[255] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_258 
+ vdd vdd vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_259 
+ vdd vdd vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_0 
+ vdd vdd vss vdd vpb vnb wl[13] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_15_1 
+ rbl rbr vss vdd vpb vnb wl[13] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_15_2 
+ bl[0] br[0] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_3 
+ bl[1] br[1] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_4 
+ bl[2] br[2] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_5 
+ bl[3] br[3] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_6 
+ bl[4] br[4] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_7 
+ bl[5] br[5] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_8 
+ bl[6] br[6] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_9 
+ bl[7] br[7] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_10 
+ bl[8] br[8] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_11 
+ bl[9] br[9] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_12 
+ bl[10] br[10] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_13 
+ bl[11] br[11] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_14 
+ bl[12] br[12] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_15 
+ bl[13] br[13] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_16 
+ bl[14] br[14] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_17 
+ bl[15] br[15] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_18 
+ bl[16] br[16] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_19 
+ bl[17] br[17] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_20 
+ bl[18] br[18] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_21 
+ bl[19] br[19] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_22 
+ bl[20] br[20] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_23 
+ bl[21] br[21] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_24 
+ bl[22] br[22] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_25 
+ bl[23] br[23] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_26 
+ bl[24] br[24] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_27 
+ bl[25] br[25] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_28 
+ bl[26] br[26] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_29 
+ bl[27] br[27] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_30 
+ bl[28] br[28] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_31 
+ bl[29] br[29] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_32 
+ bl[30] br[30] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_33 
+ bl[31] br[31] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_34 
+ bl[32] br[32] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_35 
+ bl[33] br[33] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_36 
+ bl[34] br[34] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_37 
+ bl[35] br[35] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_38 
+ bl[36] br[36] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_39 
+ bl[37] br[37] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_40 
+ bl[38] br[38] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_41 
+ bl[39] br[39] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_42 
+ bl[40] br[40] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_43 
+ bl[41] br[41] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_44 
+ bl[42] br[42] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_45 
+ bl[43] br[43] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_46 
+ bl[44] br[44] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_47 
+ bl[45] br[45] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_48 
+ bl[46] br[46] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_49 
+ bl[47] br[47] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_50 
+ bl[48] br[48] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_51 
+ bl[49] br[49] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_52 
+ bl[50] br[50] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_53 
+ bl[51] br[51] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_54 
+ bl[52] br[52] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_55 
+ bl[53] br[53] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_56 
+ bl[54] br[54] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_57 
+ bl[55] br[55] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_58 
+ bl[56] br[56] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_59 
+ bl[57] br[57] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_60 
+ bl[58] br[58] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_61 
+ bl[59] br[59] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_62 
+ bl[60] br[60] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_63 
+ bl[61] br[61] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_64 
+ bl[62] br[62] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_65 
+ bl[63] br[63] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_66 
+ bl[64] br[64] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_67 
+ bl[65] br[65] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_68 
+ bl[66] br[66] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_69 
+ bl[67] br[67] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_70 
+ bl[68] br[68] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_71 
+ bl[69] br[69] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_72 
+ bl[70] br[70] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_73 
+ bl[71] br[71] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_74 
+ bl[72] br[72] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_75 
+ bl[73] br[73] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_76 
+ bl[74] br[74] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_77 
+ bl[75] br[75] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_78 
+ bl[76] br[76] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_79 
+ bl[77] br[77] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_80 
+ bl[78] br[78] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_81 
+ bl[79] br[79] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_82 
+ bl[80] br[80] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_83 
+ bl[81] br[81] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_84 
+ bl[82] br[82] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_85 
+ bl[83] br[83] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_86 
+ bl[84] br[84] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_87 
+ bl[85] br[85] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_88 
+ bl[86] br[86] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_89 
+ bl[87] br[87] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_90 
+ bl[88] br[88] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_91 
+ bl[89] br[89] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_92 
+ bl[90] br[90] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_93 
+ bl[91] br[91] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_94 
+ bl[92] br[92] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_95 
+ bl[93] br[93] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_96 
+ bl[94] br[94] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_97 
+ bl[95] br[95] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_98 
+ bl[96] br[96] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_99 
+ bl[97] br[97] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_100 
+ bl[98] br[98] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_101 
+ bl[99] br[99] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_102 
+ bl[100] br[100] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_103 
+ bl[101] br[101] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_104 
+ bl[102] br[102] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_105 
+ bl[103] br[103] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_106 
+ bl[104] br[104] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_107 
+ bl[105] br[105] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_108 
+ bl[106] br[106] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_109 
+ bl[107] br[107] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_110 
+ bl[108] br[108] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_111 
+ bl[109] br[109] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_112 
+ bl[110] br[110] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_113 
+ bl[111] br[111] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_114 
+ bl[112] br[112] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_115 
+ bl[113] br[113] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_116 
+ bl[114] br[114] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_117 
+ bl[115] br[115] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_118 
+ bl[116] br[116] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_119 
+ bl[117] br[117] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_120 
+ bl[118] br[118] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_121 
+ bl[119] br[119] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_122 
+ bl[120] br[120] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_123 
+ bl[121] br[121] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_124 
+ bl[122] br[122] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_125 
+ bl[123] br[123] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_126 
+ bl[124] br[124] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_127 
+ bl[125] br[125] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_128 
+ bl[126] br[126] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_129 
+ bl[127] br[127] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_130 
+ bl[128] br[128] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_131 
+ bl[129] br[129] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_132 
+ bl[130] br[130] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_133 
+ bl[131] br[131] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_134 
+ bl[132] br[132] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_135 
+ bl[133] br[133] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_136 
+ bl[134] br[134] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_137 
+ bl[135] br[135] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_138 
+ bl[136] br[136] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_139 
+ bl[137] br[137] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_140 
+ bl[138] br[138] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_141 
+ bl[139] br[139] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_142 
+ bl[140] br[140] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_143 
+ bl[141] br[141] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_144 
+ bl[142] br[142] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_145 
+ bl[143] br[143] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_146 
+ bl[144] br[144] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_147 
+ bl[145] br[145] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_148 
+ bl[146] br[146] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_149 
+ bl[147] br[147] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_150 
+ bl[148] br[148] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_151 
+ bl[149] br[149] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_152 
+ bl[150] br[150] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_153 
+ bl[151] br[151] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_154 
+ bl[152] br[152] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_155 
+ bl[153] br[153] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_156 
+ bl[154] br[154] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_157 
+ bl[155] br[155] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_158 
+ bl[156] br[156] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_159 
+ bl[157] br[157] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_160 
+ bl[158] br[158] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_161 
+ bl[159] br[159] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_162 
+ bl[160] br[160] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_163 
+ bl[161] br[161] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_164 
+ bl[162] br[162] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_165 
+ bl[163] br[163] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_166 
+ bl[164] br[164] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_167 
+ bl[165] br[165] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_168 
+ bl[166] br[166] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_169 
+ bl[167] br[167] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_170 
+ bl[168] br[168] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_171 
+ bl[169] br[169] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_172 
+ bl[170] br[170] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_173 
+ bl[171] br[171] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_174 
+ bl[172] br[172] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_175 
+ bl[173] br[173] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_176 
+ bl[174] br[174] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_177 
+ bl[175] br[175] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_178 
+ bl[176] br[176] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_179 
+ bl[177] br[177] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_180 
+ bl[178] br[178] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_181 
+ bl[179] br[179] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_182 
+ bl[180] br[180] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_183 
+ bl[181] br[181] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_184 
+ bl[182] br[182] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_185 
+ bl[183] br[183] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_186 
+ bl[184] br[184] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_187 
+ bl[185] br[185] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_188 
+ bl[186] br[186] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_189 
+ bl[187] br[187] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_190 
+ bl[188] br[188] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_191 
+ bl[189] br[189] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_192 
+ bl[190] br[190] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_193 
+ bl[191] br[191] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_194 
+ bl[192] br[192] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_195 
+ bl[193] br[193] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_196 
+ bl[194] br[194] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_197 
+ bl[195] br[195] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_198 
+ bl[196] br[196] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_199 
+ bl[197] br[197] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_200 
+ bl[198] br[198] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_201 
+ bl[199] br[199] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_202 
+ bl[200] br[200] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_203 
+ bl[201] br[201] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_204 
+ bl[202] br[202] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_205 
+ bl[203] br[203] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_206 
+ bl[204] br[204] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_207 
+ bl[205] br[205] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_208 
+ bl[206] br[206] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_209 
+ bl[207] br[207] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_210 
+ bl[208] br[208] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_211 
+ bl[209] br[209] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_212 
+ bl[210] br[210] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_213 
+ bl[211] br[211] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_214 
+ bl[212] br[212] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_215 
+ bl[213] br[213] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_216 
+ bl[214] br[214] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_217 
+ bl[215] br[215] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_218 
+ bl[216] br[216] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_219 
+ bl[217] br[217] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_220 
+ bl[218] br[218] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_221 
+ bl[219] br[219] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_222 
+ bl[220] br[220] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_223 
+ bl[221] br[221] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_224 
+ bl[222] br[222] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_225 
+ bl[223] br[223] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_226 
+ bl[224] br[224] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_227 
+ bl[225] br[225] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_228 
+ bl[226] br[226] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_229 
+ bl[227] br[227] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_230 
+ bl[228] br[228] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_231 
+ bl[229] br[229] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_232 
+ bl[230] br[230] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_233 
+ bl[231] br[231] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_234 
+ bl[232] br[232] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_235 
+ bl[233] br[233] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_236 
+ bl[234] br[234] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_237 
+ bl[235] br[235] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_238 
+ bl[236] br[236] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_239 
+ bl[237] br[237] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_240 
+ bl[238] br[238] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_241 
+ bl[239] br[239] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_242 
+ bl[240] br[240] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_243 
+ bl[241] br[241] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_244 
+ bl[242] br[242] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_245 
+ bl[243] br[243] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_246 
+ bl[244] br[244] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_247 
+ bl[245] br[245] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_248 
+ bl[246] br[246] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_249 
+ bl[247] br[247] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_250 
+ bl[248] br[248] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_251 
+ bl[249] br[249] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_252 
+ bl[250] br[250] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_253 
+ bl[251] br[251] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_254 
+ bl[252] br[252] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_255 
+ bl[253] br[253] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_256 
+ bl[254] br[254] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_257 
+ bl[255] br[255] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_258 
+ vdd vdd vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_259 
+ vdd vdd vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_0 
+ vdd vdd vss vdd vpb vnb wl[14] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_16_1 
+ rbl rbr vss vdd vpb vnb wl[14] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_16_2 
+ bl[0] br[0] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_3 
+ bl[1] br[1] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_4 
+ bl[2] br[2] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_5 
+ bl[3] br[3] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_6 
+ bl[4] br[4] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_7 
+ bl[5] br[5] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_8 
+ bl[6] br[6] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_9 
+ bl[7] br[7] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_10 
+ bl[8] br[8] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_11 
+ bl[9] br[9] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_12 
+ bl[10] br[10] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_13 
+ bl[11] br[11] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_14 
+ bl[12] br[12] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_15 
+ bl[13] br[13] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_16 
+ bl[14] br[14] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_17 
+ bl[15] br[15] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_18 
+ bl[16] br[16] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_19 
+ bl[17] br[17] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_20 
+ bl[18] br[18] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_21 
+ bl[19] br[19] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_22 
+ bl[20] br[20] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_23 
+ bl[21] br[21] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_24 
+ bl[22] br[22] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_25 
+ bl[23] br[23] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_26 
+ bl[24] br[24] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_27 
+ bl[25] br[25] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_28 
+ bl[26] br[26] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_29 
+ bl[27] br[27] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_30 
+ bl[28] br[28] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_31 
+ bl[29] br[29] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_32 
+ bl[30] br[30] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_33 
+ bl[31] br[31] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_34 
+ bl[32] br[32] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_35 
+ bl[33] br[33] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_36 
+ bl[34] br[34] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_37 
+ bl[35] br[35] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_38 
+ bl[36] br[36] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_39 
+ bl[37] br[37] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_40 
+ bl[38] br[38] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_41 
+ bl[39] br[39] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_42 
+ bl[40] br[40] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_43 
+ bl[41] br[41] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_44 
+ bl[42] br[42] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_45 
+ bl[43] br[43] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_46 
+ bl[44] br[44] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_47 
+ bl[45] br[45] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_48 
+ bl[46] br[46] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_49 
+ bl[47] br[47] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_50 
+ bl[48] br[48] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_51 
+ bl[49] br[49] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_52 
+ bl[50] br[50] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_53 
+ bl[51] br[51] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_54 
+ bl[52] br[52] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_55 
+ bl[53] br[53] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_56 
+ bl[54] br[54] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_57 
+ bl[55] br[55] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_58 
+ bl[56] br[56] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_59 
+ bl[57] br[57] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_60 
+ bl[58] br[58] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_61 
+ bl[59] br[59] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_62 
+ bl[60] br[60] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_63 
+ bl[61] br[61] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_64 
+ bl[62] br[62] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_65 
+ bl[63] br[63] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_66 
+ bl[64] br[64] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_67 
+ bl[65] br[65] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_68 
+ bl[66] br[66] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_69 
+ bl[67] br[67] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_70 
+ bl[68] br[68] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_71 
+ bl[69] br[69] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_72 
+ bl[70] br[70] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_73 
+ bl[71] br[71] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_74 
+ bl[72] br[72] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_75 
+ bl[73] br[73] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_76 
+ bl[74] br[74] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_77 
+ bl[75] br[75] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_78 
+ bl[76] br[76] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_79 
+ bl[77] br[77] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_80 
+ bl[78] br[78] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_81 
+ bl[79] br[79] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_82 
+ bl[80] br[80] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_83 
+ bl[81] br[81] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_84 
+ bl[82] br[82] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_85 
+ bl[83] br[83] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_86 
+ bl[84] br[84] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_87 
+ bl[85] br[85] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_88 
+ bl[86] br[86] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_89 
+ bl[87] br[87] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_90 
+ bl[88] br[88] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_91 
+ bl[89] br[89] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_92 
+ bl[90] br[90] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_93 
+ bl[91] br[91] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_94 
+ bl[92] br[92] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_95 
+ bl[93] br[93] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_96 
+ bl[94] br[94] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_97 
+ bl[95] br[95] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_98 
+ bl[96] br[96] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_99 
+ bl[97] br[97] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_100 
+ bl[98] br[98] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_101 
+ bl[99] br[99] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_102 
+ bl[100] br[100] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_103 
+ bl[101] br[101] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_104 
+ bl[102] br[102] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_105 
+ bl[103] br[103] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_106 
+ bl[104] br[104] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_107 
+ bl[105] br[105] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_108 
+ bl[106] br[106] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_109 
+ bl[107] br[107] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_110 
+ bl[108] br[108] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_111 
+ bl[109] br[109] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_112 
+ bl[110] br[110] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_113 
+ bl[111] br[111] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_114 
+ bl[112] br[112] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_115 
+ bl[113] br[113] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_116 
+ bl[114] br[114] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_117 
+ bl[115] br[115] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_118 
+ bl[116] br[116] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_119 
+ bl[117] br[117] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_120 
+ bl[118] br[118] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_121 
+ bl[119] br[119] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_122 
+ bl[120] br[120] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_123 
+ bl[121] br[121] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_124 
+ bl[122] br[122] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_125 
+ bl[123] br[123] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_126 
+ bl[124] br[124] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_127 
+ bl[125] br[125] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_128 
+ bl[126] br[126] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_129 
+ bl[127] br[127] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_130 
+ bl[128] br[128] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_131 
+ bl[129] br[129] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_132 
+ bl[130] br[130] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_133 
+ bl[131] br[131] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_134 
+ bl[132] br[132] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_135 
+ bl[133] br[133] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_136 
+ bl[134] br[134] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_137 
+ bl[135] br[135] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_138 
+ bl[136] br[136] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_139 
+ bl[137] br[137] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_140 
+ bl[138] br[138] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_141 
+ bl[139] br[139] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_142 
+ bl[140] br[140] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_143 
+ bl[141] br[141] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_144 
+ bl[142] br[142] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_145 
+ bl[143] br[143] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_146 
+ bl[144] br[144] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_147 
+ bl[145] br[145] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_148 
+ bl[146] br[146] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_149 
+ bl[147] br[147] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_150 
+ bl[148] br[148] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_151 
+ bl[149] br[149] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_152 
+ bl[150] br[150] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_153 
+ bl[151] br[151] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_154 
+ bl[152] br[152] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_155 
+ bl[153] br[153] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_156 
+ bl[154] br[154] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_157 
+ bl[155] br[155] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_158 
+ bl[156] br[156] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_159 
+ bl[157] br[157] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_160 
+ bl[158] br[158] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_161 
+ bl[159] br[159] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_162 
+ bl[160] br[160] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_163 
+ bl[161] br[161] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_164 
+ bl[162] br[162] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_165 
+ bl[163] br[163] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_166 
+ bl[164] br[164] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_167 
+ bl[165] br[165] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_168 
+ bl[166] br[166] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_169 
+ bl[167] br[167] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_170 
+ bl[168] br[168] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_171 
+ bl[169] br[169] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_172 
+ bl[170] br[170] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_173 
+ bl[171] br[171] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_174 
+ bl[172] br[172] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_175 
+ bl[173] br[173] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_176 
+ bl[174] br[174] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_177 
+ bl[175] br[175] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_178 
+ bl[176] br[176] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_179 
+ bl[177] br[177] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_180 
+ bl[178] br[178] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_181 
+ bl[179] br[179] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_182 
+ bl[180] br[180] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_183 
+ bl[181] br[181] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_184 
+ bl[182] br[182] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_185 
+ bl[183] br[183] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_186 
+ bl[184] br[184] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_187 
+ bl[185] br[185] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_188 
+ bl[186] br[186] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_189 
+ bl[187] br[187] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_190 
+ bl[188] br[188] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_191 
+ bl[189] br[189] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_192 
+ bl[190] br[190] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_193 
+ bl[191] br[191] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_194 
+ bl[192] br[192] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_195 
+ bl[193] br[193] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_196 
+ bl[194] br[194] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_197 
+ bl[195] br[195] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_198 
+ bl[196] br[196] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_199 
+ bl[197] br[197] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_200 
+ bl[198] br[198] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_201 
+ bl[199] br[199] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_202 
+ bl[200] br[200] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_203 
+ bl[201] br[201] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_204 
+ bl[202] br[202] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_205 
+ bl[203] br[203] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_206 
+ bl[204] br[204] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_207 
+ bl[205] br[205] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_208 
+ bl[206] br[206] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_209 
+ bl[207] br[207] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_210 
+ bl[208] br[208] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_211 
+ bl[209] br[209] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_212 
+ bl[210] br[210] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_213 
+ bl[211] br[211] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_214 
+ bl[212] br[212] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_215 
+ bl[213] br[213] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_216 
+ bl[214] br[214] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_217 
+ bl[215] br[215] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_218 
+ bl[216] br[216] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_219 
+ bl[217] br[217] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_220 
+ bl[218] br[218] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_221 
+ bl[219] br[219] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_222 
+ bl[220] br[220] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_223 
+ bl[221] br[221] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_224 
+ bl[222] br[222] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_225 
+ bl[223] br[223] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_226 
+ bl[224] br[224] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_227 
+ bl[225] br[225] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_228 
+ bl[226] br[226] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_229 
+ bl[227] br[227] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_230 
+ bl[228] br[228] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_231 
+ bl[229] br[229] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_232 
+ bl[230] br[230] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_233 
+ bl[231] br[231] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_234 
+ bl[232] br[232] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_235 
+ bl[233] br[233] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_236 
+ bl[234] br[234] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_237 
+ bl[235] br[235] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_238 
+ bl[236] br[236] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_239 
+ bl[237] br[237] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_240 
+ bl[238] br[238] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_241 
+ bl[239] br[239] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_242 
+ bl[240] br[240] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_243 
+ bl[241] br[241] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_244 
+ bl[242] br[242] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_245 
+ bl[243] br[243] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_246 
+ bl[244] br[244] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_247 
+ bl[245] br[245] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_248 
+ bl[246] br[246] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_249 
+ bl[247] br[247] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_250 
+ bl[248] br[248] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_251 
+ bl[249] br[249] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_252 
+ bl[250] br[250] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_253 
+ bl[251] br[251] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_254 
+ bl[252] br[252] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_255 
+ bl[253] br[253] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_256 
+ bl[254] br[254] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_257 
+ bl[255] br[255] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_258 
+ vdd vdd vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_259 
+ vdd vdd vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_0 
+ vdd vdd vss vdd vpb vnb wl[15] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_17_1 
+ rbl rbr vss vdd vpb vnb wl[15] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_17_2 
+ bl[0] br[0] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_3 
+ bl[1] br[1] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_4 
+ bl[2] br[2] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_5 
+ bl[3] br[3] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_6 
+ bl[4] br[4] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_7 
+ bl[5] br[5] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_8 
+ bl[6] br[6] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_9 
+ bl[7] br[7] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_10 
+ bl[8] br[8] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_11 
+ bl[9] br[9] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_12 
+ bl[10] br[10] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_13 
+ bl[11] br[11] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_14 
+ bl[12] br[12] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_15 
+ bl[13] br[13] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_16 
+ bl[14] br[14] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_17 
+ bl[15] br[15] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_18 
+ bl[16] br[16] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_19 
+ bl[17] br[17] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_20 
+ bl[18] br[18] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_21 
+ bl[19] br[19] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_22 
+ bl[20] br[20] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_23 
+ bl[21] br[21] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_24 
+ bl[22] br[22] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_25 
+ bl[23] br[23] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_26 
+ bl[24] br[24] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_27 
+ bl[25] br[25] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_28 
+ bl[26] br[26] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_29 
+ bl[27] br[27] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_30 
+ bl[28] br[28] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_31 
+ bl[29] br[29] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_32 
+ bl[30] br[30] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_33 
+ bl[31] br[31] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_34 
+ bl[32] br[32] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_35 
+ bl[33] br[33] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_36 
+ bl[34] br[34] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_37 
+ bl[35] br[35] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_38 
+ bl[36] br[36] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_39 
+ bl[37] br[37] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_40 
+ bl[38] br[38] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_41 
+ bl[39] br[39] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_42 
+ bl[40] br[40] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_43 
+ bl[41] br[41] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_44 
+ bl[42] br[42] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_45 
+ bl[43] br[43] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_46 
+ bl[44] br[44] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_47 
+ bl[45] br[45] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_48 
+ bl[46] br[46] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_49 
+ bl[47] br[47] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_50 
+ bl[48] br[48] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_51 
+ bl[49] br[49] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_52 
+ bl[50] br[50] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_53 
+ bl[51] br[51] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_54 
+ bl[52] br[52] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_55 
+ bl[53] br[53] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_56 
+ bl[54] br[54] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_57 
+ bl[55] br[55] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_58 
+ bl[56] br[56] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_59 
+ bl[57] br[57] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_60 
+ bl[58] br[58] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_61 
+ bl[59] br[59] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_62 
+ bl[60] br[60] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_63 
+ bl[61] br[61] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_64 
+ bl[62] br[62] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_65 
+ bl[63] br[63] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_66 
+ bl[64] br[64] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_67 
+ bl[65] br[65] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_68 
+ bl[66] br[66] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_69 
+ bl[67] br[67] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_70 
+ bl[68] br[68] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_71 
+ bl[69] br[69] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_72 
+ bl[70] br[70] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_73 
+ bl[71] br[71] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_74 
+ bl[72] br[72] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_75 
+ bl[73] br[73] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_76 
+ bl[74] br[74] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_77 
+ bl[75] br[75] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_78 
+ bl[76] br[76] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_79 
+ bl[77] br[77] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_80 
+ bl[78] br[78] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_81 
+ bl[79] br[79] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_82 
+ bl[80] br[80] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_83 
+ bl[81] br[81] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_84 
+ bl[82] br[82] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_85 
+ bl[83] br[83] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_86 
+ bl[84] br[84] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_87 
+ bl[85] br[85] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_88 
+ bl[86] br[86] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_89 
+ bl[87] br[87] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_90 
+ bl[88] br[88] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_91 
+ bl[89] br[89] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_92 
+ bl[90] br[90] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_93 
+ bl[91] br[91] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_94 
+ bl[92] br[92] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_95 
+ bl[93] br[93] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_96 
+ bl[94] br[94] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_97 
+ bl[95] br[95] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_98 
+ bl[96] br[96] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_99 
+ bl[97] br[97] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_100 
+ bl[98] br[98] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_101 
+ bl[99] br[99] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_102 
+ bl[100] br[100] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_103 
+ bl[101] br[101] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_104 
+ bl[102] br[102] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_105 
+ bl[103] br[103] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_106 
+ bl[104] br[104] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_107 
+ bl[105] br[105] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_108 
+ bl[106] br[106] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_109 
+ bl[107] br[107] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_110 
+ bl[108] br[108] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_111 
+ bl[109] br[109] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_112 
+ bl[110] br[110] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_113 
+ bl[111] br[111] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_114 
+ bl[112] br[112] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_115 
+ bl[113] br[113] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_116 
+ bl[114] br[114] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_117 
+ bl[115] br[115] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_118 
+ bl[116] br[116] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_119 
+ bl[117] br[117] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_120 
+ bl[118] br[118] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_121 
+ bl[119] br[119] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_122 
+ bl[120] br[120] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_123 
+ bl[121] br[121] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_124 
+ bl[122] br[122] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_125 
+ bl[123] br[123] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_126 
+ bl[124] br[124] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_127 
+ bl[125] br[125] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_128 
+ bl[126] br[126] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_129 
+ bl[127] br[127] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_130 
+ bl[128] br[128] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_131 
+ bl[129] br[129] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_132 
+ bl[130] br[130] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_133 
+ bl[131] br[131] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_134 
+ bl[132] br[132] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_135 
+ bl[133] br[133] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_136 
+ bl[134] br[134] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_137 
+ bl[135] br[135] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_138 
+ bl[136] br[136] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_139 
+ bl[137] br[137] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_140 
+ bl[138] br[138] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_141 
+ bl[139] br[139] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_142 
+ bl[140] br[140] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_143 
+ bl[141] br[141] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_144 
+ bl[142] br[142] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_145 
+ bl[143] br[143] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_146 
+ bl[144] br[144] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_147 
+ bl[145] br[145] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_148 
+ bl[146] br[146] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_149 
+ bl[147] br[147] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_150 
+ bl[148] br[148] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_151 
+ bl[149] br[149] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_152 
+ bl[150] br[150] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_153 
+ bl[151] br[151] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_154 
+ bl[152] br[152] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_155 
+ bl[153] br[153] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_156 
+ bl[154] br[154] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_157 
+ bl[155] br[155] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_158 
+ bl[156] br[156] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_159 
+ bl[157] br[157] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_160 
+ bl[158] br[158] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_161 
+ bl[159] br[159] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_162 
+ bl[160] br[160] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_163 
+ bl[161] br[161] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_164 
+ bl[162] br[162] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_165 
+ bl[163] br[163] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_166 
+ bl[164] br[164] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_167 
+ bl[165] br[165] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_168 
+ bl[166] br[166] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_169 
+ bl[167] br[167] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_170 
+ bl[168] br[168] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_171 
+ bl[169] br[169] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_172 
+ bl[170] br[170] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_173 
+ bl[171] br[171] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_174 
+ bl[172] br[172] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_175 
+ bl[173] br[173] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_176 
+ bl[174] br[174] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_177 
+ bl[175] br[175] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_178 
+ bl[176] br[176] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_179 
+ bl[177] br[177] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_180 
+ bl[178] br[178] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_181 
+ bl[179] br[179] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_182 
+ bl[180] br[180] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_183 
+ bl[181] br[181] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_184 
+ bl[182] br[182] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_185 
+ bl[183] br[183] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_186 
+ bl[184] br[184] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_187 
+ bl[185] br[185] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_188 
+ bl[186] br[186] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_189 
+ bl[187] br[187] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_190 
+ bl[188] br[188] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_191 
+ bl[189] br[189] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_192 
+ bl[190] br[190] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_193 
+ bl[191] br[191] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_194 
+ bl[192] br[192] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_195 
+ bl[193] br[193] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_196 
+ bl[194] br[194] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_197 
+ bl[195] br[195] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_198 
+ bl[196] br[196] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_199 
+ bl[197] br[197] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_200 
+ bl[198] br[198] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_201 
+ bl[199] br[199] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_202 
+ bl[200] br[200] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_203 
+ bl[201] br[201] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_204 
+ bl[202] br[202] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_205 
+ bl[203] br[203] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_206 
+ bl[204] br[204] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_207 
+ bl[205] br[205] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_208 
+ bl[206] br[206] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_209 
+ bl[207] br[207] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_210 
+ bl[208] br[208] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_211 
+ bl[209] br[209] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_212 
+ bl[210] br[210] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_213 
+ bl[211] br[211] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_214 
+ bl[212] br[212] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_215 
+ bl[213] br[213] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_216 
+ bl[214] br[214] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_217 
+ bl[215] br[215] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_218 
+ bl[216] br[216] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_219 
+ bl[217] br[217] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_220 
+ bl[218] br[218] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_221 
+ bl[219] br[219] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_222 
+ bl[220] br[220] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_223 
+ bl[221] br[221] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_224 
+ bl[222] br[222] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_225 
+ bl[223] br[223] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_226 
+ bl[224] br[224] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_227 
+ bl[225] br[225] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_228 
+ bl[226] br[226] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_229 
+ bl[227] br[227] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_230 
+ bl[228] br[228] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_231 
+ bl[229] br[229] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_232 
+ bl[230] br[230] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_233 
+ bl[231] br[231] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_234 
+ bl[232] br[232] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_235 
+ bl[233] br[233] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_236 
+ bl[234] br[234] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_237 
+ bl[235] br[235] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_238 
+ bl[236] br[236] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_239 
+ bl[237] br[237] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_240 
+ bl[238] br[238] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_241 
+ bl[239] br[239] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_242 
+ bl[240] br[240] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_243 
+ bl[241] br[241] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_244 
+ bl[242] br[242] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_245 
+ bl[243] br[243] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_246 
+ bl[244] br[244] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_247 
+ bl[245] br[245] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_248 
+ bl[246] br[246] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_249 
+ bl[247] br[247] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_250 
+ bl[248] br[248] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_251 
+ bl[249] br[249] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_252 
+ bl[250] br[250] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_253 
+ bl[251] br[251] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_254 
+ bl[252] br[252] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_255 
+ bl[253] br[253] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_256 
+ bl[254] br[254] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_257 
+ bl[255] br[255] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_258 
+ vdd vdd vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_259 
+ vdd vdd vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_0 
+ vdd vdd vss vdd vpb vnb wl[16] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_18_1 
+ rbl rbr vss vdd vpb vnb wl[16] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_18_2 
+ bl[0] br[0] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_3 
+ bl[1] br[1] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_4 
+ bl[2] br[2] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_5 
+ bl[3] br[3] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_6 
+ bl[4] br[4] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_7 
+ bl[5] br[5] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_8 
+ bl[6] br[6] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_9 
+ bl[7] br[7] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_10 
+ bl[8] br[8] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_11 
+ bl[9] br[9] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_12 
+ bl[10] br[10] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_13 
+ bl[11] br[11] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_14 
+ bl[12] br[12] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_15 
+ bl[13] br[13] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_16 
+ bl[14] br[14] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_17 
+ bl[15] br[15] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_18 
+ bl[16] br[16] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_19 
+ bl[17] br[17] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_20 
+ bl[18] br[18] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_21 
+ bl[19] br[19] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_22 
+ bl[20] br[20] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_23 
+ bl[21] br[21] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_24 
+ bl[22] br[22] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_25 
+ bl[23] br[23] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_26 
+ bl[24] br[24] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_27 
+ bl[25] br[25] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_28 
+ bl[26] br[26] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_29 
+ bl[27] br[27] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_30 
+ bl[28] br[28] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_31 
+ bl[29] br[29] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_32 
+ bl[30] br[30] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_33 
+ bl[31] br[31] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_34 
+ bl[32] br[32] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_35 
+ bl[33] br[33] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_36 
+ bl[34] br[34] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_37 
+ bl[35] br[35] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_38 
+ bl[36] br[36] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_39 
+ bl[37] br[37] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_40 
+ bl[38] br[38] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_41 
+ bl[39] br[39] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_42 
+ bl[40] br[40] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_43 
+ bl[41] br[41] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_44 
+ bl[42] br[42] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_45 
+ bl[43] br[43] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_46 
+ bl[44] br[44] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_47 
+ bl[45] br[45] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_48 
+ bl[46] br[46] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_49 
+ bl[47] br[47] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_50 
+ bl[48] br[48] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_51 
+ bl[49] br[49] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_52 
+ bl[50] br[50] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_53 
+ bl[51] br[51] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_54 
+ bl[52] br[52] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_55 
+ bl[53] br[53] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_56 
+ bl[54] br[54] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_57 
+ bl[55] br[55] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_58 
+ bl[56] br[56] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_59 
+ bl[57] br[57] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_60 
+ bl[58] br[58] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_61 
+ bl[59] br[59] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_62 
+ bl[60] br[60] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_63 
+ bl[61] br[61] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_64 
+ bl[62] br[62] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_65 
+ bl[63] br[63] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_66 
+ bl[64] br[64] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_67 
+ bl[65] br[65] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_68 
+ bl[66] br[66] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_69 
+ bl[67] br[67] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_70 
+ bl[68] br[68] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_71 
+ bl[69] br[69] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_72 
+ bl[70] br[70] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_73 
+ bl[71] br[71] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_74 
+ bl[72] br[72] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_75 
+ bl[73] br[73] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_76 
+ bl[74] br[74] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_77 
+ bl[75] br[75] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_78 
+ bl[76] br[76] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_79 
+ bl[77] br[77] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_80 
+ bl[78] br[78] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_81 
+ bl[79] br[79] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_82 
+ bl[80] br[80] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_83 
+ bl[81] br[81] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_84 
+ bl[82] br[82] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_85 
+ bl[83] br[83] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_86 
+ bl[84] br[84] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_87 
+ bl[85] br[85] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_88 
+ bl[86] br[86] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_89 
+ bl[87] br[87] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_90 
+ bl[88] br[88] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_91 
+ bl[89] br[89] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_92 
+ bl[90] br[90] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_93 
+ bl[91] br[91] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_94 
+ bl[92] br[92] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_95 
+ bl[93] br[93] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_96 
+ bl[94] br[94] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_97 
+ bl[95] br[95] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_98 
+ bl[96] br[96] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_99 
+ bl[97] br[97] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_100 
+ bl[98] br[98] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_101 
+ bl[99] br[99] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_102 
+ bl[100] br[100] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_103 
+ bl[101] br[101] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_104 
+ bl[102] br[102] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_105 
+ bl[103] br[103] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_106 
+ bl[104] br[104] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_107 
+ bl[105] br[105] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_108 
+ bl[106] br[106] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_109 
+ bl[107] br[107] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_110 
+ bl[108] br[108] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_111 
+ bl[109] br[109] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_112 
+ bl[110] br[110] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_113 
+ bl[111] br[111] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_114 
+ bl[112] br[112] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_115 
+ bl[113] br[113] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_116 
+ bl[114] br[114] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_117 
+ bl[115] br[115] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_118 
+ bl[116] br[116] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_119 
+ bl[117] br[117] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_120 
+ bl[118] br[118] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_121 
+ bl[119] br[119] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_122 
+ bl[120] br[120] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_123 
+ bl[121] br[121] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_124 
+ bl[122] br[122] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_125 
+ bl[123] br[123] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_126 
+ bl[124] br[124] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_127 
+ bl[125] br[125] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_128 
+ bl[126] br[126] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_129 
+ bl[127] br[127] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_130 
+ bl[128] br[128] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_131 
+ bl[129] br[129] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_132 
+ bl[130] br[130] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_133 
+ bl[131] br[131] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_134 
+ bl[132] br[132] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_135 
+ bl[133] br[133] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_136 
+ bl[134] br[134] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_137 
+ bl[135] br[135] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_138 
+ bl[136] br[136] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_139 
+ bl[137] br[137] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_140 
+ bl[138] br[138] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_141 
+ bl[139] br[139] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_142 
+ bl[140] br[140] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_143 
+ bl[141] br[141] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_144 
+ bl[142] br[142] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_145 
+ bl[143] br[143] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_146 
+ bl[144] br[144] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_147 
+ bl[145] br[145] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_148 
+ bl[146] br[146] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_149 
+ bl[147] br[147] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_150 
+ bl[148] br[148] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_151 
+ bl[149] br[149] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_152 
+ bl[150] br[150] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_153 
+ bl[151] br[151] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_154 
+ bl[152] br[152] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_155 
+ bl[153] br[153] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_156 
+ bl[154] br[154] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_157 
+ bl[155] br[155] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_158 
+ bl[156] br[156] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_159 
+ bl[157] br[157] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_160 
+ bl[158] br[158] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_161 
+ bl[159] br[159] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_162 
+ bl[160] br[160] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_163 
+ bl[161] br[161] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_164 
+ bl[162] br[162] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_165 
+ bl[163] br[163] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_166 
+ bl[164] br[164] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_167 
+ bl[165] br[165] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_168 
+ bl[166] br[166] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_169 
+ bl[167] br[167] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_170 
+ bl[168] br[168] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_171 
+ bl[169] br[169] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_172 
+ bl[170] br[170] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_173 
+ bl[171] br[171] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_174 
+ bl[172] br[172] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_175 
+ bl[173] br[173] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_176 
+ bl[174] br[174] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_177 
+ bl[175] br[175] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_178 
+ bl[176] br[176] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_179 
+ bl[177] br[177] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_180 
+ bl[178] br[178] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_181 
+ bl[179] br[179] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_182 
+ bl[180] br[180] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_183 
+ bl[181] br[181] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_184 
+ bl[182] br[182] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_185 
+ bl[183] br[183] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_186 
+ bl[184] br[184] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_187 
+ bl[185] br[185] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_188 
+ bl[186] br[186] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_189 
+ bl[187] br[187] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_190 
+ bl[188] br[188] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_191 
+ bl[189] br[189] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_192 
+ bl[190] br[190] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_193 
+ bl[191] br[191] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_194 
+ bl[192] br[192] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_195 
+ bl[193] br[193] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_196 
+ bl[194] br[194] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_197 
+ bl[195] br[195] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_198 
+ bl[196] br[196] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_199 
+ bl[197] br[197] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_200 
+ bl[198] br[198] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_201 
+ bl[199] br[199] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_202 
+ bl[200] br[200] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_203 
+ bl[201] br[201] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_204 
+ bl[202] br[202] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_205 
+ bl[203] br[203] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_206 
+ bl[204] br[204] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_207 
+ bl[205] br[205] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_208 
+ bl[206] br[206] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_209 
+ bl[207] br[207] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_210 
+ bl[208] br[208] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_211 
+ bl[209] br[209] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_212 
+ bl[210] br[210] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_213 
+ bl[211] br[211] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_214 
+ bl[212] br[212] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_215 
+ bl[213] br[213] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_216 
+ bl[214] br[214] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_217 
+ bl[215] br[215] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_218 
+ bl[216] br[216] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_219 
+ bl[217] br[217] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_220 
+ bl[218] br[218] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_221 
+ bl[219] br[219] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_222 
+ bl[220] br[220] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_223 
+ bl[221] br[221] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_224 
+ bl[222] br[222] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_225 
+ bl[223] br[223] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_226 
+ bl[224] br[224] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_227 
+ bl[225] br[225] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_228 
+ bl[226] br[226] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_229 
+ bl[227] br[227] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_230 
+ bl[228] br[228] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_231 
+ bl[229] br[229] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_232 
+ bl[230] br[230] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_233 
+ bl[231] br[231] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_234 
+ bl[232] br[232] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_235 
+ bl[233] br[233] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_236 
+ bl[234] br[234] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_237 
+ bl[235] br[235] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_238 
+ bl[236] br[236] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_239 
+ bl[237] br[237] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_240 
+ bl[238] br[238] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_241 
+ bl[239] br[239] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_242 
+ bl[240] br[240] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_243 
+ bl[241] br[241] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_244 
+ bl[242] br[242] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_245 
+ bl[243] br[243] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_246 
+ bl[244] br[244] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_247 
+ bl[245] br[245] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_248 
+ bl[246] br[246] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_249 
+ bl[247] br[247] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_250 
+ bl[248] br[248] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_251 
+ bl[249] br[249] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_252 
+ bl[250] br[250] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_253 
+ bl[251] br[251] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_254 
+ bl[252] br[252] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_255 
+ bl[253] br[253] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_256 
+ bl[254] br[254] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_257 
+ bl[255] br[255] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_258 
+ vdd vdd vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_259 
+ vdd vdd vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_0 
+ vdd vdd vss vdd vpb vnb wl[17] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_19_1 
+ rbl rbr vss vdd vpb vnb wl[17] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_19_2 
+ bl[0] br[0] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_3 
+ bl[1] br[1] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_4 
+ bl[2] br[2] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_5 
+ bl[3] br[3] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_6 
+ bl[4] br[4] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_7 
+ bl[5] br[5] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_8 
+ bl[6] br[6] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_9 
+ bl[7] br[7] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_10 
+ bl[8] br[8] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_11 
+ bl[9] br[9] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_12 
+ bl[10] br[10] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_13 
+ bl[11] br[11] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_14 
+ bl[12] br[12] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_15 
+ bl[13] br[13] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_16 
+ bl[14] br[14] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_17 
+ bl[15] br[15] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_18 
+ bl[16] br[16] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_19 
+ bl[17] br[17] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_20 
+ bl[18] br[18] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_21 
+ bl[19] br[19] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_22 
+ bl[20] br[20] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_23 
+ bl[21] br[21] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_24 
+ bl[22] br[22] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_25 
+ bl[23] br[23] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_26 
+ bl[24] br[24] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_27 
+ bl[25] br[25] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_28 
+ bl[26] br[26] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_29 
+ bl[27] br[27] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_30 
+ bl[28] br[28] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_31 
+ bl[29] br[29] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_32 
+ bl[30] br[30] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_33 
+ bl[31] br[31] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_34 
+ bl[32] br[32] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_35 
+ bl[33] br[33] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_36 
+ bl[34] br[34] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_37 
+ bl[35] br[35] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_38 
+ bl[36] br[36] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_39 
+ bl[37] br[37] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_40 
+ bl[38] br[38] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_41 
+ bl[39] br[39] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_42 
+ bl[40] br[40] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_43 
+ bl[41] br[41] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_44 
+ bl[42] br[42] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_45 
+ bl[43] br[43] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_46 
+ bl[44] br[44] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_47 
+ bl[45] br[45] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_48 
+ bl[46] br[46] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_49 
+ bl[47] br[47] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_50 
+ bl[48] br[48] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_51 
+ bl[49] br[49] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_52 
+ bl[50] br[50] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_53 
+ bl[51] br[51] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_54 
+ bl[52] br[52] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_55 
+ bl[53] br[53] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_56 
+ bl[54] br[54] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_57 
+ bl[55] br[55] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_58 
+ bl[56] br[56] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_59 
+ bl[57] br[57] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_60 
+ bl[58] br[58] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_61 
+ bl[59] br[59] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_62 
+ bl[60] br[60] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_63 
+ bl[61] br[61] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_64 
+ bl[62] br[62] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_65 
+ bl[63] br[63] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_66 
+ bl[64] br[64] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_67 
+ bl[65] br[65] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_68 
+ bl[66] br[66] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_69 
+ bl[67] br[67] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_70 
+ bl[68] br[68] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_71 
+ bl[69] br[69] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_72 
+ bl[70] br[70] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_73 
+ bl[71] br[71] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_74 
+ bl[72] br[72] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_75 
+ bl[73] br[73] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_76 
+ bl[74] br[74] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_77 
+ bl[75] br[75] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_78 
+ bl[76] br[76] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_79 
+ bl[77] br[77] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_80 
+ bl[78] br[78] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_81 
+ bl[79] br[79] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_82 
+ bl[80] br[80] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_83 
+ bl[81] br[81] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_84 
+ bl[82] br[82] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_85 
+ bl[83] br[83] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_86 
+ bl[84] br[84] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_87 
+ bl[85] br[85] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_88 
+ bl[86] br[86] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_89 
+ bl[87] br[87] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_90 
+ bl[88] br[88] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_91 
+ bl[89] br[89] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_92 
+ bl[90] br[90] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_93 
+ bl[91] br[91] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_94 
+ bl[92] br[92] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_95 
+ bl[93] br[93] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_96 
+ bl[94] br[94] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_97 
+ bl[95] br[95] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_98 
+ bl[96] br[96] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_99 
+ bl[97] br[97] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_100 
+ bl[98] br[98] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_101 
+ bl[99] br[99] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_102 
+ bl[100] br[100] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_103 
+ bl[101] br[101] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_104 
+ bl[102] br[102] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_105 
+ bl[103] br[103] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_106 
+ bl[104] br[104] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_107 
+ bl[105] br[105] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_108 
+ bl[106] br[106] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_109 
+ bl[107] br[107] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_110 
+ bl[108] br[108] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_111 
+ bl[109] br[109] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_112 
+ bl[110] br[110] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_113 
+ bl[111] br[111] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_114 
+ bl[112] br[112] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_115 
+ bl[113] br[113] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_116 
+ bl[114] br[114] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_117 
+ bl[115] br[115] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_118 
+ bl[116] br[116] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_119 
+ bl[117] br[117] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_120 
+ bl[118] br[118] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_121 
+ bl[119] br[119] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_122 
+ bl[120] br[120] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_123 
+ bl[121] br[121] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_124 
+ bl[122] br[122] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_125 
+ bl[123] br[123] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_126 
+ bl[124] br[124] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_127 
+ bl[125] br[125] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_128 
+ bl[126] br[126] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_129 
+ bl[127] br[127] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_130 
+ bl[128] br[128] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_131 
+ bl[129] br[129] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_132 
+ bl[130] br[130] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_133 
+ bl[131] br[131] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_134 
+ bl[132] br[132] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_135 
+ bl[133] br[133] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_136 
+ bl[134] br[134] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_137 
+ bl[135] br[135] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_138 
+ bl[136] br[136] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_139 
+ bl[137] br[137] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_140 
+ bl[138] br[138] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_141 
+ bl[139] br[139] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_142 
+ bl[140] br[140] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_143 
+ bl[141] br[141] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_144 
+ bl[142] br[142] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_145 
+ bl[143] br[143] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_146 
+ bl[144] br[144] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_147 
+ bl[145] br[145] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_148 
+ bl[146] br[146] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_149 
+ bl[147] br[147] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_150 
+ bl[148] br[148] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_151 
+ bl[149] br[149] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_152 
+ bl[150] br[150] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_153 
+ bl[151] br[151] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_154 
+ bl[152] br[152] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_155 
+ bl[153] br[153] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_156 
+ bl[154] br[154] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_157 
+ bl[155] br[155] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_158 
+ bl[156] br[156] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_159 
+ bl[157] br[157] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_160 
+ bl[158] br[158] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_161 
+ bl[159] br[159] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_162 
+ bl[160] br[160] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_163 
+ bl[161] br[161] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_164 
+ bl[162] br[162] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_165 
+ bl[163] br[163] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_166 
+ bl[164] br[164] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_167 
+ bl[165] br[165] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_168 
+ bl[166] br[166] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_169 
+ bl[167] br[167] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_170 
+ bl[168] br[168] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_171 
+ bl[169] br[169] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_172 
+ bl[170] br[170] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_173 
+ bl[171] br[171] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_174 
+ bl[172] br[172] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_175 
+ bl[173] br[173] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_176 
+ bl[174] br[174] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_177 
+ bl[175] br[175] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_178 
+ bl[176] br[176] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_179 
+ bl[177] br[177] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_180 
+ bl[178] br[178] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_181 
+ bl[179] br[179] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_182 
+ bl[180] br[180] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_183 
+ bl[181] br[181] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_184 
+ bl[182] br[182] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_185 
+ bl[183] br[183] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_186 
+ bl[184] br[184] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_187 
+ bl[185] br[185] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_188 
+ bl[186] br[186] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_189 
+ bl[187] br[187] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_190 
+ bl[188] br[188] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_191 
+ bl[189] br[189] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_192 
+ bl[190] br[190] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_193 
+ bl[191] br[191] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_194 
+ bl[192] br[192] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_195 
+ bl[193] br[193] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_196 
+ bl[194] br[194] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_197 
+ bl[195] br[195] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_198 
+ bl[196] br[196] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_199 
+ bl[197] br[197] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_200 
+ bl[198] br[198] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_201 
+ bl[199] br[199] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_202 
+ bl[200] br[200] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_203 
+ bl[201] br[201] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_204 
+ bl[202] br[202] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_205 
+ bl[203] br[203] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_206 
+ bl[204] br[204] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_207 
+ bl[205] br[205] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_208 
+ bl[206] br[206] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_209 
+ bl[207] br[207] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_210 
+ bl[208] br[208] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_211 
+ bl[209] br[209] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_212 
+ bl[210] br[210] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_213 
+ bl[211] br[211] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_214 
+ bl[212] br[212] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_215 
+ bl[213] br[213] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_216 
+ bl[214] br[214] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_217 
+ bl[215] br[215] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_218 
+ bl[216] br[216] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_219 
+ bl[217] br[217] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_220 
+ bl[218] br[218] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_221 
+ bl[219] br[219] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_222 
+ bl[220] br[220] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_223 
+ bl[221] br[221] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_224 
+ bl[222] br[222] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_225 
+ bl[223] br[223] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_226 
+ bl[224] br[224] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_227 
+ bl[225] br[225] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_228 
+ bl[226] br[226] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_229 
+ bl[227] br[227] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_230 
+ bl[228] br[228] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_231 
+ bl[229] br[229] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_232 
+ bl[230] br[230] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_233 
+ bl[231] br[231] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_234 
+ bl[232] br[232] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_235 
+ bl[233] br[233] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_236 
+ bl[234] br[234] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_237 
+ bl[235] br[235] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_238 
+ bl[236] br[236] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_239 
+ bl[237] br[237] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_240 
+ bl[238] br[238] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_241 
+ bl[239] br[239] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_242 
+ bl[240] br[240] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_243 
+ bl[241] br[241] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_244 
+ bl[242] br[242] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_245 
+ bl[243] br[243] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_246 
+ bl[244] br[244] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_247 
+ bl[245] br[245] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_248 
+ bl[246] br[246] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_249 
+ bl[247] br[247] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_250 
+ bl[248] br[248] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_251 
+ bl[249] br[249] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_252 
+ bl[250] br[250] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_253 
+ bl[251] br[251] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_254 
+ bl[252] br[252] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_255 
+ bl[253] br[253] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_256 
+ bl[254] br[254] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_257 
+ bl[255] br[255] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_258 
+ vdd vdd vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_259 
+ vdd vdd vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_0 
+ vdd vdd vss vdd vpb vnb wl[18] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_20_1 
+ rbl rbr vss vdd vpb vnb wl[18] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_20_2 
+ bl[0] br[0] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_3 
+ bl[1] br[1] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_4 
+ bl[2] br[2] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_5 
+ bl[3] br[3] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_6 
+ bl[4] br[4] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_7 
+ bl[5] br[5] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_8 
+ bl[6] br[6] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_9 
+ bl[7] br[7] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_10 
+ bl[8] br[8] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_11 
+ bl[9] br[9] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_12 
+ bl[10] br[10] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_13 
+ bl[11] br[11] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_14 
+ bl[12] br[12] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_15 
+ bl[13] br[13] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_16 
+ bl[14] br[14] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_17 
+ bl[15] br[15] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_18 
+ bl[16] br[16] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_19 
+ bl[17] br[17] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_20 
+ bl[18] br[18] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_21 
+ bl[19] br[19] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_22 
+ bl[20] br[20] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_23 
+ bl[21] br[21] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_24 
+ bl[22] br[22] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_25 
+ bl[23] br[23] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_26 
+ bl[24] br[24] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_27 
+ bl[25] br[25] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_28 
+ bl[26] br[26] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_29 
+ bl[27] br[27] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_30 
+ bl[28] br[28] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_31 
+ bl[29] br[29] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_32 
+ bl[30] br[30] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_33 
+ bl[31] br[31] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_34 
+ bl[32] br[32] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_35 
+ bl[33] br[33] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_36 
+ bl[34] br[34] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_37 
+ bl[35] br[35] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_38 
+ bl[36] br[36] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_39 
+ bl[37] br[37] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_40 
+ bl[38] br[38] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_41 
+ bl[39] br[39] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_42 
+ bl[40] br[40] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_43 
+ bl[41] br[41] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_44 
+ bl[42] br[42] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_45 
+ bl[43] br[43] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_46 
+ bl[44] br[44] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_47 
+ bl[45] br[45] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_48 
+ bl[46] br[46] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_49 
+ bl[47] br[47] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_50 
+ bl[48] br[48] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_51 
+ bl[49] br[49] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_52 
+ bl[50] br[50] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_53 
+ bl[51] br[51] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_54 
+ bl[52] br[52] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_55 
+ bl[53] br[53] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_56 
+ bl[54] br[54] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_57 
+ bl[55] br[55] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_58 
+ bl[56] br[56] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_59 
+ bl[57] br[57] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_60 
+ bl[58] br[58] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_61 
+ bl[59] br[59] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_62 
+ bl[60] br[60] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_63 
+ bl[61] br[61] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_64 
+ bl[62] br[62] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_65 
+ bl[63] br[63] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_66 
+ bl[64] br[64] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_67 
+ bl[65] br[65] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_68 
+ bl[66] br[66] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_69 
+ bl[67] br[67] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_70 
+ bl[68] br[68] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_71 
+ bl[69] br[69] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_72 
+ bl[70] br[70] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_73 
+ bl[71] br[71] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_74 
+ bl[72] br[72] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_75 
+ bl[73] br[73] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_76 
+ bl[74] br[74] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_77 
+ bl[75] br[75] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_78 
+ bl[76] br[76] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_79 
+ bl[77] br[77] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_80 
+ bl[78] br[78] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_81 
+ bl[79] br[79] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_82 
+ bl[80] br[80] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_83 
+ bl[81] br[81] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_84 
+ bl[82] br[82] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_85 
+ bl[83] br[83] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_86 
+ bl[84] br[84] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_87 
+ bl[85] br[85] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_88 
+ bl[86] br[86] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_89 
+ bl[87] br[87] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_90 
+ bl[88] br[88] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_91 
+ bl[89] br[89] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_92 
+ bl[90] br[90] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_93 
+ bl[91] br[91] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_94 
+ bl[92] br[92] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_95 
+ bl[93] br[93] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_96 
+ bl[94] br[94] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_97 
+ bl[95] br[95] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_98 
+ bl[96] br[96] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_99 
+ bl[97] br[97] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_100 
+ bl[98] br[98] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_101 
+ bl[99] br[99] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_102 
+ bl[100] br[100] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_103 
+ bl[101] br[101] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_104 
+ bl[102] br[102] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_105 
+ bl[103] br[103] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_106 
+ bl[104] br[104] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_107 
+ bl[105] br[105] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_108 
+ bl[106] br[106] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_109 
+ bl[107] br[107] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_110 
+ bl[108] br[108] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_111 
+ bl[109] br[109] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_112 
+ bl[110] br[110] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_113 
+ bl[111] br[111] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_114 
+ bl[112] br[112] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_115 
+ bl[113] br[113] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_116 
+ bl[114] br[114] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_117 
+ bl[115] br[115] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_118 
+ bl[116] br[116] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_119 
+ bl[117] br[117] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_120 
+ bl[118] br[118] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_121 
+ bl[119] br[119] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_122 
+ bl[120] br[120] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_123 
+ bl[121] br[121] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_124 
+ bl[122] br[122] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_125 
+ bl[123] br[123] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_126 
+ bl[124] br[124] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_127 
+ bl[125] br[125] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_128 
+ bl[126] br[126] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_129 
+ bl[127] br[127] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_130 
+ bl[128] br[128] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_131 
+ bl[129] br[129] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_132 
+ bl[130] br[130] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_133 
+ bl[131] br[131] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_134 
+ bl[132] br[132] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_135 
+ bl[133] br[133] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_136 
+ bl[134] br[134] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_137 
+ bl[135] br[135] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_138 
+ bl[136] br[136] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_139 
+ bl[137] br[137] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_140 
+ bl[138] br[138] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_141 
+ bl[139] br[139] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_142 
+ bl[140] br[140] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_143 
+ bl[141] br[141] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_144 
+ bl[142] br[142] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_145 
+ bl[143] br[143] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_146 
+ bl[144] br[144] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_147 
+ bl[145] br[145] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_148 
+ bl[146] br[146] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_149 
+ bl[147] br[147] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_150 
+ bl[148] br[148] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_151 
+ bl[149] br[149] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_152 
+ bl[150] br[150] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_153 
+ bl[151] br[151] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_154 
+ bl[152] br[152] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_155 
+ bl[153] br[153] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_156 
+ bl[154] br[154] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_157 
+ bl[155] br[155] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_158 
+ bl[156] br[156] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_159 
+ bl[157] br[157] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_160 
+ bl[158] br[158] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_161 
+ bl[159] br[159] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_162 
+ bl[160] br[160] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_163 
+ bl[161] br[161] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_164 
+ bl[162] br[162] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_165 
+ bl[163] br[163] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_166 
+ bl[164] br[164] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_167 
+ bl[165] br[165] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_168 
+ bl[166] br[166] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_169 
+ bl[167] br[167] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_170 
+ bl[168] br[168] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_171 
+ bl[169] br[169] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_172 
+ bl[170] br[170] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_173 
+ bl[171] br[171] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_174 
+ bl[172] br[172] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_175 
+ bl[173] br[173] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_176 
+ bl[174] br[174] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_177 
+ bl[175] br[175] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_178 
+ bl[176] br[176] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_179 
+ bl[177] br[177] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_180 
+ bl[178] br[178] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_181 
+ bl[179] br[179] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_182 
+ bl[180] br[180] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_183 
+ bl[181] br[181] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_184 
+ bl[182] br[182] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_185 
+ bl[183] br[183] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_186 
+ bl[184] br[184] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_187 
+ bl[185] br[185] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_188 
+ bl[186] br[186] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_189 
+ bl[187] br[187] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_190 
+ bl[188] br[188] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_191 
+ bl[189] br[189] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_192 
+ bl[190] br[190] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_193 
+ bl[191] br[191] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_194 
+ bl[192] br[192] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_195 
+ bl[193] br[193] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_196 
+ bl[194] br[194] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_197 
+ bl[195] br[195] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_198 
+ bl[196] br[196] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_199 
+ bl[197] br[197] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_200 
+ bl[198] br[198] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_201 
+ bl[199] br[199] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_202 
+ bl[200] br[200] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_203 
+ bl[201] br[201] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_204 
+ bl[202] br[202] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_205 
+ bl[203] br[203] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_206 
+ bl[204] br[204] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_207 
+ bl[205] br[205] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_208 
+ bl[206] br[206] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_209 
+ bl[207] br[207] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_210 
+ bl[208] br[208] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_211 
+ bl[209] br[209] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_212 
+ bl[210] br[210] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_213 
+ bl[211] br[211] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_214 
+ bl[212] br[212] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_215 
+ bl[213] br[213] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_216 
+ bl[214] br[214] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_217 
+ bl[215] br[215] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_218 
+ bl[216] br[216] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_219 
+ bl[217] br[217] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_220 
+ bl[218] br[218] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_221 
+ bl[219] br[219] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_222 
+ bl[220] br[220] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_223 
+ bl[221] br[221] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_224 
+ bl[222] br[222] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_225 
+ bl[223] br[223] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_226 
+ bl[224] br[224] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_227 
+ bl[225] br[225] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_228 
+ bl[226] br[226] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_229 
+ bl[227] br[227] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_230 
+ bl[228] br[228] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_231 
+ bl[229] br[229] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_232 
+ bl[230] br[230] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_233 
+ bl[231] br[231] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_234 
+ bl[232] br[232] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_235 
+ bl[233] br[233] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_236 
+ bl[234] br[234] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_237 
+ bl[235] br[235] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_238 
+ bl[236] br[236] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_239 
+ bl[237] br[237] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_240 
+ bl[238] br[238] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_241 
+ bl[239] br[239] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_242 
+ bl[240] br[240] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_243 
+ bl[241] br[241] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_244 
+ bl[242] br[242] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_245 
+ bl[243] br[243] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_246 
+ bl[244] br[244] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_247 
+ bl[245] br[245] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_248 
+ bl[246] br[246] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_249 
+ bl[247] br[247] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_250 
+ bl[248] br[248] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_251 
+ bl[249] br[249] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_252 
+ bl[250] br[250] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_253 
+ bl[251] br[251] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_254 
+ bl[252] br[252] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_255 
+ bl[253] br[253] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_256 
+ bl[254] br[254] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_257 
+ bl[255] br[255] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_258 
+ vdd vdd vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_259 
+ vdd vdd vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_0 
+ vdd vdd vss vdd vpb vnb wl[19] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_21_1 
+ rbl rbr vss vdd vpb vnb wl[19] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_21_2 
+ bl[0] br[0] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_3 
+ bl[1] br[1] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_4 
+ bl[2] br[2] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_5 
+ bl[3] br[3] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_6 
+ bl[4] br[4] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_7 
+ bl[5] br[5] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_8 
+ bl[6] br[6] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_9 
+ bl[7] br[7] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_10 
+ bl[8] br[8] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_11 
+ bl[9] br[9] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_12 
+ bl[10] br[10] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_13 
+ bl[11] br[11] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_14 
+ bl[12] br[12] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_15 
+ bl[13] br[13] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_16 
+ bl[14] br[14] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_17 
+ bl[15] br[15] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_18 
+ bl[16] br[16] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_19 
+ bl[17] br[17] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_20 
+ bl[18] br[18] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_21 
+ bl[19] br[19] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_22 
+ bl[20] br[20] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_23 
+ bl[21] br[21] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_24 
+ bl[22] br[22] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_25 
+ bl[23] br[23] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_26 
+ bl[24] br[24] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_27 
+ bl[25] br[25] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_28 
+ bl[26] br[26] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_29 
+ bl[27] br[27] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_30 
+ bl[28] br[28] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_31 
+ bl[29] br[29] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_32 
+ bl[30] br[30] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_33 
+ bl[31] br[31] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_34 
+ bl[32] br[32] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_35 
+ bl[33] br[33] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_36 
+ bl[34] br[34] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_37 
+ bl[35] br[35] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_38 
+ bl[36] br[36] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_39 
+ bl[37] br[37] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_40 
+ bl[38] br[38] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_41 
+ bl[39] br[39] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_42 
+ bl[40] br[40] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_43 
+ bl[41] br[41] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_44 
+ bl[42] br[42] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_45 
+ bl[43] br[43] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_46 
+ bl[44] br[44] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_47 
+ bl[45] br[45] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_48 
+ bl[46] br[46] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_49 
+ bl[47] br[47] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_50 
+ bl[48] br[48] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_51 
+ bl[49] br[49] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_52 
+ bl[50] br[50] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_53 
+ bl[51] br[51] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_54 
+ bl[52] br[52] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_55 
+ bl[53] br[53] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_56 
+ bl[54] br[54] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_57 
+ bl[55] br[55] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_58 
+ bl[56] br[56] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_59 
+ bl[57] br[57] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_60 
+ bl[58] br[58] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_61 
+ bl[59] br[59] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_62 
+ bl[60] br[60] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_63 
+ bl[61] br[61] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_64 
+ bl[62] br[62] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_65 
+ bl[63] br[63] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_66 
+ bl[64] br[64] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_67 
+ bl[65] br[65] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_68 
+ bl[66] br[66] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_69 
+ bl[67] br[67] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_70 
+ bl[68] br[68] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_71 
+ bl[69] br[69] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_72 
+ bl[70] br[70] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_73 
+ bl[71] br[71] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_74 
+ bl[72] br[72] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_75 
+ bl[73] br[73] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_76 
+ bl[74] br[74] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_77 
+ bl[75] br[75] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_78 
+ bl[76] br[76] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_79 
+ bl[77] br[77] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_80 
+ bl[78] br[78] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_81 
+ bl[79] br[79] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_82 
+ bl[80] br[80] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_83 
+ bl[81] br[81] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_84 
+ bl[82] br[82] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_85 
+ bl[83] br[83] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_86 
+ bl[84] br[84] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_87 
+ bl[85] br[85] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_88 
+ bl[86] br[86] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_89 
+ bl[87] br[87] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_90 
+ bl[88] br[88] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_91 
+ bl[89] br[89] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_92 
+ bl[90] br[90] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_93 
+ bl[91] br[91] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_94 
+ bl[92] br[92] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_95 
+ bl[93] br[93] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_96 
+ bl[94] br[94] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_97 
+ bl[95] br[95] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_98 
+ bl[96] br[96] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_99 
+ bl[97] br[97] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_100 
+ bl[98] br[98] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_101 
+ bl[99] br[99] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_102 
+ bl[100] br[100] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_103 
+ bl[101] br[101] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_104 
+ bl[102] br[102] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_105 
+ bl[103] br[103] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_106 
+ bl[104] br[104] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_107 
+ bl[105] br[105] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_108 
+ bl[106] br[106] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_109 
+ bl[107] br[107] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_110 
+ bl[108] br[108] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_111 
+ bl[109] br[109] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_112 
+ bl[110] br[110] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_113 
+ bl[111] br[111] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_114 
+ bl[112] br[112] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_115 
+ bl[113] br[113] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_116 
+ bl[114] br[114] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_117 
+ bl[115] br[115] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_118 
+ bl[116] br[116] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_119 
+ bl[117] br[117] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_120 
+ bl[118] br[118] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_121 
+ bl[119] br[119] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_122 
+ bl[120] br[120] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_123 
+ bl[121] br[121] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_124 
+ bl[122] br[122] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_125 
+ bl[123] br[123] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_126 
+ bl[124] br[124] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_127 
+ bl[125] br[125] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_128 
+ bl[126] br[126] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_129 
+ bl[127] br[127] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_130 
+ bl[128] br[128] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_131 
+ bl[129] br[129] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_132 
+ bl[130] br[130] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_133 
+ bl[131] br[131] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_134 
+ bl[132] br[132] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_135 
+ bl[133] br[133] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_136 
+ bl[134] br[134] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_137 
+ bl[135] br[135] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_138 
+ bl[136] br[136] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_139 
+ bl[137] br[137] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_140 
+ bl[138] br[138] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_141 
+ bl[139] br[139] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_142 
+ bl[140] br[140] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_143 
+ bl[141] br[141] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_144 
+ bl[142] br[142] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_145 
+ bl[143] br[143] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_146 
+ bl[144] br[144] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_147 
+ bl[145] br[145] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_148 
+ bl[146] br[146] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_149 
+ bl[147] br[147] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_150 
+ bl[148] br[148] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_151 
+ bl[149] br[149] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_152 
+ bl[150] br[150] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_153 
+ bl[151] br[151] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_154 
+ bl[152] br[152] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_155 
+ bl[153] br[153] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_156 
+ bl[154] br[154] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_157 
+ bl[155] br[155] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_158 
+ bl[156] br[156] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_159 
+ bl[157] br[157] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_160 
+ bl[158] br[158] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_161 
+ bl[159] br[159] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_162 
+ bl[160] br[160] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_163 
+ bl[161] br[161] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_164 
+ bl[162] br[162] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_165 
+ bl[163] br[163] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_166 
+ bl[164] br[164] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_167 
+ bl[165] br[165] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_168 
+ bl[166] br[166] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_169 
+ bl[167] br[167] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_170 
+ bl[168] br[168] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_171 
+ bl[169] br[169] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_172 
+ bl[170] br[170] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_173 
+ bl[171] br[171] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_174 
+ bl[172] br[172] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_175 
+ bl[173] br[173] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_176 
+ bl[174] br[174] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_177 
+ bl[175] br[175] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_178 
+ bl[176] br[176] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_179 
+ bl[177] br[177] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_180 
+ bl[178] br[178] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_181 
+ bl[179] br[179] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_182 
+ bl[180] br[180] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_183 
+ bl[181] br[181] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_184 
+ bl[182] br[182] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_185 
+ bl[183] br[183] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_186 
+ bl[184] br[184] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_187 
+ bl[185] br[185] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_188 
+ bl[186] br[186] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_189 
+ bl[187] br[187] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_190 
+ bl[188] br[188] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_191 
+ bl[189] br[189] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_192 
+ bl[190] br[190] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_193 
+ bl[191] br[191] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_194 
+ bl[192] br[192] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_195 
+ bl[193] br[193] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_196 
+ bl[194] br[194] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_197 
+ bl[195] br[195] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_198 
+ bl[196] br[196] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_199 
+ bl[197] br[197] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_200 
+ bl[198] br[198] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_201 
+ bl[199] br[199] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_202 
+ bl[200] br[200] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_203 
+ bl[201] br[201] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_204 
+ bl[202] br[202] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_205 
+ bl[203] br[203] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_206 
+ bl[204] br[204] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_207 
+ bl[205] br[205] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_208 
+ bl[206] br[206] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_209 
+ bl[207] br[207] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_210 
+ bl[208] br[208] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_211 
+ bl[209] br[209] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_212 
+ bl[210] br[210] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_213 
+ bl[211] br[211] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_214 
+ bl[212] br[212] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_215 
+ bl[213] br[213] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_216 
+ bl[214] br[214] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_217 
+ bl[215] br[215] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_218 
+ bl[216] br[216] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_219 
+ bl[217] br[217] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_220 
+ bl[218] br[218] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_221 
+ bl[219] br[219] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_222 
+ bl[220] br[220] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_223 
+ bl[221] br[221] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_224 
+ bl[222] br[222] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_225 
+ bl[223] br[223] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_226 
+ bl[224] br[224] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_227 
+ bl[225] br[225] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_228 
+ bl[226] br[226] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_229 
+ bl[227] br[227] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_230 
+ bl[228] br[228] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_231 
+ bl[229] br[229] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_232 
+ bl[230] br[230] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_233 
+ bl[231] br[231] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_234 
+ bl[232] br[232] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_235 
+ bl[233] br[233] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_236 
+ bl[234] br[234] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_237 
+ bl[235] br[235] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_238 
+ bl[236] br[236] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_239 
+ bl[237] br[237] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_240 
+ bl[238] br[238] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_241 
+ bl[239] br[239] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_242 
+ bl[240] br[240] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_243 
+ bl[241] br[241] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_244 
+ bl[242] br[242] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_245 
+ bl[243] br[243] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_246 
+ bl[244] br[244] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_247 
+ bl[245] br[245] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_248 
+ bl[246] br[246] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_249 
+ bl[247] br[247] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_250 
+ bl[248] br[248] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_251 
+ bl[249] br[249] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_252 
+ bl[250] br[250] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_253 
+ bl[251] br[251] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_254 
+ bl[252] br[252] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_255 
+ bl[253] br[253] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_256 
+ bl[254] br[254] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_257 
+ bl[255] br[255] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_258 
+ vdd vdd vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_259 
+ vdd vdd vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_0 
+ vdd vdd vss vdd vpb vnb wl[20] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_22_1 
+ rbl rbr vss vdd vpb vnb wl[20] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_22_2 
+ bl[0] br[0] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_3 
+ bl[1] br[1] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_4 
+ bl[2] br[2] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_5 
+ bl[3] br[3] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_6 
+ bl[4] br[4] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_7 
+ bl[5] br[5] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_8 
+ bl[6] br[6] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_9 
+ bl[7] br[7] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_10 
+ bl[8] br[8] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_11 
+ bl[9] br[9] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_12 
+ bl[10] br[10] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_13 
+ bl[11] br[11] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_14 
+ bl[12] br[12] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_15 
+ bl[13] br[13] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_16 
+ bl[14] br[14] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_17 
+ bl[15] br[15] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_18 
+ bl[16] br[16] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_19 
+ bl[17] br[17] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_20 
+ bl[18] br[18] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_21 
+ bl[19] br[19] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_22 
+ bl[20] br[20] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_23 
+ bl[21] br[21] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_24 
+ bl[22] br[22] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_25 
+ bl[23] br[23] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_26 
+ bl[24] br[24] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_27 
+ bl[25] br[25] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_28 
+ bl[26] br[26] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_29 
+ bl[27] br[27] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_30 
+ bl[28] br[28] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_31 
+ bl[29] br[29] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_32 
+ bl[30] br[30] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_33 
+ bl[31] br[31] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_34 
+ bl[32] br[32] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_35 
+ bl[33] br[33] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_36 
+ bl[34] br[34] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_37 
+ bl[35] br[35] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_38 
+ bl[36] br[36] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_39 
+ bl[37] br[37] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_40 
+ bl[38] br[38] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_41 
+ bl[39] br[39] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_42 
+ bl[40] br[40] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_43 
+ bl[41] br[41] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_44 
+ bl[42] br[42] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_45 
+ bl[43] br[43] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_46 
+ bl[44] br[44] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_47 
+ bl[45] br[45] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_48 
+ bl[46] br[46] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_49 
+ bl[47] br[47] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_50 
+ bl[48] br[48] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_51 
+ bl[49] br[49] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_52 
+ bl[50] br[50] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_53 
+ bl[51] br[51] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_54 
+ bl[52] br[52] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_55 
+ bl[53] br[53] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_56 
+ bl[54] br[54] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_57 
+ bl[55] br[55] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_58 
+ bl[56] br[56] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_59 
+ bl[57] br[57] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_60 
+ bl[58] br[58] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_61 
+ bl[59] br[59] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_62 
+ bl[60] br[60] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_63 
+ bl[61] br[61] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_64 
+ bl[62] br[62] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_65 
+ bl[63] br[63] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_66 
+ bl[64] br[64] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_67 
+ bl[65] br[65] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_68 
+ bl[66] br[66] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_69 
+ bl[67] br[67] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_70 
+ bl[68] br[68] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_71 
+ bl[69] br[69] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_72 
+ bl[70] br[70] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_73 
+ bl[71] br[71] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_74 
+ bl[72] br[72] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_75 
+ bl[73] br[73] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_76 
+ bl[74] br[74] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_77 
+ bl[75] br[75] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_78 
+ bl[76] br[76] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_79 
+ bl[77] br[77] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_80 
+ bl[78] br[78] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_81 
+ bl[79] br[79] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_82 
+ bl[80] br[80] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_83 
+ bl[81] br[81] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_84 
+ bl[82] br[82] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_85 
+ bl[83] br[83] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_86 
+ bl[84] br[84] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_87 
+ bl[85] br[85] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_88 
+ bl[86] br[86] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_89 
+ bl[87] br[87] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_90 
+ bl[88] br[88] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_91 
+ bl[89] br[89] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_92 
+ bl[90] br[90] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_93 
+ bl[91] br[91] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_94 
+ bl[92] br[92] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_95 
+ bl[93] br[93] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_96 
+ bl[94] br[94] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_97 
+ bl[95] br[95] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_98 
+ bl[96] br[96] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_99 
+ bl[97] br[97] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_100 
+ bl[98] br[98] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_101 
+ bl[99] br[99] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_102 
+ bl[100] br[100] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_103 
+ bl[101] br[101] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_104 
+ bl[102] br[102] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_105 
+ bl[103] br[103] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_106 
+ bl[104] br[104] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_107 
+ bl[105] br[105] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_108 
+ bl[106] br[106] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_109 
+ bl[107] br[107] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_110 
+ bl[108] br[108] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_111 
+ bl[109] br[109] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_112 
+ bl[110] br[110] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_113 
+ bl[111] br[111] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_114 
+ bl[112] br[112] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_115 
+ bl[113] br[113] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_116 
+ bl[114] br[114] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_117 
+ bl[115] br[115] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_118 
+ bl[116] br[116] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_119 
+ bl[117] br[117] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_120 
+ bl[118] br[118] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_121 
+ bl[119] br[119] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_122 
+ bl[120] br[120] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_123 
+ bl[121] br[121] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_124 
+ bl[122] br[122] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_125 
+ bl[123] br[123] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_126 
+ bl[124] br[124] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_127 
+ bl[125] br[125] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_128 
+ bl[126] br[126] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_129 
+ bl[127] br[127] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_130 
+ bl[128] br[128] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_131 
+ bl[129] br[129] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_132 
+ bl[130] br[130] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_133 
+ bl[131] br[131] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_134 
+ bl[132] br[132] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_135 
+ bl[133] br[133] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_136 
+ bl[134] br[134] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_137 
+ bl[135] br[135] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_138 
+ bl[136] br[136] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_139 
+ bl[137] br[137] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_140 
+ bl[138] br[138] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_141 
+ bl[139] br[139] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_142 
+ bl[140] br[140] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_143 
+ bl[141] br[141] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_144 
+ bl[142] br[142] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_145 
+ bl[143] br[143] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_146 
+ bl[144] br[144] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_147 
+ bl[145] br[145] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_148 
+ bl[146] br[146] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_149 
+ bl[147] br[147] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_150 
+ bl[148] br[148] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_151 
+ bl[149] br[149] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_152 
+ bl[150] br[150] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_153 
+ bl[151] br[151] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_154 
+ bl[152] br[152] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_155 
+ bl[153] br[153] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_156 
+ bl[154] br[154] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_157 
+ bl[155] br[155] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_158 
+ bl[156] br[156] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_159 
+ bl[157] br[157] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_160 
+ bl[158] br[158] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_161 
+ bl[159] br[159] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_162 
+ bl[160] br[160] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_163 
+ bl[161] br[161] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_164 
+ bl[162] br[162] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_165 
+ bl[163] br[163] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_166 
+ bl[164] br[164] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_167 
+ bl[165] br[165] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_168 
+ bl[166] br[166] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_169 
+ bl[167] br[167] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_170 
+ bl[168] br[168] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_171 
+ bl[169] br[169] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_172 
+ bl[170] br[170] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_173 
+ bl[171] br[171] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_174 
+ bl[172] br[172] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_175 
+ bl[173] br[173] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_176 
+ bl[174] br[174] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_177 
+ bl[175] br[175] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_178 
+ bl[176] br[176] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_179 
+ bl[177] br[177] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_180 
+ bl[178] br[178] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_181 
+ bl[179] br[179] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_182 
+ bl[180] br[180] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_183 
+ bl[181] br[181] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_184 
+ bl[182] br[182] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_185 
+ bl[183] br[183] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_186 
+ bl[184] br[184] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_187 
+ bl[185] br[185] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_188 
+ bl[186] br[186] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_189 
+ bl[187] br[187] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_190 
+ bl[188] br[188] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_191 
+ bl[189] br[189] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_192 
+ bl[190] br[190] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_193 
+ bl[191] br[191] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_194 
+ bl[192] br[192] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_195 
+ bl[193] br[193] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_196 
+ bl[194] br[194] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_197 
+ bl[195] br[195] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_198 
+ bl[196] br[196] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_199 
+ bl[197] br[197] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_200 
+ bl[198] br[198] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_201 
+ bl[199] br[199] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_202 
+ bl[200] br[200] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_203 
+ bl[201] br[201] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_204 
+ bl[202] br[202] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_205 
+ bl[203] br[203] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_206 
+ bl[204] br[204] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_207 
+ bl[205] br[205] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_208 
+ bl[206] br[206] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_209 
+ bl[207] br[207] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_210 
+ bl[208] br[208] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_211 
+ bl[209] br[209] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_212 
+ bl[210] br[210] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_213 
+ bl[211] br[211] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_214 
+ bl[212] br[212] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_215 
+ bl[213] br[213] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_216 
+ bl[214] br[214] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_217 
+ bl[215] br[215] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_218 
+ bl[216] br[216] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_219 
+ bl[217] br[217] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_220 
+ bl[218] br[218] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_221 
+ bl[219] br[219] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_222 
+ bl[220] br[220] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_223 
+ bl[221] br[221] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_224 
+ bl[222] br[222] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_225 
+ bl[223] br[223] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_226 
+ bl[224] br[224] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_227 
+ bl[225] br[225] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_228 
+ bl[226] br[226] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_229 
+ bl[227] br[227] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_230 
+ bl[228] br[228] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_231 
+ bl[229] br[229] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_232 
+ bl[230] br[230] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_233 
+ bl[231] br[231] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_234 
+ bl[232] br[232] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_235 
+ bl[233] br[233] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_236 
+ bl[234] br[234] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_237 
+ bl[235] br[235] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_238 
+ bl[236] br[236] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_239 
+ bl[237] br[237] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_240 
+ bl[238] br[238] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_241 
+ bl[239] br[239] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_242 
+ bl[240] br[240] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_243 
+ bl[241] br[241] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_244 
+ bl[242] br[242] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_245 
+ bl[243] br[243] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_246 
+ bl[244] br[244] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_247 
+ bl[245] br[245] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_248 
+ bl[246] br[246] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_249 
+ bl[247] br[247] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_250 
+ bl[248] br[248] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_251 
+ bl[249] br[249] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_252 
+ bl[250] br[250] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_253 
+ bl[251] br[251] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_254 
+ bl[252] br[252] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_255 
+ bl[253] br[253] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_256 
+ bl[254] br[254] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_257 
+ bl[255] br[255] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_258 
+ vdd vdd vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_259 
+ vdd vdd vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_0 
+ vdd vdd vss vdd vpb vnb wl[21] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_23_1 
+ rbl rbr vss vdd vpb vnb wl[21] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_23_2 
+ bl[0] br[0] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_3 
+ bl[1] br[1] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_4 
+ bl[2] br[2] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_5 
+ bl[3] br[3] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_6 
+ bl[4] br[4] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_7 
+ bl[5] br[5] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_8 
+ bl[6] br[6] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_9 
+ bl[7] br[7] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_10 
+ bl[8] br[8] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_11 
+ bl[9] br[9] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_12 
+ bl[10] br[10] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_13 
+ bl[11] br[11] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_14 
+ bl[12] br[12] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_15 
+ bl[13] br[13] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_16 
+ bl[14] br[14] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_17 
+ bl[15] br[15] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_18 
+ bl[16] br[16] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_19 
+ bl[17] br[17] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_20 
+ bl[18] br[18] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_21 
+ bl[19] br[19] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_22 
+ bl[20] br[20] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_23 
+ bl[21] br[21] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_24 
+ bl[22] br[22] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_25 
+ bl[23] br[23] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_26 
+ bl[24] br[24] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_27 
+ bl[25] br[25] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_28 
+ bl[26] br[26] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_29 
+ bl[27] br[27] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_30 
+ bl[28] br[28] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_31 
+ bl[29] br[29] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_32 
+ bl[30] br[30] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_33 
+ bl[31] br[31] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_34 
+ bl[32] br[32] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_35 
+ bl[33] br[33] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_36 
+ bl[34] br[34] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_37 
+ bl[35] br[35] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_38 
+ bl[36] br[36] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_39 
+ bl[37] br[37] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_40 
+ bl[38] br[38] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_41 
+ bl[39] br[39] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_42 
+ bl[40] br[40] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_43 
+ bl[41] br[41] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_44 
+ bl[42] br[42] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_45 
+ bl[43] br[43] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_46 
+ bl[44] br[44] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_47 
+ bl[45] br[45] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_48 
+ bl[46] br[46] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_49 
+ bl[47] br[47] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_50 
+ bl[48] br[48] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_51 
+ bl[49] br[49] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_52 
+ bl[50] br[50] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_53 
+ bl[51] br[51] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_54 
+ bl[52] br[52] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_55 
+ bl[53] br[53] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_56 
+ bl[54] br[54] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_57 
+ bl[55] br[55] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_58 
+ bl[56] br[56] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_59 
+ bl[57] br[57] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_60 
+ bl[58] br[58] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_61 
+ bl[59] br[59] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_62 
+ bl[60] br[60] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_63 
+ bl[61] br[61] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_64 
+ bl[62] br[62] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_65 
+ bl[63] br[63] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_66 
+ bl[64] br[64] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_67 
+ bl[65] br[65] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_68 
+ bl[66] br[66] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_69 
+ bl[67] br[67] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_70 
+ bl[68] br[68] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_71 
+ bl[69] br[69] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_72 
+ bl[70] br[70] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_73 
+ bl[71] br[71] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_74 
+ bl[72] br[72] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_75 
+ bl[73] br[73] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_76 
+ bl[74] br[74] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_77 
+ bl[75] br[75] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_78 
+ bl[76] br[76] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_79 
+ bl[77] br[77] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_80 
+ bl[78] br[78] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_81 
+ bl[79] br[79] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_82 
+ bl[80] br[80] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_83 
+ bl[81] br[81] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_84 
+ bl[82] br[82] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_85 
+ bl[83] br[83] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_86 
+ bl[84] br[84] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_87 
+ bl[85] br[85] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_88 
+ bl[86] br[86] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_89 
+ bl[87] br[87] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_90 
+ bl[88] br[88] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_91 
+ bl[89] br[89] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_92 
+ bl[90] br[90] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_93 
+ bl[91] br[91] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_94 
+ bl[92] br[92] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_95 
+ bl[93] br[93] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_96 
+ bl[94] br[94] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_97 
+ bl[95] br[95] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_98 
+ bl[96] br[96] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_99 
+ bl[97] br[97] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_100 
+ bl[98] br[98] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_101 
+ bl[99] br[99] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_102 
+ bl[100] br[100] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_103 
+ bl[101] br[101] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_104 
+ bl[102] br[102] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_105 
+ bl[103] br[103] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_106 
+ bl[104] br[104] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_107 
+ bl[105] br[105] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_108 
+ bl[106] br[106] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_109 
+ bl[107] br[107] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_110 
+ bl[108] br[108] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_111 
+ bl[109] br[109] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_112 
+ bl[110] br[110] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_113 
+ bl[111] br[111] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_114 
+ bl[112] br[112] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_115 
+ bl[113] br[113] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_116 
+ bl[114] br[114] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_117 
+ bl[115] br[115] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_118 
+ bl[116] br[116] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_119 
+ bl[117] br[117] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_120 
+ bl[118] br[118] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_121 
+ bl[119] br[119] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_122 
+ bl[120] br[120] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_123 
+ bl[121] br[121] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_124 
+ bl[122] br[122] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_125 
+ bl[123] br[123] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_126 
+ bl[124] br[124] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_127 
+ bl[125] br[125] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_128 
+ bl[126] br[126] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_129 
+ bl[127] br[127] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_130 
+ bl[128] br[128] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_131 
+ bl[129] br[129] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_132 
+ bl[130] br[130] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_133 
+ bl[131] br[131] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_134 
+ bl[132] br[132] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_135 
+ bl[133] br[133] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_136 
+ bl[134] br[134] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_137 
+ bl[135] br[135] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_138 
+ bl[136] br[136] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_139 
+ bl[137] br[137] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_140 
+ bl[138] br[138] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_141 
+ bl[139] br[139] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_142 
+ bl[140] br[140] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_143 
+ bl[141] br[141] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_144 
+ bl[142] br[142] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_145 
+ bl[143] br[143] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_146 
+ bl[144] br[144] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_147 
+ bl[145] br[145] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_148 
+ bl[146] br[146] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_149 
+ bl[147] br[147] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_150 
+ bl[148] br[148] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_151 
+ bl[149] br[149] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_152 
+ bl[150] br[150] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_153 
+ bl[151] br[151] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_154 
+ bl[152] br[152] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_155 
+ bl[153] br[153] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_156 
+ bl[154] br[154] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_157 
+ bl[155] br[155] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_158 
+ bl[156] br[156] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_159 
+ bl[157] br[157] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_160 
+ bl[158] br[158] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_161 
+ bl[159] br[159] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_162 
+ bl[160] br[160] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_163 
+ bl[161] br[161] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_164 
+ bl[162] br[162] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_165 
+ bl[163] br[163] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_166 
+ bl[164] br[164] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_167 
+ bl[165] br[165] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_168 
+ bl[166] br[166] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_169 
+ bl[167] br[167] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_170 
+ bl[168] br[168] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_171 
+ bl[169] br[169] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_172 
+ bl[170] br[170] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_173 
+ bl[171] br[171] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_174 
+ bl[172] br[172] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_175 
+ bl[173] br[173] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_176 
+ bl[174] br[174] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_177 
+ bl[175] br[175] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_178 
+ bl[176] br[176] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_179 
+ bl[177] br[177] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_180 
+ bl[178] br[178] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_181 
+ bl[179] br[179] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_182 
+ bl[180] br[180] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_183 
+ bl[181] br[181] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_184 
+ bl[182] br[182] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_185 
+ bl[183] br[183] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_186 
+ bl[184] br[184] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_187 
+ bl[185] br[185] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_188 
+ bl[186] br[186] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_189 
+ bl[187] br[187] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_190 
+ bl[188] br[188] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_191 
+ bl[189] br[189] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_192 
+ bl[190] br[190] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_193 
+ bl[191] br[191] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_194 
+ bl[192] br[192] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_195 
+ bl[193] br[193] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_196 
+ bl[194] br[194] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_197 
+ bl[195] br[195] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_198 
+ bl[196] br[196] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_199 
+ bl[197] br[197] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_200 
+ bl[198] br[198] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_201 
+ bl[199] br[199] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_202 
+ bl[200] br[200] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_203 
+ bl[201] br[201] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_204 
+ bl[202] br[202] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_205 
+ bl[203] br[203] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_206 
+ bl[204] br[204] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_207 
+ bl[205] br[205] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_208 
+ bl[206] br[206] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_209 
+ bl[207] br[207] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_210 
+ bl[208] br[208] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_211 
+ bl[209] br[209] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_212 
+ bl[210] br[210] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_213 
+ bl[211] br[211] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_214 
+ bl[212] br[212] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_215 
+ bl[213] br[213] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_216 
+ bl[214] br[214] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_217 
+ bl[215] br[215] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_218 
+ bl[216] br[216] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_219 
+ bl[217] br[217] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_220 
+ bl[218] br[218] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_221 
+ bl[219] br[219] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_222 
+ bl[220] br[220] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_223 
+ bl[221] br[221] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_224 
+ bl[222] br[222] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_225 
+ bl[223] br[223] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_226 
+ bl[224] br[224] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_227 
+ bl[225] br[225] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_228 
+ bl[226] br[226] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_229 
+ bl[227] br[227] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_230 
+ bl[228] br[228] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_231 
+ bl[229] br[229] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_232 
+ bl[230] br[230] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_233 
+ bl[231] br[231] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_234 
+ bl[232] br[232] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_235 
+ bl[233] br[233] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_236 
+ bl[234] br[234] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_237 
+ bl[235] br[235] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_238 
+ bl[236] br[236] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_239 
+ bl[237] br[237] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_240 
+ bl[238] br[238] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_241 
+ bl[239] br[239] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_242 
+ bl[240] br[240] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_243 
+ bl[241] br[241] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_244 
+ bl[242] br[242] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_245 
+ bl[243] br[243] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_246 
+ bl[244] br[244] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_247 
+ bl[245] br[245] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_248 
+ bl[246] br[246] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_249 
+ bl[247] br[247] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_250 
+ bl[248] br[248] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_251 
+ bl[249] br[249] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_252 
+ bl[250] br[250] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_253 
+ bl[251] br[251] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_254 
+ bl[252] br[252] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_255 
+ bl[253] br[253] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_256 
+ bl[254] br[254] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_257 
+ bl[255] br[255] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_258 
+ vdd vdd vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_259 
+ vdd vdd vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_0 
+ vdd vdd vss vdd vpb vnb wl[22] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_24_1 
+ rbl rbr vss vdd vpb vnb wl[22] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_24_2 
+ bl[0] br[0] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_3 
+ bl[1] br[1] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_4 
+ bl[2] br[2] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_5 
+ bl[3] br[3] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_6 
+ bl[4] br[4] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_7 
+ bl[5] br[5] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_8 
+ bl[6] br[6] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_9 
+ bl[7] br[7] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_10 
+ bl[8] br[8] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_11 
+ bl[9] br[9] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_12 
+ bl[10] br[10] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_13 
+ bl[11] br[11] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_14 
+ bl[12] br[12] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_15 
+ bl[13] br[13] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_16 
+ bl[14] br[14] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_17 
+ bl[15] br[15] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_18 
+ bl[16] br[16] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_19 
+ bl[17] br[17] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_20 
+ bl[18] br[18] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_21 
+ bl[19] br[19] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_22 
+ bl[20] br[20] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_23 
+ bl[21] br[21] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_24 
+ bl[22] br[22] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_25 
+ bl[23] br[23] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_26 
+ bl[24] br[24] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_27 
+ bl[25] br[25] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_28 
+ bl[26] br[26] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_29 
+ bl[27] br[27] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_30 
+ bl[28] br[28] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_31 
+ bl[29] br[29] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_32 
+ bl[30] br[30] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_33 
+ bl[31] br[31] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_34 
+ bl[32] br[32] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_35 
+ bl[33] br[33] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_36 
+ bl[34] br[34] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_37 
+ bl[35] br[35] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_38 
+ bl[36] br[36] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_39 
+ bl[37] br[37] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_40 
+ bl[38] br[38] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_41 
+ bl[39] br[39] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_42 
+ bl[40] br[40] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_43 
+ bl[41] br[41] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_44 
+ bl[42] br[42] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_45 
+ bl[43] br[43] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_46 
+ bl[44] br[44] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_47 
+ bl[45] br[45] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_48 
+ bl[46] br[46] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_49 
+ bl[47] br[47] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_50 
+ bl[48] br[48] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_51 
+ bl[49] br[49] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_52 
+ bl[50] br[50] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_53 
+ bl[51] br[51] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_54 
+ bl[52] br[52] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_55 
+ bl[53] br[53] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_56 
+ bl[54] br[54] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_57 
+ bl[55] br[55] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_58 
+ bl[56] br[56] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_59 
+ bl[57] br[57] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_60 
+ bl[58] br[58] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_61 
+ bl[59] br[59] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_62 
+ bl[60] br[60] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_63 
+ bl[61] br[61] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_64 
+ bl[62] br[62] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_65 
+ bl[63] br[63] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_66 
+ bl[64] br[64] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_67 
+ bl[65] br[65] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_68 
+ bl[66] br[66] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_69 
+ bl[67] br[67] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_70 
+ bl[68] br[68] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_71 
+ bl[69] br[69] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_72 
+ bl[70] br[70] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_73 
+ bl[71] br[71] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_74 
+ bl[72] br[72] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_75 
+ bl[73] br[73] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_76 
+ bl[74] br[74] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_77 
+ bl[75] br[75] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_78 
+ bl[76] br[76] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_79 
+ bl[77] br[77] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_80 
+ bl[78] br[78] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_81 
+ bl[79] br[79] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_82 
+ bl[80] br[80] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_83 
+ bl[81] br[81] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_84 
+ bl[82] br[82] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_85 
+ bl[83] br[83] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_86 
+ bl[84] br[84] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_87 
+ bl[85] br[85] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_88 
+ bl[86] br[86] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_89 
+ bl[87] br[87] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_90 
+ bl[88] br[88] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_91 
+ bl[89] br[89] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_92 
+ bl[90] br[90] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_93 
+ bl[91] br[91] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_94 
+ bl[92] br[92] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_95 
+ bl[93] br[93] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_96 
+ bl[94] br[94] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_97 
+ bl[95] br[95] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_98 
+ bl[96] br[96] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_99 
+ bl[97] br[97] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_100 
+ bl[98] br[98] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_101 
+ bl[99] br[99] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_102 
+ bl[100] br[100] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_103 
+ bl[101] br[101] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_104 
+ bl[102] br[102] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_105 
+ bl[103] br[103] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_106 
+ bl[104] br[104] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_107 
+ bl[105] br[105] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_108 
+ bl[106] br[106] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_109 
+ bl[107] br[107] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_110 
+ bl[108] br[108] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_111 
+ bl[109] br[109] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_112 
+ bl[110] br[110] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_113 
+ bl[111] br[111] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_114 
+ bl[112] br[112] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_115 
+ bl[113] br[113] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_116 
+ bl[114] br[114] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_117 
+ bl[115] br[115] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_118 
+ bl[116] br[116] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_119 
+ bl[117] br[117] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_120 
+ bl[118] br[118] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_121 
+ bl[119] br[119] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_122 
+ bl[120] br[120] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_123 
+ bl[121] br[121] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_124 
+ bl[122] br[122] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_125 
+ bl[123] br[123] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_126 
+ bl[124] br[124] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_127 
+ bl[125] br[125] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_128 
+ bl[126] br[126] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_129 
+ bl[127] br[127] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_130 
+ bl[128] br[128] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_131 
+ bl[129] br[129] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_132 
+ bl[130] br[130] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_133 
+ bl[131] br[131] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_134 
+ bl[132] br[132] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_135 
+ bl[133] br[133] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_136 
+ bl[134] br[134] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_137 
+ bl[135] br[135] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_138 
+ bl[136] br[136] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_139 
+ bl[137] br[137] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_140 
+ bl[138] br[138] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_141 
+ bl[139] br[139] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_142 
+ bl[140] br[140] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_143 
+ bl[141] br[141] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_144 
+ bl[142] br[142] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_145 
+ bl[143] br[143] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_146 
+ bl[144] br[144] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_147 
+ bl[145] br[145] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_148 
+ bl[146] br[146] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_149 
+ bl[147] br[147] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_150 
+ bl[148] br[148] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_151 
+ bl[149] br[149] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_152 
+ bl[150] br[150] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_153 
+ bl[151] br[151] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_154 
+ bl[152] br[152] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_155 
+ bl[153] br[153] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_156 
+ bl[154] br[154] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_157 
+ bl[155] br[155] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_158 
+ bl[156] br[156] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_159 
+ bl[157] br[157] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_160 
+ bl[158] br[158] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_161 
+ bl[159] br[159] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_162 
+ bl[160] br[160] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_163 
+ bl[161] br[161] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_164 
+ bl[162] br[162] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_165 
+ bl[163] br[163] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_166 
+ bl[164] br[164] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_167 
+ bl[165] br[165] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_168 
+ bl[166] br[166] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_169 
+ bl[167] br[167] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_170 
+ bl[168] br[168] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_171 
+ bl[169] br[169] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_172 
+ bl[170] br[170] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_173 
+ bl[171] br[171] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_174 
+ bl[172] br[172] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_175 
+ bl[173] br[173] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_176 
+ bl[174] br[174] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_177 
+ bl[175] br[175] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_178 
+ bl[176] br[176] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_179 
+ bl[177] br[177] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_180 
+ bl[178] br[178] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_181 
+ bl[179] br[179] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_182 
+ bl[180] br[180] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_183 
+ bl[181] br[181] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_184 
+ bl[182] br[182] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_185 
+ bl[183] br[183] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_186 
+ bl[184] br[184] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_187 
+ bl[185] br[185] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_188 
+ bl[186] br[186] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_189 
+ bl[187] br[187] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_190 
+ bl[188] br[188] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_191 
+ bl[189] br[189] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_192 
+ bl[190] br[190] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_193 
+ bl[191] br[191] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_194 
+ bl[192] br[192] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_195 
+ bl[193] br[193] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_196 
+ bl[194] br[194] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_197 
+ bl[195] br[195] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_198 
+ bl[196] br[196] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_199 
+ bl[197] br[197] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_200 
+ bl[198] br[198] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_201 
+ bl[199] br[199] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_202 
+ bl[200] br[200] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_203 
+ bl[201] br[201] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_204 
+ bl[202] br[202] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_205 
+ bl[203] br[203] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_206 
+ bl[204] br[204] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_207 
+ bl[205] br[205] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_208 
+ bl[206] br[206] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_209 
+ bl[207] br[207] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_210 
+ bl[208] br[208] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_211 
+ bl[209] br[209] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_212 
+ bl[210] br[210] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_213 
+ bl[211] br[211] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_214 
+ bl[212] br[212] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_215 
+ bl[213] br[213] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_216 
+ bl[214] br[214] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_217 
+ bl[215] br[215] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_218 
+ bl[216] br[216] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_219 
+ bl[217] br[217] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_220 
+ bl[218] br[218] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_221 
+ bl[219] br[219] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_222 
+ bl[220] br[220] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_223 
+ bl[221] br[221] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_224 
+ bl[222] br[222] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_225 
+ bl[223] br[223] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_226 
+ bl[224] br[224] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_227 
+ bl[225] br[225] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_228 
+ bl[226] br[226] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_229 
+ bl[227] br[227] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_230 
+ bl[228] br[228] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_231 
+ bl[229] br[229] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_232 
+ bl[230] br[230] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_233 
+ bl[231] br[231] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_234 
+ bl[232] br[232] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_235 
+ bl[233] br[233] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_236 
+ bl[234] br[234] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_237 
+ bl[235] br[235] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_238 
+ bl[236] br[236] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_239 
+ bl[237] br[237] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_240 
+ bl[238] br[238] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_241 
+ bl[239] br[239] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_242 
+ bl[240] br[240] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_243 
+ bl[241] br[241] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_244 
+ bl[242] br[242] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_245 
+ bl[243] br[243] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_246 
+ bl[244] br[244] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_247 
+ bl[245] br[245] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_248 
+ bl[246] br[246] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_249 
+ bl[247] br[247] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_250 
+ bl[248] br[248] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_251 
+ bl[249] br[249] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_252 
+ bl[250] br[250] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_253 
+ bl[251] br[251] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_254 
+ bl[252] br[252] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_255 
+ bl[253] br[253] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_256 
+ bl[254] br[254] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_257 
+ bl[255] br[255] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_258 
+ vdd vdd vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_259 
+ vdd vdd vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_0 
+ vdd vdd vss vdd vpb vnb wl[23] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_25_1 
+ rbl rbr vss vdd vpb vnb wl[23] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_25_2 
+ bl[0] br[0] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_3 
+ bl[1] br[1] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_4 
+ bl[2] br[2] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_5 
+ bl[3] br[3] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_6 
+ bl[4] br[4] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_7 
+ bl[5] br[5] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_8 
+ bl[6] br[6] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_9 
+ bl[7] br[7] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_10 
+ bl[8] br[8] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_11 
+ bl[9] br[9] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_12 
+ bl[10] br[10] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_13 
+ bl[11] br[11] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_14 
+ bl[12] br[12] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_15 
+ bl[13] br[13] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_16 
+ bl[14] br[14] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_17 
+ bl[15] br[15] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_18 
+ bl[16] br[16] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_19 
+ bl[17] br[17] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_20 
+ bl[18] br[18] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_21 
+ bl[19] br[19] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_22 
+ bl[20] br[20] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_23 
+ bl[21] br[21] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_24 
+ bl[22] br[22] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_25 
+ bl[23] br[23] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_26 
+ bl[24] br[24] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_27 
+ bl[25] br[25] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_28 
+ bl[26] br[26] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_29 
+ bl[27] br[27] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_30 
+ bl[28] br[28] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_31 
+ bl[29] br[29] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_32 
+ bl[30] br[30] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_33 
+ bl[31] br[31] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_34 
+ bl[32] br[32] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_35 
+ bl[33] br[33] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_36 
+ bl[34] br[34] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_37 
+ bl[35] br[35] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_38 
+ bl[36] br[36] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_39 
+ bl[37] br[37] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_40 
+ bl[38] br[38] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_41 
+ bl[39] br[39] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_42 
+ bl[40] br[40] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_43 
+ bl[41] br[41] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_44 
+ bl[42] br[42] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_45 
+ bl[43] br[43] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_46 
+ bl[44] br[44] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_47 
+ bl[45] br[45] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_48 
+ bl[46] br[46] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_49 
+ bl[47] br[47] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_50 
+ bl[48] br[48] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_51 
+ bl[49] br[49] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_52 
+ bl[50] br[50] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_53 
+ bl[51] br[51] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_54 
+ bl[52] br[52] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_55 
+ bl[53] br[53] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_56 
+ bl[54] br[54] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_57 
+ bl[55] br[55] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_58 
+ bl[56] br[56] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_59 
+ bl[57] br[57] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_60 
+ bl[58] br[58] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_61 
+ bl[59] br[59] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_62 
+ bl[60] br[60] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_63 
+ bl[61] br[61] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_64 
+ bl[62] br[62] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_65 
+ bl[63] br[63] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_66 
+ bl[64] br[64] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_67 
+ bl[65] br[65] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_68 
+ bl[66] br[66] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_69 
+ bl[67] br[67] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_70 
+ bl[68] br[68] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_71 
+ bl[69] br[69] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_72 
+ bl[70] br[70] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_73 
+ bl[71] br[71] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_74 
+ bl[72] br[72] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_75 
+ bl[73] br[73] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_76 
+ bl[74] br[74] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_77 
+ bl[75] br[75] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_78 
+ bl[76] br[76] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_79 
+ bl[77] br[77] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_80 
+ bl[78] br[78] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_81 
+ bl[79] br[79] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_82 
+ bl[80] br[80] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_83 
+ bl[81] br[81] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_84 
+ bl[82] br[82] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_85 
+ bl[83] br[83] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_86 
+ bl[84] br[84] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_87 
+ bl[85] br[85] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_88 
+ bl[86] br[86] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_89 
+ bl[87] br[87] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_90 
+ bl[88] br[88] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_91 
+ bl[89] br[89] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_92 
+ bl[90] br[90] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_93 
+ bl[91] br[91] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_94 
+ bl[92] br[92] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_95 
+ bl[93] br[93] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_96 
+ bl[94] br[94] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_97 
+ bl[95] br[95] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_98 
+ bl[96] br[96] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_99 
+ bl[97] br[97] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_100 
+ bl[98] br[98] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_101 
+ bl[99] br[99] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_102 
+ bl[100] br[100] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_103 
+ bl[101] br[101] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_104 
+ bl[102] br[102] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_105 
+ bl[103] br[103] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_106 
+ bl[104] br[104] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_107 
+ bl[105] br[105] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_108 
+ bl[106] br[106] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_109 
+ bl[107] br[107] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_110 
+ bl[108] br[108] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_111 
+ bl[109] br[109] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_112 
+ bl[110] br[110] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_113 
+ bl[111] br[111] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_114 
+ bl[112] br[112] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_115 
+ bl[113] br[113] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_116 
+ bl[114] br[114] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_117 
+ bl[115] br[115] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_118 
+ bl[116] br[116] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_119 
+ bl[117] br[117] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_120 
+ bl[118] br[118] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_121 
+ bl[119] br[119] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_122 
+ bl[120] br[120] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_123 
+ bl[121] br[121] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_124 
+ bl[122] br[122] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_125 
+ bl[123] br[123] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_126 
+ bl[124] br[124] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_127 
+ bl[125] br[125] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_128 
+ bl[126] br[126] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_129 
+ bl[127] br[127] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_130 
+ bl[128] br[128] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_131 
+ bl[129] br[129] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_132 
+ bl[130] br[130] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_133 
+ bl[131] br[131] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_134 
+ bl[132] br[132] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_135 
+ bl[133] br[133] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_136 
+ bl[134] br[134] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_137 
+ bl[135] br[135] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_138 
+ bl[136] br[136] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_139 
+ bl[137] br[137] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_140 
+ bl[138] br[138] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_141 
+ bl[139] br[139] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_142 
+ bl[140] br[140] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_143 
+ bl[141] br[141] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_144 
+ bl[142] br[142] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_145 
+ bl[143] br[143] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_146 
+ bl[144] br[144] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_147 
+ bl[145] br[145] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_148 
+ bl[146] br[146] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_149 
+ bl[147] br[147] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_150 
+ bl[148] br[148] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_151 
+ bl[149] br[149] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_152 
+ bl[150] br[150] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_153 
+ bl[151] br[151] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_154 
+ bl[152] br[152] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_155 
+ bl[153] br[153] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_156 
+ bl[154] br[154] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_157 
+ bl[155] br[155] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_158 
+ bl[156] br[156] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_159 
+ bl[157] br[157] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_160 
+ bl[158] br[158] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_161 
+ bl[159] br[159] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_162 
+ bl[160] br[160] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_163 
+ bl[161] br[161] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_164 
+ bl[162] br[162] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_165 
+ bl[163] br[163] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_166 
+ bl[164] br[164] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_167 
+ bl[165] br[165] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_168 
+ bl[166] br[166] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_169 
+ bl[167] br[167] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_170 
+ bl[168] br[168] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_171 
+ bl[169] br[169] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_172 
+ bl[170] br[170] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_173 
+ bl[171] br[171] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_174 
+ bl[172] br[172] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_175 
+ bl[173] br[173] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_176 
+ bl[174] br[174] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_177 
+ bl[175] br[175] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_178 
+ bl[176] br[176] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_179 
+ bl[177] br[177] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_180 
+ bl[178] br[178] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_181 
+ bl[179] br[179] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_182 
+ bl[180] br[180] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_183 
+ bl[181] br[181] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_184 
+ bl[182] br[182] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_185 
+ bl[183] br[183] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_186 
+ bl[184] br[184] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_187 
+ bl[185] br[185] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_188 
+ bl[186] br[186] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_189 
+ bl[187] br[187] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_190 
+ bl[188] br[188] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_191 
+ bl[189] br[189] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_192 
+ bl[190] br[190] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_193 
+ bl[191] br[191] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_194 
+ bl[192] br[192] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_195 
+ bl[193] br[193] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_196 
+ bl[194] br[194] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_197 
+ bl[195] br[195] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_198 
+ bl[196] br[196] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_199 
+ bl[197] br[197] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_200 
+ bl[198] br[198] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_201 
+ bl[199] br[199] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_202 
+ bl[200] br[200] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_203 
+ bl[201] br[201] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_204 
+ bl[202] br[202] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_205 
+ bl[203] br[203] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_206 
+ bl[204] br[204] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_207 
+ bl[205] br[205] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_208 
+ bl[206] br[206] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_209 
+ bl[207] br[207] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_210 
+ bl[208] br[208] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_211 
+ bl[209] br[209] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_212 
+ bl[210] br[210] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_213 
+ bl[211] br[211] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_214 
+ bl[212] br[212] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_215 
+ bl[213] br[213] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_216 
+ bl[214] br[214] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_217 
+ bl[215] br[215] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_218 
+ bl[216] br[216] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_219 
+ bl[217] br[217] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_220 
+ bl[218] br[218] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_221 
+ bl[219] br[219] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_222 
+ bl[220] br[220] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_223 
+ bl[221] br[221] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_224 
+ bl[222] br[222] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_225 
+ bl[223] br[223] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_226 
+ bl[224] br[224] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_227 
+ bl[225] br[225] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_228 
+ bl[226] br[226] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_229 
+ bl[227] br[227] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_230 
+ bl[228] br[228] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_231 
+ bl[229] br[229] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_232 
+ bl[230] br[230] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_233 
+ bl[231] br[231] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_234 
+ bl[232] br[232] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_235 
+ bl[233] br[233] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_236 
+ bl[234] br[234] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_237 
+ bl[235] br[235] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_238 
+ bl[236] br[236] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_239 
+ bl[237] br[237] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_240 
+ bl[238] br[238] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_241 
+ bl[239] br[239] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_242 
+ bl[240] br[240] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_243 
+ bl[241] br[241] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_244 
+ bl[242] br[242] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_245 
+ bl[243] br[243] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_246 
+ bl[244] br[244] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_247 
+ bl[245] br[245] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_248 
+ bl[246] br[246] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_249 
+ bl[247] br[247] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_250 
+ bl[248] br[248] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_251 
+ bl[249] br[249] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_252 
+ bl[250] br[250] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_253 
+ bl[251] br[251] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_254 
+ bl[252] br[252] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_255 
+ bl[253] br[253] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_256 
+ bl[254] br[254] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_257 
+ bl[255] br[255] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_258 
+ vdd vdd vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_259 
+ vdd vdd vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_0 
+ vdd vdd vss vdd vpb vnb wl[24] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_26_1 
+ rbl rbr vss vdd vpb vnb wl[24] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_26_2 
+ bl[0] br[0] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_3 
+ bl[1] br[1] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_4 
+ bl[2] br[2] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_5 
+ bl[3] br[3] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_6 
+ bl[4] br[4] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_7 
+ bl[5] br[5] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_8 
+ bl[6] br[6] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_9 
+ bl[7] br[7] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_10 
+ bl[8] br[8] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_11 
+ bl[9] br[9] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_12 
+ bl[10] br[10] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_13 
+ bl[11] br[11] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_14 
+ bl[12] br[12] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_15 
+ bl[13] br[13] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_16 
+ bl[14] br[14] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_17 
+ bl[15] br[15] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_18 
+ bl[16] br[16] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_19 
+ bl[17] br[17] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_20 
+ bl[18] br[18] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_21 
+ bl[19] br[19] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_22 
+ bl[20] br[20] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_23 
+ bl[21] br[21] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_24 
+ bl[22] br[22] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_25 
+ bl[23] br[23] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_26 
+ bl[24] br[24] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_27 
+ bl[25] br[25] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_28 
+ bl[26] br[26] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_29 
+ bl[27] br[27] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_30 
+ bl[28] br[28] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_31 
+ bl[29] br[29] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_32 
+ bl[30] br[30] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_33 
+ bl[31] br[31] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_34 
+ bl[32] br[32] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_35 
+ bl[33] br[33] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_36 
+ bl[34] br[34] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_37 
+ bl[35] br[35] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_38 
+ bl[36] br[36] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_39 
+ bl[37] br[37] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_40 
+ bl[38] br[38] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_41 
+ bl[39] br[39] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_42 
+ bl[40] br[40] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_43 
+ bl[41] br[41] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_44 
+ bl[42] br[42] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_45 
+ bl[43] br[43] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_46 
+ bl[44] br[44] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_47 
+ bl[45] br[45] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_48 
+ bl[46] br[46] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_49 
+ bl[47] br[47] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_50 
+ bl[48] br[48] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_51 
+ bl[49] br[49] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_52 
+ bl[50] br[50] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_53 
+ bl[51] br[51] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_54 
+ bl[52] br[52] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_55 
+ bl[53] br[53] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_56 
+ bl[54] br[54] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_57 
+ bl[55] br[55] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_58 
+ bl[56] br[56] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_59 
+ bl[57] br[57] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_60 
+ bl[58] br[58] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_61 
+ bl[59] br[59] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_62 
+ bl[60] br[60] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_63 
+ bl[61] br[61] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_64 
+ bl[62] br[62] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_65 
+ bl[63] br[63] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_66 
+ bl[64] br[64] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_67 
+ bl[65] br[65] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_68 
+ bl[66] br[66] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_69 
+ bl[67] br[67] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_70 
+ bl[68] br[68] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_71 
+ bl[69] br[69] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_72 
+ bl[70] br[70] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_73 
+ bl[71] br[71] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_74 
+ bl[72] br[72] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_75 
+ bl[73] br[73] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_76 
+ bl[74] br[74] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_77 
+ bl[75] br[75] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_78 
+ bl[76] br[76] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_79 
+ bl[77] br[77] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_80 
+ bl[78] br[78] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_81 
+ bl[79] br[79] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_82 
+ bl[80] br[80] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_83 
+ bl[81] br[81] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_84 
+ bl[82] br[82] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_85 
+ bl[83] br[83] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_86 
+ bl[84] br[84] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_87 
+ bl[85] br[85] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_88 
+ bl[86] br[86] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_89 
+ bl[87] br[87] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_90 
+ bl[88] br[88] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_91 
+ bl[89] br[89] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_92 
+ bl[90] br[90] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_93 
+ bl[91] br[91] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_94 
+ bl[92] br[92] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_95 
+ bl[93] br[93] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_96 
+ bl[94] br[94] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_97 
+ bl[95] br[95] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_98 
+ bl[96] br[96] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_99 
+ bl[97] br[97] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_100 
+ bl[98] br[98] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_101 
+ bl[99] br[99] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_102 
+ bl[100] br[100] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_103 
+ bl[101] br[101] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_104 
+ bl[102] br[102] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_105 
+ bl[103] br[103] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_106 
+ bl[104] br[104] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_107 
+ bl[105] br[105] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_108 
+ bl[106] br[106] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_109 
+ bl[107] br[107] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_110 
+ bl[108] br[108] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_111 
+ bl[109] br[109] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_112 
+ bl[110] br[110] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_113 
+ bl[111] br[111] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_114 
+ bl[112] br[112] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_115 
+ bl[113] br[113] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_116 
+ bl[114] br[114] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_117 
+ bl[115] br[115] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_118 
+ bl[116] br[116] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_119 
+ bl[117] br[117] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_120 
+ bl[118] br[118] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_121 
+ bl[119] br[119] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_122 
+ bl[120] br[120] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_123 
+ bl[121] br[121] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_124 
+ bl[122] br[122] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_125 
+ bl[123] br[123] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_126 
+ bl[124] br[124] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_127 
+ bl[125] br[125] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_128 
+ bl[126] br[126] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_129 
+ bl[127] br[127] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_130 
+ bl[128] br[128] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_131 
+ bl[129] br[129] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_132 
+ bl[130] br[130] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_133 
+ bl[131] br[131] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_134 
+ bl[132] br[132] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_135 
+ bl[133] br[133] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_136 
+ bl[134] br[134] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_137 
+ bl[135] br[135] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_138 
+ bl[136] br[136] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_139 
+ bl[137] br[137] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_140 
+ bl[138] br[138] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_141 
+ bl[139] br[139] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_142 
+ bl[140] br[140] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_143 
+ bl[141] br[141] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_144 
+ bl[142] br[142] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_145 
+ bl[143] br[143] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_146 
+ bl[144] br[144] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_147 
+ bl[145] br[145] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_148 
+ bl[146] br[146] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_149 
+ bl[147] br[147] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_150 
+ bl[148] br[148] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_151 
+ bl[149] br[149] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_152 
+ bl[150] br[150] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_153 
+ bl[151] br[151] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_154 
+ bl[152] br[152] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_155 
+ bl[153] br[153] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_156 
+ bl[154] br[154] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_157 
+ bl[155] br[155] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_158 
+ bl[156] br[156] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_159 
+ bl[157] br[157] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_160 
+ bl[158] br[158] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_161 
+ bl[159] br[159] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_162 
+ bl[160] br[160] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_163 
+ bl[161] br[161] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_164 
+ bl[162] br[162] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_165 
+ bl[163] br[163] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_166 
+ bl[164] br[164] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_167 
+ bl[165] br[165] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_168 
+ bl[166] br[166] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_169 
+ bl[167] br[167] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_170 
+ bl[168] br[168] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_171 
+ bl[169] br[169] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_172 
+ bl[170] br[170] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_173 
+ bl[171] br[171] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_174 
+ bl[172] br[172] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_175 
+ bl[173] br[173] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_176 
+ bl[174] br[174] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_177 
+ bl[175] br[175] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_178 
+ bl[176] br[176] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_179 
+ bl[177] br[177] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_180 
+ bl[178] br[178] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_181 
+ bl[179] br[179] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_182 
+ bl[180] br[180] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_183 
+ bl[181] br[181] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_184 
+ bl[182] br[182] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_185 
+ bl[183] br[183] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_186 
+ bl[184] br[184] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_187 
+ bl[185] br[185] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_188 
+ bl[186] br[186] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_189 
+ bl[187] br[187] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_190 
+ bl[188] br[188] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_191 
+ bl[189] br[189] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_192 
+ bl[190] br[190] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_193 
+ bl[191] br[191] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_194 
+ bl[192] br[192] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_195 
+ bl[193] br[193] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_196 
+ bl[194] br[194] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_197 
+ bl[195] br[195] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_198 
+ bl[196] br[196] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_199 
+ bl[197] br[197] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_200 
+ bl[198] br[198] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_201 
+ bl[199] br[199] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_202 
+ bl[200] br[200] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_203 
+ bl[201] br[201] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_204 
+ bl[202] br[202] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_205 
+ bl[203] br[203] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_206 
+ bl[204] br[204] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_207 
+ bl[205] br[205] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_208 
+ bl[206] br[206] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_209 
+ bl[207] br[207] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_210 
+ bl[208] br[208] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_211 
+ bl[209] br[209] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_212 
+ bl[210] br[210] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_213 
+ bl[211] br[211] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_214 
+ bl[212] br[212] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_215 
+ bl[213] br[213] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_216 
+ bl[214] br[214] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_217 
+ bl[215] br[215] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_218 
+ bl[216] br[216] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_219 
+ bl[217] br[217] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_220 
+ bl[218] br[218] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_221 
+ bl[219] br[219] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_222 
+ bl[220] br[220] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_223 
+ bl[221] br[221] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_224 
+ bl[222] br[222] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_225 
+ bl[223] br[223] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_226 
+ bl[224] br[224] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_227 
+ bl[225] br[225] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_228 
+ bl[226] br[226] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_229 
+ bl[227] br[227] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_230 
+ bl[228] br[228] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_231 
+ bl[229] br[229] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_232 
+ bl[230] br[230] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_233 
+ bl[231] br[231] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_234 
+ bl[232] br[232] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_235 
+ bl[233] br[233] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_236 
+ bl[234] br[234] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_237 
+ bl[235] br[235] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_238 
+ bl[236] br[236] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_239 
+ bl[237] br[237] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_240 
+ bl[238] br[238] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_241 
+ bl[239] br[239] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_242 
+ bl[240] br[240] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_243 
+ bl[241] br[241] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_244 
+ bl[242] br[242] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_245 
+ bl[243] br[243] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_246 
+ bl[244] br[244] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_247 
+ bl[245] br[245] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_248 
+ bl[246] br[246] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_249 
+ bl[247] br[247] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_250 
+ bl[248] br[248] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_251 
+ bl[249] br[249] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_252 
+ bl[250] br[250] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_253 
+ bl[251] br[251] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_254 
+ bl[252] br[252] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_255 
+ bl[253] br[253] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_256 
+ bl[254] br[254] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_257 
+ bl[255] br[255] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_258 
+ vdd vdd vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_259 
+ vdd vdd vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_0 
+ vdd vdd vss vdd vpb vnb wl[25] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_27_1 
+ rbl rbr vss vdd vpb vnb wl[25] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_27_2 
+ bl[0] br[0] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_3 
+ bl[1] br[1] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_4 
+ bl[2] br[2] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_5 
+ bl[3] br[3] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_6 
+ bl[4] br[4] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_7 
+ bl[5] br[5] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_8 
+ bl[6] br[6] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_9 
+ bl[7] br[7] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_10 
+ bl[8] br[8] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_11 
+ bl[9] br[9] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_12 
+ bl[10] br[10] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_13 
+ bl[11] br[11] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_14 
+ bl[12] br[12] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_15 
+ bl[13] br[13] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_16 
+ bl[14] br[14] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_17 
+ bl[15] br[15] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_18 
+ bl[16] br[16] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_19 
+ bl[17] br[17] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_20 
+ bl[18] br[18] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_21 
+ bl[19] br[19] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_22 
+ bl[20] br[20] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_23 
+ bl[21] br[21] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_24 
+ bl[22] br[22] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_25 
+ bl[23] br[23] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_26 
+ bl[24] br[24] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_27 
+ bl[25] br[25] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_28 
+ bl[26] br[26] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_29 
+ bl[27] br[27] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_30 
+ bl[28] br[28] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_31 
+ bl[29] br[29] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_32 
+ bl[30] br[30] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_33 
+ bl[31] br[31] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_34 
+ bl[32] br[32] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_35 
+ bl[33] br[33] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_36 
+ bl[34] br[34] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_37 
+ bl[35] br[35] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_38 
+ bl[36] br[36] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_39 
+ bl[37] br[37] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_40 
+ bl[38] br[38] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_41 
+ bl[39] br[39] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_42 
+ bl[40] br[40] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_43 
+ bl[41] br[41] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_44 
+ bl[42] br[42] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_45 
+ bl[43] br[43] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_46 
+ bl[44] br[44] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_47 
+ bl[45] br[45] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_48 
+ bl[46] br[46] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_49 
+ bl[47] br[47] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_50 
+ bl[48] br[48] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_51 
+ bl[49] br[49] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_52 
+ bl[50] br[50] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_53 
+ bl[51] br[51] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_54 
+ bl[52] br[52] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_55 
+ bl[53] br[53] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_56 
+ bl[54] br[54] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_57 
+ bl[55] br[55] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_58 
+ bl[56] br[56] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_59 
+ bl[57] br[57] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_60 
+ bl[58] br[58] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_61 
+ bl[59] br[59] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_62 
+ bl[60] br[60] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_63 
+ bl[61] br[61] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_64 
+ bl[62] br[62] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_65 
+ bl[63] br[63] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_66 
+ bl[64] br[64] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_67 
+ bl[65] br[65] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_68 
+ bl[66] br[66] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_69 
+ bl[67] br[67] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_70 
+ bl[68] br[68] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_71 
+ bl[69] br[69] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_72 
+ bl[70] br[70] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_73 
+ bl[71] br[71] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_74 
+ bl[72] br[72] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_75 
+ bl[73] br[73] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_76 
+ bl[74] br[74] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_77 
+ bl[75] br[75] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_78 
+ bl[76] br[76] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_79 
+ bl[77] br[77] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_80 
+ bl[78] br[78] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_81 
+ bl[79] br[79] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_82 
+ bl[80] br[80] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_83 
+ bl[81] br[81] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_84 
+ bl[82] br[82] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_85 
+ bl[83] br[83] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_86 
+ bl[84] br[84] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_87 
+ bl[85] br[85] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_88 
+ bl[86] br[86] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_89 
+ bl[87] br[87] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_90 
+ bl[88] br[88] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_91 
+ bl[89] br[89] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_92 
+ bl[90] br[90] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_93 
+ bl[91] br[91] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_94 
+ bl[92] br[92] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_95 
+ bl[93] br[93] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_96 
+ bl[94] br[94] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_97 
+ bl[95] br[95] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_98 
+ bl[96] br[96] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_99 
+ bl[97] br[97] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_100 
+ bl[98] br[98] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_101 
+ bl[99] br[99] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_102 
+ bl[100] br[100] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_103 
+ bl[101] br[101] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_104 
+ bl[102] br[102] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_105 
+ bl[103] br[103] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_106 
+ bl[104] br[104] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_107 
+ bl[105] br[105] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_108 
+ bl[106] br[106] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_109 
+ bl[107] br[107] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_110 
+ bl[108] br[108] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_111 
+ bl[109] br[109] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_112 
+ bl[110] br[110] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_113 
+ bl[111] br[111] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_114 
+ bl[112] br[112] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_115 
+ bl[113] br[113] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_116 
+ bl[114] br[114] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_117 
+ bl[115] br[115] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_118 
+ bl[116] br[116] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_119 
+ bl[117] br[117] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_120 
+ bl[118] br[118] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_121 
+ bl[119] br[119] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_122 
+ bl[120] br[120] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_123 
+ bl[121] br[121] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_124 
+ bl[122] br[122] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_125 
+ bl[123] br[123] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_126 
+ bl[124] br[124] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_127 
+ bl[125] br[125] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_128 
+ bl[126] br[126] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_129 
+ bl[127] br[127] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_130 
+ bl[128] br[128] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_131 
+ bl[129] br[129] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_132 
+ bl[130] br[130] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_133 
+ bl[131] br[131] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_134 
+ bl[132] br[132] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_135 
+ bl[133] br[133] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_136 
+ bl[134] br[134] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_137 
+ bl[135] br[135] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_138 
+ bl[136] br[136] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_139 
+ bl[137] br[137] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_140 
+ bl[138] br[138] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_141 
+ bl[139] br[139] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_142 
+ bl[140] br[140] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_143 
+ bl[141] br[141] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_144 
+ bl[142] br[142] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_145 
+ bl[143] br[143] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_146 
+ bl[144] br[144] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_147 
+ bl[145] br[145] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_148 
+ bl[146] br[146] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_149 
+ bl[147] br[147] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_150 
+ bl[148] br[148] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_151 
+ bl[149] br[149] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_152 
+ bl[150] br[150] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_153 
+ bl[151] br[151] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_154 
+ bl[152] br[152] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_155 
+ bl[153] br[153] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_156 
+ bl[154] br[154] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_157 
+ bl[155] br[155] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_158 
+ bl[156] br[156] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_159 
+ bl[157] br[157] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_160 
+ bl[158] br[158] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_161 
+ bl[159] br[159] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_162 
+ bl[160] br[160] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_163 
+ bl[161] br[161] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_164 
+ bl[162] br[162] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_165 
+ bl[163] br[163] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_166 
+ bl[164] br[164] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_167 
+ bl[165] br[165] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_168 
+ bl[166] br[166] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_169 
+ bl[167] br[167] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_170 
+ bl[168] br[168] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_171 
+ bl[169] br[169] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_172 
+ bl[170] br[170] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_173 
+ bl[171] br[171] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_174 
+ bl[172] br[172] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_175 
+ bl[173] br[173] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_176 
+ bl[174] br[174] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_177 
+ bl[175] br[175] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_178 
+ bl[176] br[176] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_179 
+ bl[177] br[177] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_180 
+ bl[178] br[178] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_181 
+ bl[179] br[179] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_182 
+ bl[180] br[180] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_183 
+ bl[181] br[181] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_184 
+ bl[182] br[182] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_185 
+ bl[183] br[183] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_186 
+ bl[184] br[184] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_187 
+ bl[185] br[185] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_188 
+ bl[186] br[186] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_189 
+ bl[187] br[187] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_190 
+ bl[188] br[188] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_191 
+ bl[189] br[189] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_192 
+ bl[190] br[190] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_193 
+ bl[191] br[191] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_194 
+ bl[192] br[192] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_195 
+ bl[193] br[193] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_196 
+ bl[194] br[194] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_197 
+ bl[195] br[195] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_198 
+ bl[196] br[196] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_199 
+ bl[197] br[197] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_200 
+ bl[198] br[198] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_201 
+ bl[199] br[199] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_202 
+ bl[200] br[200] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_203 
+ bl[201] br[201] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_204 
+ bl[202] br[202] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_205 
+ bl[203] br[203] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_206 
+ bl[204] br[204] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_207 
+ bl[205] br[205] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_208 
+ bl[206] br[206] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_209 
+ bl[207] br[207] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_210 
+ bl[208] br[208] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_211 
+ bl[209] br[209] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_212 
+ bl[210] br[210] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_213 
+ bl[211] br[211] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_214 
+ bl[212] br[212] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_215 
+ bl[213] br[213] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_216 
+ bl[214] br[214] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_217 
+ bl[215] br[215] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_218 
+ bl[216] br[216] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_219 
+ bl[217] br[217] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_220 
+ bl[218] br[218] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_221 
+ bl[219] br[219] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_222 
+ bl[220] br[220] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_223 
+ bl[221] br[221] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_224 
+ bl[222] br[222] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_225 
+ bl[223] br[223] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_226 
+ bl[224] br[224] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_227 
+ bl[225] br[225] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_228 
+ bl[226] br[226] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_229 
+ bl[227] br[227] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_230 
+ bl[228] br[228] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_231 
+ bl[229] br[229] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_232 
+ bl[230] br[230] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_233 
+ bl[231] br[231] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_234 
+ bl[232] br[232] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_235 
+ bl[233] br[233] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_236 
+ bl[234] br[234] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_237 
+ bl[235] br[235] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_238 
+ bl[236] br[236] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_239 
+ bl[237] br[237] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_240 
+ bl[238] br[238] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_241 
+ bl[239] br[239] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_242 
+ bl[240] br[240] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_243 
+ bl[241] br[241] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_244 
+ bl[242] br[242] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_245 
+ bl[243] br[243] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_246 
+ bl[244] br[244] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_247 
+ bl[245] br[245] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_248 
+ bl[246] br[246] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_249 
+ bl[247] br[247] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_250 
+ bl[248] br[248] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_251 
+ bl[249] br[249] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_252 
+ bl[250] br[250] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_253 
+ bl[251] br[251] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_254 
+ bl[252] br[252] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_255 
+ bl[253] br[253] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_256 
+ bl[254] br[254] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_257 
+ bl[255] br[255] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_258 
+ vdd vdd vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_259 
+ vdd vdd vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_0 
+ vdd vdd vss vdd vpb vnb wl[26] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_28_1 
+ rbl rbr vss vdd vpb vnb wl[26] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_28_2 
+ bl[0] br[0] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_3 
+ bl[1] br[1] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_4 
+ bl[2] br[2] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_5 
+ bl[3] br[3] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_6 
+ bl[4] br[4] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_7 
+ bl[5] br[5] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_8 
+ bl[6] br[6] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_9 
+ bl[7] br[7] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_10 
+ bl[8] br[8] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_11 
+ bl[9] br[9] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_12 
+ bl[10] br[10] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_13 
+ bl[11] br[11] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_14 
+ bl[12] br[12] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_15 
+ bl[13] br[13] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_16 
+ bl[14] br[14] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_17 
+ bl[15] br[15] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_18 
+ bl[16] br[16] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_19 
+ bl[17] br[17] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_20 
+ bl[18] br[18] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_21 
+ bl[19] br[19] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_22 
+ bl[20] br[20] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_23 
+ bl[21] br[21] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_24 
+ bl[22] br[22] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_25 
+ bl[23] br[23] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_26 
+ bl[24] br[24] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_27 
+ bl[25] br[25] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_28 
+ bl[26] br[26] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_29 
+ bl[27] br[27] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_30 
+ bl[28] br[28] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_31 
+ bl[29] br[29] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_32 
+ bl[30] br[30] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_33 
+ bl[31] br[31] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_34 
+ bl[32] br[32] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_35 
+ bl[33] br[33] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_36 
+ bl[34] br[34] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_37 
+ bl[35] br[35] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_38 
+ bl[36] br[36] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_39 
+ bl[37] br[37] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_40 
+ bl[38] br[38] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_41 
+ bl[39] br[39] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_42 
+ bl[40] br[40] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_43 
+ bl[41] br[41] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_44 
+ bl[42] br[42] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_45 
+ bl[43] br[43] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_46 
+ bl[44] br[44] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_47 
+ bl[45] br[45] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_48 
+ bl[46] br[46] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_49 
+ bl[47] br[47] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_50 
+ bl[48] br[48] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_51 
+ bl[49] br[49] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_52 
+ bl[50] br[50] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_53 
+ bl[51] br[51] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_54 
+ bl[52] br[52] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_55 
+ bl[53] br[53] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_56 
+ bl[54] br[54] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_57 
+ bl[55] br[55] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_58 
+ bl[56] br[56] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_59 
+ bl[57] br[57] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_60 
+ bl[58] br[58] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_61 
+ bl[59] br[59] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_62 
+ bl[60] br[60] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_63 
+ bl[61] br[61] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_64 
+ bl[62] br[62] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_65 
+ bl[63] br[63] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_66 
+ bl[64] br[64] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_67 
+ bl[65] br[65] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_68 
+ bl[66] br[66] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_69 
+ bl[67] br[67] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_70 
+ bl[68] br[68] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_71 
+ bl[69] br[69] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_72 
+ bl[70] br[70] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_73 
+ bl[71] br[71] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_74 
+ bl[72] br[72] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_75 
+ bl[73] br[73] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_76 
+ bl[74] br[74] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_77 
+ bl[75] br[75] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_78 
+ bl[76] br[76] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_79 
+ bl[77] br[77] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_80 
+ bl[78] br[78] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_81 
+ bl[79] br[79] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_82 
+ bl[80] br[80] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_83 
+ bl[81] br[81] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_84 
+ bl[82] br[82] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_85 
+ bl[83] br[83] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_86 
+ bl[84] br[84] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_87 
+ bl[85] br[85] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_88 
+ bl[86] br[86] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_89 
+ bl[87] br[87] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_90 
+ bl[88] br[88] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_91 
+ bl[89] br[89] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_92 
+ bl[90] br[90] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_93 
+ bl[91] br[91] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_94 
+ bl[92] br[92] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_95 
+ bl[93] br[93] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_96 
+ bl[94] br[94] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_97 
+ bl[95] br[95] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_98 
+ bl[96] br[96] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_99 
+ bl[97] br[97] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_100 
+ bl[98] br[98] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_101 
+ bl[99] br[99] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_102 
+ bl[100] br[100] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_103 
+ bl[101] br[101] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_104 
+ bl[102] br[102] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_105 
+ bl[103] br[103] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_106 
+ bl[104] br[104] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_107 
+ bl[105] br[105] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_108 
+ bl[106] br[106] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_109 
+ bl[107] br[107] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_110 
+ bl[108] br[108] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_111 
+ bl[109] br[109] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_112 
+ bl[110] br[110] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_113 
+ bl[111] br[111] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_114 
+ bl[112] br[112] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_115 
+ bl[113] br[113] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_116 
+ bl[114] br[114] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_117 
+ bl[115] br[115] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_118 
+ bl[116] br[116] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_119 
+ bl[117] br[117] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_120 
+ bl[118] br[118] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_121 
+ bl[119] br[119] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_122 
+ bl[120] br[120] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_123 
+ bl[121] br[121] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_124 
+ bl[122] br[122] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_125 
+ bl[123] br[123] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_126 
+ bl[124] br[124] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_127 
+ bl[125] br[125] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_128 
+ bl[126] br[126] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_129 
+ bl[127] br[127] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_130 
+ bl[128] br[128] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_131 
+ bl[129] br[129] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_132 
+ bl[130] br[130] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_133 
+ bl[131] br[131] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_134 
+ bl[132] br[132] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_135 
+ bl[133] br[133] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_136 
+ bl[134] br[134] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_137 
+ bl[135] br[135] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_138 
+ bl[136] br[136] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_139 
+ bl[137] br[137] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_140 
+ bl[138] br[138] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_141 
+ bl[139] br[139] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_142 
+ bl[140] br[140] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_143 
+ bl[141] br[141] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_144 
+ bl[142] br[142] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_145 
+ bl[143] br[143] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_146 
+ bl[144] br[144] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_147 
+ bl[145] br[145] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_148 
+ bl[146] br[146] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_149 
+ bl[147] br[147] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_150 
+ bl[148] br[148] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_151 
+ bl[149] br[149] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_152 
+ bl[150] br[150] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_153 
+ bl[151] br[151] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_154 
+ bl[152] br[152] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_155 
+ bl[153] br[153] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_156 
+ bl[154] br[154] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_157 
+ bl[155] br[155] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_158 
+ bl[156] br[156] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_159 
+ bl[157] br[157] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_160 
+ bl[158] br[158] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_161 
+ bl[159] br[159] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_162 
+ bl[160] br[160] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_163 
+ bl[161] br[161] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_164 
+ bl[162] br[162] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_165 
+ bl[163] br[163] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_166 
+ bl[164] br[164] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_167 
+ bl[165] br[165] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_168 
+ bl[166] br[166] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_169 
+ bl[167] br[167] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_170 
+ bl[168] br[168] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_171 
+ bl[169] br[169] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_172 
+ bl[170] br[170] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_173 
+ bl[171] br[171] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_174 
+ bl[172] br[172] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_175 
+ bl[173] br[173] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_176 
+ bl[174] br[174] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_177 
+ bl[175] br[175] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_178 
+ bl[176] br[176] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_179 
+ bl[177] br[177] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_180 
+ bl[178] br[178] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_181 
+ bl[179] br[179] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_182 
+ bl[180] br[180] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_183 
+ bl[181] br[181] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_184 
+ bl[182] br[182] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_185 
+ bl[183] br[183] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_186 
+ bl[184] br[184] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_187 
+ bl[185] br[185] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_188 
+ bl[186] br[186] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_189 
+ bl[187] br[187] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_190 
+ bl[188] br[188] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_191 
+ bl[189] br[189] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_192 
+ bl[190] br[190] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_193 
+ bl[191] br[191] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_194 
+ bl[192] br[192] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_195 
+ bl[193] br[193] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_196 
+ bl[194] br[194] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_197 
+ bl[195] br[195] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_198 
+ bl[196] br[196] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_199 
+ bl[197] br[197] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_200 
+ bl[198] br[198] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_201 
+ bl[199] br[199] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_202 
+ bl[200] br[200] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_203 
+ bl[201] br[201] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_204 
+ bl[202] br[202] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_205 
+ bl[203] br[203] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_206 
+ bl[204] br[204] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_207 
+ bl[205] br[205] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_208 
+ bl[206] br[206] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_209 
+ bl[207] br[207] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_210 
+ bl[208] br[208] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_211 
+ bl[209] br[209] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_212 
+ bl[210] br[210] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_213 
+ bl[211] br[211] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_214 
+ bl[212] br[212] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_215 
+ bl[213] br[213] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_216 
+ bl[214] br[214] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_217 
+ bl[215] br[215] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_218 
+ bl[216] br[216] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_219 
+ bl[217] br[217] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_220 
+ bl[218] br[218] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_221 
+ bl[219] br[219] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_222 
+ bl[220] br[220] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_223 
+ bl[221] br[221] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_224 
+ bl[222] br[222] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_225 
+ bl[223] br[223] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_226 
+ bl[224] br[224] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_227 
+ bl[225] br[225] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_228 
+ bl[226] br[226] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_229 
+ bl[227] br[227] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_230 
+ bl[228] br[228] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_231 
+ bl[229] br[229] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_232 
+ bl[230] br[230] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_233 
+ bl[231] br[231] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_234 
+ bl[232] br[232] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_235 
+ bl[233] br[233] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_236 
+ bl[234] br[234] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_237 
+ bl[235] br[235] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_238 
+ bl[236] br[236] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_239 
+ bl[237] br[237] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_240 
+ bl[238] br[238] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_241 
+ bl[239] br[239] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_242 
+ bl[240] br[240] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_243 
+ bl[241] br[241] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_244 
+ bl[242] br[242] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_245 
+ bl[243] br[243] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_246 
+ bl[244] br[244] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_247 
+ bl[245] br[245] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_248 
+ bl[246] br[246] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_249 
+ bl[247] br[247] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_250 
+ bl[248] br[248] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_251 
+ bl[249] br[249] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_252 
+ bl[250] br[250] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_253 
+ bl[251] br[251] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_254 
+ bl[252] br[252] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_255 
+ bl[253] br[253] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_256 
+ bl[254] br[254] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_257 
+ bl[255] br[255] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_258 
+ vdd vdd vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_259 
+ vdd vdd vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_0 
+ vdd vdd vss vdd vpb vnb wl[27] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_29_1 
+ rbl rbr vss vdd vpb vnb wl[27] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_29_2 
+ bl[0] br[0] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_3 
+ bl[1] br[1] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_4 
+ bl[2] br[2] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_5 
+ bl[3] br[3] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_6 
+ bl[4] br[4] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_7 
+ bl[5] br[5] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_8 
+ bl[6] br[6] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_9 
+ bl[7] br[7] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_10 
+ bl[8] br[8] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_11 
+ bl[9] br[9] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_12 
+ bl[10] br[10] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_13 
+ bl[11] br[11] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_14 
+ bl[12] br[12] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_15 
+ bl[13] br[13] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_16 
+ bl[14] br[14] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_17 
+ bl[15] br[15] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_18 
+ bl[16] br[16] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_19 
+ bl[17] br[17] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_20 
+ bl[18] br[18] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_21 
+ bl[19] br[19] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_22 
+ bl[20] br[20] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_23 
+ bl[21] br[21] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_24 
+ bl[22] br[22] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_25 
+ bl[23] br[23] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_26 
+ bl[24] br[24] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_27 
+ bl[25] br[25] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_28 
+ bl[26] br[26] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_29 
+ bl[27] br[27] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_30 
+ bl[28] br[28] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_31 
+ bl[29] br[29] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_32 
+ bl[30] br[30] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_33 
+ bl[31] br[31] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_34 
+ bl[32] br[32] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_35 
+ bl[33] br[33] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_36 
+ bl[34] br[34] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_37 
+ bl[35] br[35] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_38 
+ bl[36] br[36] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_39 
+ bl[37] br[37] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_40 
+ bl[38] br[38] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_41 
+ bl[39] br[39] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_42 
+ bl[40] br[40] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_43 
+ bl[41] br[41] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_44 
+ bl[42] br[42] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_45 
+ bl[43] br[43] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_46 
+ bl[44] br[44] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_47 
+ bl[45] br[45] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_48 
+ bl[46] br[46] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_49 
+ bl[47] br[47] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_50 
+ bl[48] br[48] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_51 
+ bl[49] br[49] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_52 
+ bl[50] br[50] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_53 
+ bl[51] br[51] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_54 
+ bl[52] br[52] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_55 
+ bl[53] br[53] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_56 
+ bl[54] br[54] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_57 
+ bl[55] br[55] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_58 
+ bl[56] br[56] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_59 
+ bl[57] br[57] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_60 
+ bl[58] br[58] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_61 
+ bl[59] br[59] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_62 
+ bl[60] br[60] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_63 
+ bl[61] br[61] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_64 
+ bl[62] br[62] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_65 
+ bl[63] br[63] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_66 
+ bl[64] br[64] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_67 
+ bl[65] br[65] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_68 
+ bl[66] br[66] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_69 
+ bl[67] br[67] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_70 
+ bl[68] br[68] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_71 
+ bl[69] br[69] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_72 
+ bl[70] br[70] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_73 
+ bl[71] br[71] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_74 
+ bl[72] br[72] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_75 
+ bl[73] br[73] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_76 
+ bl[74] br[74] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_77 
+ bl[75] br[75] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_78 
+ bl[76] br[76] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_79 
+ bl[77] br[77] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_80 
+ bl[78] br[78] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_81 
+ bl[79] br[79] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_82 
+ bl[80] br[80] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_83 
+ bl[81] br[81] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_84 
+ bl[82] br[82] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_85 
+ bl[83] br[83] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_86 
+ bl[84] br[84] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_87 
+ bl[85] br[85] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_88 
+ bl[86] br[86] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_89 
+ bl[87] br[87] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_90 
+ bl[88] br[88] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_91 
+ bl[89] br[89] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_92 
+ bl[90] br[90] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_93 
+ bl[91] br[91] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_94 
+ bl[92] br[92] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_95 
+ bl[93] br[93] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_96 
+ bl[94] br[94] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_97 
+ bl[95] br[95] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_98 
+ bl[96] br[96] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_99 
+ bl[97] br[97] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_100 
+ bl[98] br[98] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_101 
+ bl[99] br[99] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_102 
+ bl[100] br[100] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_103 
+ bl[101] br[101] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_104 
+ bl[102] br[102] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_105 
+ bl[103] br[103] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_106 
+ bl[104] br[104] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_107 
+ bl[105] br[105] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_108 
+ bl[106] br[106] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_109 
+ bl[107] br[107] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_110 
+ bl[108] br[108] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_111 
+ bl[109] br[109] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_112 
+ bl[110] br[110] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_113 
+ bl[111] br[111] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_114 
+ bl[112] br[112] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_115 
+ bl[113] br[113] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_116 
+ bl[114] br[114] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_117 
+ bl[115] br[115] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_118 
+ bl[116] br[116] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_119 
+ bl[117] br[117] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_120 
+ bl[118] br[118] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_121 
+ bl[119] br[119] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_122 
+ bl[120] br[120] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_123 
+ bl[121] br[121] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_124 
+ bl[122] br[122] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_125 
+ bl[123] br[123] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_126 
+ bl[124] br[124] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_127 
+ bl[125] br[125] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_128 
+ bl[126] br[126] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_129 
+ bl[127] br[127] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_130 
+ bl[128] br[128] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_131 
+ bl[129] br[129] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_132 
+ bl[130] br[130] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_133 
+ bl[131] br[131] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_134 
+ bl[132] br[132] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_135 
+ bl[133] br[133] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_136 
+ bl[134] br[134] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_137 
+ bl[135] br[135] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_138 
+ bl[136] br[136] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_139 
+ bl[137] br[137] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_140 
+ bl[138] br[138] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_141 
+ bl[139] br[139] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_142 
+ bl[140] br[140] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_143 
+ bl[141] br[141] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_144 
+ bl[142] br[142] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_145 
+ bl[143] br[143] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_146 
+ bl[144] br[144] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_147 
+ bl[145] br[145] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_148 
+ bl[146] br[146] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_149 
+ bl[147] br[147] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_150 
+ bl[148] br[148] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_151 
+ bl[149] br[149] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_152 
+ bl[150] br[150] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_153 
+ bl[151] br[151] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_154 
+ bl[152] br[152] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_155 
+ bl[153] br[153] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_156 
+ bl[154] br[154] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_157 
+ bl[155] br[155] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_158 
+ bl[156] br[156] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_159 
+ bl[157] br[157] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_160 
+ bl[158] br[158] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_161 
+ bl[159] br[159] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_162 
+ bl[160] br[160] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_163 
+ bl[161] br[161] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_164 
+ bl[162] br[162] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_165 
+ bl[163] br[163] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_166 
+ bl[164] br[164] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_167 
+ bl[165] br[165] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_168 
+ bl[166] br[166] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_169 
+ bl[167] br[167] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_170 
+ bl[168] br[168] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_171 
+ bl[169] br[169] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_172 
+ bl[170] br[170] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_173 
+ bl[171] br[171] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_174 
+ bl[172] br[172] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_175 
+ bl[173] br[173] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_176 
+ bl[174] br[174] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_177 
+ bl[175] br[175] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_178 
+ bl[176] br[176] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_179 
+ bl[177] br[177] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_180 
+ bl[178] br[178] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_181 
+ bl[179] br[179] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_182 
+ bl[180] br[180] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_183 
+ bl[181] br[181] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_184 
+ bl[182] br[182] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_185 
+ bl[183] br[183] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_186 
+ bl[184] br[184] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_187 
+ bl[185] br[185] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_188 
+ bl[186] br[186] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_189 
+ bl[187] br[187] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_190 
+ bl[188] br[188] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_191 
+ bl[189] br[189] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_192 
+ bl[190] br[190] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_193 
+ bl[191] br[191] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_194 
+ bl[192] br[192] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_195 
+ bl[193] br[193] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_196 
+ bl[194] br[194] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_197 
+ bl[195] br[195] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_198 
+ bl[196] br[196] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_199 
+ bl[197] br[197] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_200 
+ bl[198] br[198] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_201 
+ bl[199] br[199] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_202 
+ bl[200] br[200] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_203 
+ bl[201] br[201] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_204 
+ bl[202] br[202] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_205 
+ bl[203] br[203] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_206 
+ bl[204] br[204] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_207 
+ bl[205] br[205] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_208 
+ bl[206] br[206] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_209 
+ bl[207] br[207] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_210 
+ bl[208] br[208] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_211 
+ bl[209] br[209] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_212 
+ bl[210] br[210] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_213 
+ bl[211] br[211] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_214 
+ bl[212] br[212] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_215 
+ bl[213] br[213] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_216 
+ bl[214] br[214] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_217 
+ bl[215] br[215] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_218 
+ bl[216] br[216] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_219 
+ bl[217] br[217] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_220 
+ bl[218] br[218] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_221 
+ bl[219] br[219] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_222 
+ bl[220] br[220] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_223 
+ bl[221] br[221] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_224 
+ bl[222] br[222] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_225 
+ bl[223] br[223] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_226 
+ bl[224] br[224] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_227 
+ bl[225] br[225] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_228 
+ bl[226] br[226] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_229 
+ bl[227] br[227] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_230 
+ bl[228] br[228] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_231 
+ bl[229] br[229] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_232 
+ bl[230] br[230] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_233 
+ bl[231] br[231] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_234 
+ bl[232] br[232] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_235 
+ bl[233] br[233] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_236 
+ bl[234] br[234] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_237 
+ bl[235] br[235] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_238 
+ bl[236] br[236] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_239 
+ bl[237] br[237] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_240 
+ bl[238] br[238] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_241 
+ bl[239] br[239] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_242 
+ bl[240] br[240] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_243 
+ bl[241] br[241] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_244 
+ bl[242] br[242] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_245 
+ bl[243] br[243] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_246 
+ bl[244] br[244] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_247 
+ bl[245] br[245] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_248 
+ bl[246] br[246] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_249 
+ bl[247] br[247] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_250 
+ bl[248] br[248] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_251 
+ bl[249] br[249] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_252 
+ bl[250] br[250] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_253 
+ bl[251] br[251] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_254 
+ bl[252] br[252] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_255 
+ bl[253] br[253] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_256 
+ bl[254] br[254] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_257 
+ bl[255] br[255] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_258 
+ vdd vdd vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_259 
+ vdd vdd vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_0 
+ vdd vdd vss vdd vpb vnb wl[28] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_30_1 
+ rbl rbr vss vdd vpb vnb wl[28] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_30_2 
+ bl[0] br[0] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_3 
+ bl[1] br[1] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_4 
+ bl[2] br[2] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_5 
+ bl[3] br[3] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_6 
+ bl[4] br[4] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_7 
+ bl[5] br[5] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_8 
+ bl[6] br[6] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_9 
+ bl[7] br[7] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_10 
+ bl[8] br[8] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_11 
+ bl[9] br[9] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_12 
+ bl[10] br[10] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_13 
+ bl[11] br[11] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_14 
+ bl[12] br[12] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_15 
+ bl[13] br[13] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_16 
+ bl[14] br[14] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_17 
+ bl[15] br[15] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_18 
+ bl[16] br[16] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_19 
+ bl[17] br[17] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_20 
+ bl[18] br[18] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_21 
+ bl[19] br[19] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_22 
+ bl[20] br[20] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_23 
+ bl[21] br[21] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_24 
+ bl[22] br[22] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_25 
+ bl[23] br[23] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_26 
+ bl[24] br[24] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_27 
+ bl[25] br[25] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_28 
+ bl[26] br[26] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_29 
+ bl[27] br[27] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_30 
+ bl[28] br[28] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_31 
+ bl[29] br[29] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_32 
+ bl[30] br[30] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_33 
+ bl[31] br[31] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_34 
+ bl[32] br[32] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_35 
+ bl[33] br[33] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_36 
+ bl[34] br[34] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_37 
+ bl[35] br[35] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_38 
+ bl[36] br[36] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_39 
+ bl[37] br[37] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_40 
+ bl[38] br[38] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_41 
+ bl[39] br[39] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_42 
+ bl[40] br[40] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_43 
+ bl[41] br[41] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_44 
+ bl[42] br[42] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_45 
+ bl[43] br[43] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_46 
+ bl[44] br[44] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_47 
+ bl[45] br[45] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_48 
+ bl[46] br[46] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_49 
+ bl[47] br[47] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_50 
+ bl[48] br[48] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_51 
+ bl[49] br[49] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_52 
+ bl[50] br[50] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_53 
+ bl[51] br[51] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_54 
+ bl[52] br[52] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_55 
+ bl[53] br[53] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_56 
+ bl[54] br[54] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_57 
+ bl[55] br[55] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_58 
+ bl[56] br[56] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_59 
+ bl[57] br[57] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_60 
+ bl[58] br[58] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_61 
+ bl[59] br[59] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_62 
+ bl[60] br[60] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_63 
+ bl[61] br[61] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_64 
+ bl[62] br[62] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_65 
+ bl[63] br[63] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_66 
+ bl[64] br[64] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_67 
+ bl[65] br[65] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_68 
+ bl[66] br[66] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_69 
+ bl[67] br[67] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_70 
+ bl[68] br[68] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_71 
+ bl[69] br[69] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_72 
+ bl[70] br[70] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_73 
+ bl[71] br[71] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_74 
+ bl[72] br[72] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_75 
+ bl[73] br[73] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_76 
+ bl[74] br[74] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_77 
+ bl[75] br[75] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_78 
+ bl[76] br[76] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_79 
+ bl[77] br[77] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_80 
+ bl[78] br[78] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_81 
+ bl[79] br[79] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_82 
+ bl[80] br[80] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_83 
+ bl[81] br[81] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_84 
+ bl[82] br[82] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_85 
+ bl[83] br[83] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_86 
+ bl[84] br[84] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_87 
+ bl[85] br[85] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_88 
+ bl[86] br[86] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_89 
+ bl[87] br[87] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_90 
+ bl[88] br[88] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_91 
+ bl[89] br[89] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_92 
+ bl[90] br[90] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_93 
+ bl[91] br[91] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_94 
+ bl[92] br[92] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_95 
+ bl[93] br[93] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_96 
+ bl[94] br[94] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_97 
+ bl[95] br[95] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_98 
+ bl[96] br[96] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_99 
+ bl[97] br[97] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_100 
+ bl[98] br[98] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_101 
+ bl[99] br[99] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_102 
+ bl[100] br[100] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_103 
+ bl[101] br[101] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_104 
+ bl[102] br[102] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_105 
+ bl[103] br[103] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_106 
+ bl[104] br[104] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_107 
+ bl[105] br[105] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_108 
+ bl[106] br[106] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_109 
+ bl[107] br[107] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_110 
+ bl[108] br[108] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_111 
+ bl[109] br[109] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_112 
+ bl[110] br[110] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_113 
+ bl[111] br[111] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_114 
+ bl[112] br[112] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_115 
+ bl[113] br[113] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_116 
+ bl[114] br[114] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_117 
+ bl[115] br[115] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_118 
+ bl[116] br[116] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_119 
+ bl[117] br[117] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_120 
+ bl[118] br[118] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_121 
+ bl[119] br[119] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_122 
+ bl[120] br[120] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_123 
+ bl[121] br[121] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_124 
+ bl[122] br[122] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_125 
+ bl[123] br[123] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_126 
+ bl[124] br[124] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_127 
+ bl[125] br[125] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_128 
+ bl[126] br[126] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_129 
+ bl[127] br[127] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_130 
+ bl[128] br[128] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_131 
+ bl[129] br[129] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_132 
+ bl[130] br[130] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_133 
+ bl[131] br[131] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_134 
+ bl[132] br[132] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_135 
+ bl[133] br[133] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_136 
+ bl[134] br[134] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_137 
+ bl[135] br[135] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_138 
+ bl[136] br[136] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_139 
+ bl[137] br[137] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_140 
+ bl[138] br[138] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_141 
+ bl[139] br[139] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_142 
+ bl[140] br[140] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_143 
+ bl[141] br[141] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_144 
+ bl[142] br[142] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_145 
+ bl[143] br[143] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_146 
+ bl[144] br[144] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_147 
+ bl[145] br[145] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_148 
+ bl[146] br[146] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_149 
+ bl[147] br[147] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_150 
+ bl[148] br[148] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_151 
+ bl[149] br[149] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_152 
+ bl[150] br[150] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_153 
+ bl[151] br[151] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_154 
+ bl[152] br[152] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_155 
+ bl[153] br[153] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_156 
+ bl[154] br[154] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_157 
+ bl[155] br[155] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_158 
+ bl[156] br[156] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_159 
+ bl[157] br[157] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_160 
+ bl[158] br[158] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_161 
+ bl[159] br[159] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_162 
+ bl[160] br[160] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_163 
+ bl[161] br[161] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_164 
+ bl[162] br[162] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_165 
+ bl[163] br[163] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_166 
+ bl[164] br[164] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_167 
+ bl[165] br[165] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_168 
+ bl[166] br[166] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_169 
+ bl[167] br[167] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_170 
+ bl[168] br[168] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_171 
+ bl[169] br[169] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_172 
+ bl[170] br[170] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_173 
+ bl[171] br[171] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_174 
+ bl[172] br[172] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_175 
+ bl[173] br[173] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_176 
+ bl[174] br[174] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_177 
+ bl[175] br[175] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_178 
+ bl[176] br[176] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_179 
+ bl[177] br[177] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_180 
+ bl[178] br[178] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_181 
+ bl[179] br[179] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_182 
+ bl[180] br[180] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_183 
+ bl[181] br[181] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_184 
+ bl[182] br[182] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_185 
+ bl[183] br[183] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_186 
+ bl[184] br[184] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_187 
+ bl[185] br[185] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_188 
+ bl[186] br[186] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_189 
+ bl[187] br[187] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_190 
+ bl[188] br[188] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_191 
+ bl[189] br[189] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_192 
+ bl[190] br[190] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_193 
+ bl[191] br[191] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_194 
+ bl[192] br[192] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_195 
+ bl[193] br[193] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_196 
+ bl[194] br[194] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_197 
+ bl[195] br[195] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_198 
+ bl[196] br[196] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_199 
+ bl[197] br[197] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_200 
+ bl[198] br[198] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_201 
+ bl[199] br[199] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_202 
+ bl[200] br[200] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_203 
+ bl[201] br[201] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_204 
+ bl[202] br[202] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_205 
+ bl[203] br[203] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_206 
+ bl[204] br[204] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_207 
+ bl[205] br[205] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_208 
+ bl[206] br[206] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_209 
+ bl[207] br[207] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_210 
+ bl[208] br[208] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_211 
+ bl[209] br[209] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_212 
+ bl[210] br[210] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_213 
+ bl[211] br[211] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_214 
+ bl[212] br[212] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_215 
+ bl[213] br[213] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_216 
+ bl[214] br[214] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_217 
+ bl[215] br[215] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_218 
+ bl[216] br[216] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_219 
+ bl[217] br[217] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_220 
+ bl[218] br[218] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_221 
+ bl[219] br[219] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_222 
+ bl[220] br[220] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_223 
+ bl[221] br[221] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_224 
+ bl[222] br[222] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_225 
+ bl[223] br[223] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_226 
+ bl[224] br[224] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_227 
+ bl[225] br[225] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_228 
+ bl[226] br[226] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_229 
+ bl[227] br[227] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_230 
+ bl[228] br[228] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_231 
+ bl[229] br[229] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_232 
+ bl[230] br[230] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_233 
+ bl[231] br[231] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_234 
+ bl[232] br[232] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_235 
+ bl[233] br[233] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_236 
+ bl[234] br[234] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_237 
+ bl[235] br[235] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_238 
+ bl[236] br[236] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_239 
+ bl[237] br[237] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_240 
+ bl[238] br[238] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_241 
+ bl[239] br[239] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_242 
+ bl[240] br[240] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_243 
+ bl[241] br[241] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_244 
+ bl[242] br[242] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_245 
+ bl[243] br[243] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_246 
+ bl[244] br[244] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_247 
+ bl[245] br[245] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_248 
+ bl[246] br[246] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_249 
+ bl[247] br[247] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_250 
+ bl[248] br[248] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_251 
+ bl[249] br[249] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_252 
+ bl[250] br[250] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_253 
+ bl[251] br[251] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_254 
+ bl[252] br[252] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_255 
+ bl[253] br[253] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_256 
+ bl[254] br[254] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_257 
+ bl[255] br[255] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_258 
+ vdd vdd vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_259 
+ vdd vdd vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_0 
+ vdd vdd vss vdd vpb vnb wl[29] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_31_1 
+ rbl rbr vss vdd vpb vnb wl[29] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_31_2 
+ bl[0] br[0] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_3 
+ bl[1] br[1] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_4 
+ bl[2] br[2] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_5 
+ bl[3] br[3] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_6 
+ bl[4] br[4] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_7 
+ bl[5] br[5] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_8 
+ bl[6] br[6] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_9 
+ bl[7] br[7] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_10 
+ bl[8] br[8] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_11 
+ bl[9] br[9] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_12 
+ bl[10] br[10] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_13 
+ bl[11] br[11] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_14 
+ bl[12] br[12] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_15 
+ bl[13] br[13] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_16 
+ bl[14] br[14] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_17 
+ bl[15] br[15] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_18 
+ bl[16] br[16] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_19 
+ bl[17] br[17] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_20 
+ bl[18] br[18] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_21 
+ bl[19] br[19] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_22 
+ bl[20] br[20] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_23 
+ bl[21] br[21] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_24 
+ bl[22] br[22] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_25 
+ bl[23] br[23] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_26 
+ bl[24] br[24] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_27 
+ bl[25] br[25] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_28 
+ bl[26] br[26] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_29 
+ bl[27] br[27] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_30 
+ bl[28] br[28] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_31 
+ bl[29] br[29] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_32 
+ bl[30] br[30] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_33 
+ bl[31] br[31] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_34 
+ bl[32] br[32] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_35 
+ bl[33] br[33] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_36 
+ bl[34] br[34] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_37 
+ bl[35] br[35] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_38 
+ bl[36] br[36] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_39 
+ bl[37] br[37] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_40 
+ bl[38] br[38] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_41 
+ bl[39] br[39] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_42 
+ bl[40] br[40] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_43 
+ bl[41] br[41] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_44 
+ bl[42] br[42] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_45 
+ bl[43] br[43] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_46 
+ bl[44] br[44] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_47 
+ bl[45] br[45] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_48 
+ bl[46] br[46] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_49 
+ bl[47] br[47] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_50 
+ bl[48] br[48] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_51 
+ bl[49] br[49] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_52 
+ bl[50] br[50] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_53 
+ bl[51] br[51] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_54 
+ bl[52] br[52] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_55 
+ bl[53] br[53] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_56 
+ bl[54] br[54] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_57 
+ bl[55] br[55] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_58 
+ bl[56] br[56] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_59 
+ bl[57] br[57] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_60 
+ bl[58] br[58] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_61 
+ bl[59] br[59] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_62 
+ bl[60] br[60] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_63 
+ bl[61] br[61] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_64 
+ bl[62] br[62] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_65 
+ bl[63] br[63] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_66 
+ bl[64] br[64] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_67 
+ bl[65] br[65] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_68 
+ bl[66] br[66] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_69 
+ bl[67] br[67] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_70 
+ bl[68] br[68] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_71 
+ bl[69] br[69] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_72 
+ bl[70] br[70] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_73 
+ bl[71] br[71] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_74 
+ bl[72] br[72] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_75 
+ bl[73] br[73] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_76 
+ bl[74] br[74] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_77 
+ bl[75] br[75] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_78 
+ bl[76] br[76] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_79 
+ bl[77] br[77] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_80 
+ bl[78] br[78] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_81 
+ bl[79] br[79] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_82 
+ bl[80] br[80] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_83 
+ bl[81] br[81] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_84 
+ bl[82] br[82] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_85 
+ bl[83] br[83] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_86 
+ bl[84] br[84] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_87 
+ bl[85] br[85] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_88 
+ bl[86] br[86] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_89 
+ bl[87] br[87] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_90 
+ bl[88] br[88] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_91 
+ bl[89] br[89] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_92 
+ bl[90] br[90] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_93 
+ bl[91] br[91] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_94 
+ bl[92] br[92] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_95 
+ bl[93] br[93] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_96 
+ bl[94] br[94] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_97 
+ bl[95] br[95] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_98 
+ bl[96] br[96] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_99 
+ bl[97] br[97] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_100 
+ bl[98] br[98] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_101 
+ bl[99] br[99] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_102 
+ bl[100] br[100] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_103 
+ bl[101] br[101] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_104 
+ bl[102] br[102] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_105 
+ bl[103] br[103] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_106 
+ bl[104] br[104] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_107 
+ bl[105] br[105] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_108 
+ bl[106] br[106] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_109 
+ bl[107] br[107] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_110 
+ bl[108] br[108] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_111 
+ bl[109] br[109] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_112 
+ bl[110] br[110] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_113 
+ bl[111] br[111] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_114 
+ bl[112] br[112] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_115 
+ bl[113] br[113] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_116 
+ bl[114] br[114] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_117 
+ bl[115] br[115] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_118 
+ bl[116] br[116] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_119 
+ bl[117] br[117] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_120 
+ bl[118] br[118] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_121 
+ bl[119] br[119] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_122 
+ bl[120] br[120] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_123 
+ bl[121] br[121] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_124 
+ bl[122] br[122] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_125 
+ bl[123] br[123] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_126 
+ bl[124] br[124] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_127 
+ bl[125] br[125] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_128 
+ bl[126] br[126] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_129 
+ bl[127] br[127] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_130 
+ bl[128] br[128] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_131 
+ bl[129] br[129] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_132 
+ bl[130] br[130] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_133 
+ bl[131] br[131] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_134 
+ bl[132] br[132] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_135 
+ bl[133] br[133] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_136 
+ bl[134] br[134] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_137 
+ bl[135] br[135] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_138 
+ bl[136] br[136] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_139 
+ bl[137] br[137] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_140 
+ bl[138] br[138] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_141 
+ bl[139] br[139] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_142 
+ bl[140] br[140] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_143 
+ bl[141] br[141] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_144 
+ bl[142] br[142] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_145 
+ bl[143] br[143] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_146 
+ bl[144] br[144] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_147 
+ bl[145] br[145] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_148 
+ bl[146] br[146] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_149 
+ bl[147] br[147] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_150 
+ bl[148] br[148] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_151 
+ bl[149] br[149] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_152 
+ bl[150] br[150] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_153 
+ bl[151] br[151] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_154 
+ bl[152] br[152] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_155 
+ bl[153] br[153] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_156 
+ bl[154] br[154] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_157 
+ bl[155] br[155] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_158 
+ bl[156] br[156] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_159 
+ bl[157] br[157] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_160 
+ bl[158] br[158] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_161 
+ bl[159] br[159] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_162 
+ bl[160] br[160] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_163 
+ bl[161] br[161] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_164 
+ bl[162] br[162] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_165 
+ bl[163] br[163] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_166 
+ bl[164] br[164] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_167 
+ bl[165] br[165] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_168 
+ bl[166] br[166] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_169 
+ bl[167] br[167] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_170 
+ bl[168] br[168] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_171 
+ bl[169] br[169] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_172 
+ bl[170] br[170] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_173 
+ bl[171] br[171] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_174 
+ bl[172] br[172] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_175 
+ bl[173] br[173] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_176 
+ bl[174] br[174] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_177 
+ bl[175] br[175] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_178 
+ bl[176] br[176] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_179 
+ bl[177] br[177] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_180 
+ bl[178] br[178] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_181 
+ bl[179] br[179] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_182 
+ bl[180] br[180] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_183 
+ bl[181] br[181] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_184 
+ bl[182] br[182] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_185 
+ bl[183] br[183] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_186 
+ bl[184] br[184] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_187 
+ bl[185] br[185] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_188 
+ bl[186] br[186] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_189 
+ bl[187] br[187] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_190 
+ bl[188] br[188] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_191 
+ bl[189] br[189] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_192 
+ bl[190] br[190] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_193 
+ bl[191] br[191] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_194 
+ bl[192] br[192] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_195 
+ bl[193] br[193] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_196 
+ bl[194] br[194] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_197 
+ bl[195] br[195] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_198 
+ bl[196] br[196] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_199 
+ bl[197] br[197] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_200 
+ bl[198] br[198] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_201 
+ bl[199] br[199] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_202 
+ bl[200] br[200] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_203 
+ bl[201] br[201] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_204 
+ bl[202] br[202] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_205 
+ bl[203] br[203] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_206 
+ bl[204] br[204] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_207 
+ bl[205] br[205] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_208 
+ bl[206] br[206] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_209 
+ bl[207] br[207] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_210 
+ bl[208] br[208] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_211 
+ bl[209] br[209] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_212 
+ bl[210] br[210] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_213 
+ bl[211] br[211] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_214 
+ bl[212] br[212] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_215 
+ bl[213] br[213] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_216 
+ bl[214] br[214] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_217 
+ bl[215] br[215] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_218 
+ bl[216] br[216] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_219 
+ bl[217] br[217] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_220 
+ bl[218] br[218] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_221 
+ bl[219] br[219] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_222 
+ bl[220] br[220] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_223 
+ bl[221] br[221] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_224 
+ bl[222] br[222] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_225 
+ bl[223] br[223] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_226 
+ bl[224] br[224] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_227 
+ bl[225] br[225] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_228 
+ bl[226] br[226] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_229 
+ bl[227] br[227] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_230 
+ bl[228] br[228] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_231 
+ bl[229] br[229] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_232 
+ bl[230] br[230] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_233 
+ bl[231] br[231] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_234 
+ bl[232] br[232] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_235 
+ bl[233] br[233] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_236 
+ bl[234] br[234] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_237 
+ bl[235] br[235] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_238 
+ bl[236] br[236] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_239 
+ bl[237] br[237] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_240 
+ bl[238] br[238] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_241 
+ bl[239] br[239] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_242 
+ bl[240] br[240] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_243 
+ bl[241] br[241] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_244 
+ bl[242] br[242] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_245 
+ bl[243] br[243] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_246 
+ bl[244] br[244] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_247 
+ bl[245] br[245] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_248 
+ bl[246] br[246] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_249 
+ bl[247] br[247] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_250 
+ bl[248] br[248] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_251 
+ bl[249] br[249] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_252 
+ bl[250] br[250] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_253 
+ bl[251] br[251] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_254 
+ bl[252] br[252] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_255 
+ bl[253] br[253] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_256 
+ bl[254] br[254] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_257 
+ bl[255] br[255] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_258 
+ vdd vdd vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_259 
+ vdd vdd vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_0 
+ vdd vdd vss vdd vpb vnb wl[30] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_32_1 
+ rbl rbr vss vdd vpb vnb wl[30] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_32_2 
+ bl[0] br[0] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_3 
+ bl[1] br[1] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_4 
+ bl[2] br[2] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_5 
+ bl[3] br[3] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_6 
+ bl[4] br[4] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_7 
+ bl[5] br[5] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_8 
+ bl[6] br[6] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_9 
+ bl[7] br[7] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_10 
+ bl[8] br[8] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_11 
+ bl[9] br[9] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_12 
+ bl[10] br[10] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_13 
+ bl[11] br[11] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_14 
+ bl[12] br[12] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_15 
+ bl[13] br[13] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_16 
+ bl[14] br[14] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_17 
+ bl[15] br[15] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_18 
+ bl[16] br[16] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_19 
+ bl[17] br[17] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_20 
+ bl[18] br[18] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_21 
+ bl[19] br[19] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_22 
+ bl[20] br[20] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_23 
+ bl[21] br[21] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_24 
+ bl[22] br[22] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_25 
+ bl[23] br[23] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_26 
+ bl[24] br[24] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_27 
+ bl[25] br[25] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_28 
+ bl[26] br[26] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_29 
+ bl[27] br[27] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_30 
+ bl[28] br[28] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_31 
+ bl[29] br[29] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_32 
+ bl[30] br[30] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_33 
+ bl[31] br[31] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_34 
+ bl[32] br[32] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_35 
+ bl[33] br[33] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_36 
+ bl[34] br[34] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_37 
+ bl[35] br[35] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_38 
+ bl[36] br[36] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_39 
+ bl[37] br[37] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_40 
+ bl[38] br[38] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_41 
+ bl[39] br[39] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_42 
+ bl[40] br[40] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_43 
+ bl[41] br[41] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_44 
+ bl[42] br[42] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_45 
+ bl[43] br[43] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_46 
+ bl[44] br[44] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_47 
+ bl[45] br[45] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_48 
+ bl[46] br[46] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_49 
+ bl[47] br[47] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_50 
+ bl[48] br[48] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_51 
+ bl[49] br[49] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_52 
+ bl[50] br[50] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_53 
+ bl[51] br[51] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_54 
+ bl[52] br[52] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_55 
+ bl[53] br[53] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_56 
+ bl[54] br[54] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_57 
+ bl[55] br[55] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_58 
+ bl[56] br[56] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_59 
+ bl[57] br[57] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_60 
+ bl[58] br[58] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_61 
+ bl[59] br[59] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_62 
+ bl[60] br[60] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_63 
+ bl[61] br[61] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_64 
+ bl[62] br[62] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_65 
+ bl[63] br[63] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_66 
+ bl[64] br[64] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_67 
+ bl[65] br[65] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_68 
+ bl[66] br[66] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_69 
+ bl[67] br[67] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_70 
+ bl[68] br[68] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_71 
+ bl[69] br[69] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_72 
+ bl[70] br[70] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_73 
+ bl[71] br[71] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_74 
+ bl[72] br[72] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_75 
+ bl[73] br[73] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_76 
+ bl[74] br[74] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_77 
+ bl[75] br[75] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_78 
+ bl[76] br[76] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_79 
+ bl[77] br[77] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_80 
+ bl[78] br[78] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_81 
+ bl[79] br[79] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_82 
+ bl[80] br[80] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_83 
+ bl[81] br[81] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_84 
+ bl[82] br[82] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_85 
+ bl[83] br[83] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_86 
+ bl[84] br[84] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_87 
+ bl[85] br[85] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_88 
+ bl[86] br[86] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_89 
+ bl[87] br[87] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_90 
+ bl[88] br[88] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_91 
+ bl[89] br[89] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_92 
+ bl[90] br[90] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_93 
+ bl[91] br[91] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_94 
+ bl[92] br[92] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_95 
+ bl[93] br[93] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_96 
+ bl[94] br[94] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_97 
+ bl[95] br[95] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_98 
+ bl[96] br[96] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_99 
+ bl[97] br[97] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_100 
+ bl[98] br[98] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_101 
+ bl[99] br[99] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_102 
+ bl[100] br[100] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_103 
+ bl[101] br[101] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_104 
+ bl[102] br[102] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_105 
+ bl[103] br[103] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_106 
+ bl[104] br[104] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_107 
+ bl[105] br[105] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_108 
+ bl[106] br[106] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_109 
+ bl[107] br[107] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_110 
+ bl[108] br[108] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_111 
+ bl[109] br[109] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_112 
+ bl[110] br[110] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_113 
+ bl[111] br[111] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_114 
+ bl[112] br[112] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_115 
+ bl[113] br[113] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_116 
+ bl[114] br[114] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_117 
+ bl[115] br[115] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_118 
+ bl[116] br[116] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_119 
+ bl[117] br[117] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_120 
+ bl[118] br[118] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_121 
+ bl[119] br[119] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_122 
+ bl[120] br[120] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_123 
+ bl[121] br[121] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_124 
+ bl[122] br[122] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_125 
+ bl[123] br[123] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_126 
+ bl[124] br[124] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_127 
+ bl[125] br[125] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_128 
+ bl[126] br[126] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_129 
+ bl[127] br[127] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_130 
+ bl[128] br[128] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_131 
+ bl[129] br[129] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_132 
+ bl[130] br[130] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_133 
+ bl[131] br[131] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_134 
+ bl[132] br[132] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_135 
+ bl[133] br[133] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_136 
+ bl[134] br[134] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_137 
+ bl[135] br[135] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_138 
+ bl[136] br[136] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_139 
+ bl[137] br[137] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_140 
+ bl[138] br[138] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_141 
+ bl[139] br[139] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_142 
+ bl[140] br[140] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_143 
+ bl[141] br[141] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_144 
+ bl[142] br[142] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_145 
+ bl[143] br[143] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_146 
+ bl[144] br[144] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_147 
+ bl[145] br[145] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_148 
+ bl[146] br[146] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_149 
+ bl[147] br[147] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_150 
+ bl[148] br[148] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_151 
+ bl[149] br[149] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_152 
+ bl[150] br[150] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_153 
+ bl[151] br[151] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_154 
+ bl[152] br[152] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_155 
+ bl[153] br[153] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_156 
+ bl[154] br[154] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_157 
+ bl[155] br[155] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_158 
+ bl[156] br[156] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_159 
+ bl[157] br[157] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_160 
+ bl[158] br[158] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_161 
+ bl[159] br[159] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_162 
+ bl[160] br[160] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_163 
+ bl[161] br[161] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_164 
+ bl[162] br[162] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_165 
+ bl[163] br[163] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_166 
+ bl[164] br[164] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_167 
+ bl[165] br[165] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_168 
+ bl[166] br[166] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_169 
+ bl[167] br[167] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_170 
+ bl[168] br[168] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_171 
+ bl[169] br[169] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_172 
+ bl[170] br[170] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_173 
+ bl[171] br[171] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_174 
+ bl[172] br[172] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_175 
+ bl[173] br[173] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_176 
+ bl[174] br[174] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_177 
+ bl[175] br[175] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_178 
+ bl[176] br[176] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_179 
+ bl[177] br[177] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_180 
+ bl[178] br[178] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_181 
+ bl[179] br[179] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_182 
+ bl[180] br[180] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_183 
+ bl[181] br[181] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_184 
+ bl[182] br[182] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_185 
+ bl[183] br[183] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_186 
+ bl[184] br[184] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_187 
+ bl[185] br[185] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_188 
+ bl[186] br[186] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_189 
+ bl[187] br[187] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_190 
+ bl[188] br[188] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_191 
+ bl[189] br[189] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_192 
+ bl[190] br[190] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_193 
+ bl[191] br[191] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_194 
+ bl[192] br[192] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_195 
+ bl[193] br[193] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_196 
+ bl[194] br[194] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_197 
+ bl[195] br[195] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_198 
+ bl[196] br[196] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_199 
+ bl[197] br[197] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_200 
+ bl[198] br[198] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_201 
+ bl[199] br[199] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_202 
+ bl[200] br[200] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_203 
+ bl[201] br[201] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_204 
+ bl[202] br[202] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_205 
+ bl[203] br[203] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_206 
+ bl[204] br[204] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_207 
+ bl[205] br[205] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_208 
+ bl[206] br[206] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_209 
+ bl[207] br[207] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_210 
+ bl[208] br[208] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_211 
+ bl[209] br[209] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_212 
+ bl[210] br[210] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_213 
+ bl[211] br[211] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_214 
+ bl[212] br[212] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_215 
+ bl[213] br[213] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_216 
+ bl[214] br[214] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_217 
+ bl[215] br[215] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_218 
+ bl[216] br[216] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_219 
+ bl[217] br[217] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_220 
+ bl[218] br[218] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_221 
+ bl[219] br[219] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_222 
+ bl[220] br[220] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_223 
+ bl[221] br[221] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_224 
+ bl[222] br[222] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_225 
+ bl[223] br[223] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_226 
+ bl[224] br[224] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_227 
+ bl[225] br[225] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_228 
+ bl[226] br[226] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_229 
+ bl[227] br[227] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_230 
+ bl[228] br[228] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_231 
+ bl[229] br[229] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_232 
+ bl[230] br[230] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_233 
+ bl[231] br[231] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_234 
+ bl[232] br[232] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_235 
+ bl[233] br[233] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_236 
+ bl[234] br[234] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_237 
+ bl[235] br[235] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_238 
+ bl[236] br[236] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_239 
+ bl[237] br[237] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_240 
+ bl[238] br[238] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_241 
+ bl[239] br[239] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_242 
+ bl[240] br[240] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_243 
+ bl[241] br[241] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_244 
+ bl[242] br[242] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_245 
+ bl[243] br[243] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_246 
+ bl[244] br[244] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_247 
+ bl[245] br[245] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_248 
+ bl[246] br[246] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_249 
+ bl[247] br[247] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_250 
+ bl[248] br[248] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_251 
+ bl[249] br[249] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_252 
+ bl[250] br[250] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_253 
+ bl[251] br[251] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_254 
+ bl[252] br[252] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_255 
+ bl[253] br[253] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_256 
+ bl[254] br[254] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_257 
+ bl[255] br[255] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_258 
+ vdd vdd vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_259 
+ vdd vdd vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_0 
+ vdd vdd vss vdd vpb vnb wl[31] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_33_1 
+ rbl rbr vss vdd vpb vnb wl[31] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_33_2 
+ bl[0] br[0] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_3 
+ bl[1] br[1] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_4 
+ bl[2] br[2] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_5 
+ bl[3] br[3] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_6 
+ bl[4] br[4] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_7 
+ bl[5] br[5] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_8 
+ bl[6] br[6] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_9 
+ bl[7] br[7] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_10 
+ bl[8] br[8] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_11 
+ bl[9] br[9] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_12 
+ bl[10] br[10] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_13 
+ bl[11] br[11] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_14 
+ bl[12] br[12] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_15 
+ bl[13] br[13] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_16 
+ bl[14] br[14] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_17 
+ bl[15] br[15] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_18 
+ bl[16] br[16] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_19 
+ bl[17] br[17] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_20 
+ bl[18] br[18] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_21 
+ bl[19] br[19] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_22 
+ bl[20] br[20] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_23 
+ bl[21] br[21] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_24 
+ bl[22] br[22] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_25 
+ bl[23] br[23] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_26 
+ bl[24] br[24] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_27 
+ bl[25] br[25] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_28 
+ bl[26] br[26] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_29 
+ bl[27] br[27] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_30 
+ bl[28] br[28] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_31 
+ bl[29] br[29] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_32 
+ bl[30] br[30] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_33 
+ bl[31] br[31] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_34 
+ bl[32] br[32] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_35 
+ bl[33] br[33] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_36 
+ bl[34] br[34] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_37 
+ bl[35] br[35] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_38 
+ bl[36] br[36] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_39 
+ bl[37] br[37] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_40 
+ bl[38] br[38] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_41 
+ bl[39] br[39] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_42 
+ bl[40] br[40] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_43 
+ bl[41] br[41] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_44 
+ bl[42] br[42] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_45 
+ bl[43] br[43] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_46 
+ bl[44] br[44] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_47 
+ bl[45] br[45] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_48 
+ bl[46] br[46] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_49 
+ bl[47] br[47] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_50 
+ bl[48] br[48] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_51 
+ bl[49] br[49] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_52 
+ bl[50] br[50] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_53 
+ bl[51] br[51] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_54 
+ bl[52] br[52] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_55 
+ bl[53] br[53] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_56 
+ bl[54] br[54] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_57 
+ bl[55] br[55] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_58 
+ bl[56] br[56] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_59 
+ bl[57] br[57] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_60 
+ bl[58] br[58] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_61 
+ bl[59] br[59] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_62 
+ bl[60] br[60] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_63 
+ bl[61] br[61] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_64 
+ bl[62] br[62] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_65 
+ bl[63] br[63] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_66 
+ bl[64] br[64] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_67 
+ bl[65] br[65] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_68 
+ bl[66] br[66] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_69 
+ bl[67] br[67] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_70 
+ bl[68] br[68] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_71 
+ bl[69] br[69] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_72 
+ bl[70] br[70] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_73 
+ bl[71] br[71] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_74 
+ bl[72] br[72] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_75 
+ bl[73] br[73] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_76 
+ bl[74] br[74] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_77 
+ bl[75] br[75] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_78 
+ bl[76] br[76] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_79 
+ bl[77] br[77] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_80 
+ bl[78] br[78] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_81 
+ bl[79] br[79] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_82 
+ bl[80] br[80] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_83 
+ bl[81] br[81] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_84 
+ bl[82] br[82] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_85 
+ bl[83] br[83] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_86 
+ bl[84] br[84] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_87 
+ bl[85] br[85] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_88 
+ bl[86] br[86] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_89 
+ bl[87] br[87] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_90 
+ bl[88] br[88] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_91 
+ bl[89] br[89] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_92 
+ bl[90] br[90] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_93 
+ bl[91] br[91] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_94 
+ bl[92] br[92] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_95 
+ bl[93] br[93] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_96 
+ bl[94] br[94] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_97 
+ bl[95] br[95] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_98 
+ bl[96] br[96] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_99 
+ bl[97] br[97] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_100 
+ bl[98] br[98] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_101 
+ bl[99] br[99] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_102 
+ bl[100] br[100] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_103 
+ bl[101] br[101] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_104 
+ bl[102] br[102] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_105 
+ bl[103] br[103] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_106 
+ bl[104] br[104] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_107 
+ bl[105] br[105] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_108 
+ bl[106] br[106] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_109 
+ bl[107] br[107] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_110 
+ bl[108] br[108] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_111 
+ bl[109] br[109] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_112 
+ bl[110] br[110] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_113 
+ bl[111] br[111] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_114 
+ bl[112] br[112] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_115 
+ bl[113] br[113] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_116 
+ bl[114] br[114] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_117 
+ bl[115] br[115] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_118 
+ bl[116] br[116] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_119 
+ bl[117] br[117] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_120 
+ bl[118] br[118] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_121 
+ bl[119] br[119] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_122 
+ bl[120] br[120] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_123 
+ bl[121] br[121] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_124 
+ bl[122] br[122] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_125 
+ bl[123] br[123] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_126 
+ bl[124] br[124] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_127 
+ bl[125] br[125] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_128 
+ bl[126] br[126] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_129 
+ bl[127] br[127] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_130 
+ bl[128] br[128] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_131 
+ bl[129] br[129] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_132 
+ bl[130] br[130] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_133 
+ bl[131] br[131] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_134 
+ bl[132] br[132] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_135 
+ bl[133] br[133] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_136 
+ bl[134] br[134] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_137 
+ bl[135] br[135] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_138 
+ bl[136] br[136] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_139 
+ bl[137] br[137] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_140 
+ bl[138] br[138] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_141 
+ bl[139] br[139] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_142 
+ bl[140] br[140] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_143 
+ bl[141] br[141] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_144 
+ bl[142] br[142] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_145 
+ bl[143] br[143] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_146 
+ bl[144] br[144] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_147 
+ bl[145] br[145] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_148 
+ bl[146] br[146] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_149 
+ bl[147] br[147] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_150 
+ bl[148] br[148] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_151 
+ bl[149] br[149] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_152 
+ bl[150] br[150] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_153 
+ bl[151] br[151] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_154 
+ bl[152] br[152] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_155 
+ bl[153] br[153] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_156 
+ bl[154] br[154] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_157 
+ bl[155] br[155] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_158 
+ bl[156] br[156] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_159 
+ bl[157] br[157] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_160 
+ bl[158] br[158] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_161 
+ bl[159] br[159] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_162 
+ bl[160] br[160] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_163 
+ bl[161] br[161] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_164 
+ bl[162] br[162] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_165 
+ bl[163] br[163] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_166 
+ bl[164] br[164] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_167 
+ bl[165] br[165] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_168 
+ bl[166] br[166] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_169 
+ bl[167] br[167] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_170 
+ bl[168] br[168] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_171 
+ bl[169] br[169] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_172 
+ bl[170] br[170] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_173 
+ bl[171] br[171] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_174 
+ bl[172] br[172] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_175 
+ bl[173] br[173] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_176 
+ bl[174] br[174] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_177 
+ bl[175] br[175] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_178 
+ bl[176] br[176] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_179 
+ bl[177] br[177] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_180 
+ bl[178] br[178] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_181 
+ bl[179] br[179] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_182 
+ bl[180] br[180] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_183 
+ bl[181] br[181] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_184 
+ bl[182] br[182] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_185 
+ bl[183] br[183] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_186 
+ bl[184] br[184] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_187 
+ bl[185] br[185] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_188 
+ bl[186] br[186] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_189 
+ bl[187] br[187] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_190 
+ bl[188] br[188] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_191 
+ bl[189] br[189] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_192 
+ bl[190] br[190] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_193 
+ bl[191] br[191] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_194 
+ bl[192] br[192] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_195 
+ bl[193] br[193] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_196 
+ bl[194] br[194] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_197 
+ bl[195] br[195] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_198 
+ bl[196] br[196] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_199 
+ bl[197] br[197] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_200 
+ bl[198] br[198] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_201 
+ bl[199] br[199] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_202 
+ bl[200] br[200] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_203 
+ bl[201] br[201] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_204 
+ bl[202] br[202] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_205 
+ bl[203] br[203] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_206 
+ bl[204] br[204] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_207 
+ bl[205] br[205] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_208 
+ bl[206] br[206] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_209 
+ bl[207] br[207] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_210 
+ bl[208] br[208] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_211 
+ bl[209] br[209] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_212 
+ bl[210] br[210] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_213 
+ bl[211] br[211] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_214 
+ bl[212] br[212] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_215 
+ bl[213] br[213] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_216 
+ bl[214] br[214] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_217 
+ bl[215] br[215] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_218 
+ bl[216] br[216] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_219 
+ bl[217] br[217] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_220 
+ bl[218] br[218] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_221 
+ bl[219] br[219] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_222 
+ bl[220] br[220] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_223 
+ bl[221] br[221] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_224 
+ bl[222] br[222] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_225 
+ bl[223] br[223] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_226 
+ bl[224] br[224] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_227 
+ bl[225] br[225] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_228 
+ bl[226] br[226] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_229 
+ bl[227] br[227] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_230 
+ bl[228] br[228] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_231 
+ bl[229] br[229] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_232 
+ bl[230] br[230] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_233 
+ bl[231] br[231] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_234 
+ bl[232] br[232] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_235 
+ bl[233] br[233] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_236 
+ bl[234] br[234] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_237 
+ bl[235] br[235] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_238 
+ bl[236] br[236] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_239 
+ bl[237] br[237] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_240 
+ bl[238] br[238] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_241 
+ bl[239] br[239] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_242 
+ bl[240] br[240] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_243 
+ bl[241] br[241] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_244 
+ bl[242] br[242] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_245 
+ bl[243] br[243] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_246 
+ bl[244] br[244] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_247 
+ bl[245] br[245] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_248 
+ bl[246] br[246] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_249 
+ bl[247] br[247] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_250 
+ bl[248] br[248] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_251 
+ bl[249] br[249] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_252 
+ bl[250] br[250] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_253 
+ bl[251] br[251] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_254 
+ bl[252] br[252] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_255 
+ bl[253] br[253] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_256 
+ bl[254] br[254] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_257 
+ bl[255] br[255] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_258 
+ vdd vdd vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_259 
+ vdd vdd vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_0 
+ vdd vdd vss vdd vpb vnb wl[32] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_34_1 
+ rbl rbr vss vdd vpb vnb wl[32] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_34_2 
+ bl[0] br[0] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_3 
+ bl[1] br[1] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_4 
+ bl[2] br[2] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_5 
+ bl[3] br[3] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_6 
+ bl[4] br[4] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_7 
+ bl[5] br[5] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_8 
+ bl[6] br[6] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_9 
+ bl[7] br[7] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_10 
+ bl[8] br[8] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_11 
+ bl[9] br[9] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_12 
+ bl[10] br[10] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_13 
+ bl[11] br[11] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_14 
+ bl[12] br[12] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_15 
+ bl[13] br[13] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_16 
+ bl[14] br[14] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_17 
+ bl[15] br[15] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_18 
+ bl[16] br[16] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_19 
+ bl[17] br[17] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_20 
+ bl[18] br[18] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_21 
+ bl[19] br[19] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_22 
+ bl[20] br[20] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_23 
+ bl[21] br[21] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_24 
+ bl[22] br[22] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_25 
+ bl[23] br[23] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_26 
+ bl[24] br[24] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_27 
+ bl[25] br[25] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_28 
+ bl[26] br[26] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_29 
+ bl[27] br[27] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_30 
+ bl[28] br[28] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_31 
+ bl[29] br[29] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_32 
+ bl[30] br[30] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_33 
+ bl[31] br[31] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_34 
+ bl[32] br[32] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_35 
+ bl[33] br[33] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_36 
+ bl[34] br[34] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_37 
+ bl[35] br[35] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_38 
+ bl[36] br[36] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_39 
+ bl[37] br[37] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_40 
+ bl[38] br[38] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_41 
+ bl[39] br[39] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_42 
+ bl[40] br[40] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_43 
+ bl[41] br[41] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_44 
+ bl[42] br[42] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_45 
+ bl[43] br[43] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_46 
+ bl[44] br[44] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_47 
+ bl[45] br[45] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_48 
+ bl[46] br[46] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_49 
+ bl[47] br[47] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_50 
+ bl[48] br[48] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_51 
+ bl[49] br[49] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_52 
+ bl[50] br[50] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_53 
+ bl[51] br[51] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_54 
+ bl[52] br[52] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_55 
+ bl[53] br[53] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_56 
+ bl[54] br[54] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_57 
+ bl[55] br[55] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_58 
+ bl[56] br[56] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_59 
+ bl[57] br[57] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_60 
+ bl[58] br[58] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_61 
+ bl[59] br[59] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_62 
+ bl[60] br[60] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_63 
+ bl[61] br[61] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_64 
+ bl[62] br[62] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_65 
+ bl[63] br[63] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_66 
+ bl[64] br[64] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_67 
+ bl[65] br[65] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_68 
+ bl[66] br[66] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_69 
+ bl[67] br[67] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_70 
+ bl[68] br[68] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_71 
+ bl[69] br[69] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_72 
+ bl[70] br[70] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_73 
+ bl[71] br[71] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_74 
+ bl[72] br[72] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_75 
+ bl[73] br[73] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_76 
+ bl[74] br[74] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_77 
+ bl[75] br[75] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_78 
+ bl[76] br[76] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_79 
+ bl[77] br[77] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_80 
+ bl[78] br[78] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_81 
+ bl[79] br[79] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_82 
+ bl[80] br[80] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_83 
+ bl[81] br[81] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_84 
+ bl[82] br[82] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_85 
+ bl[83] br[83] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_86 
+ bl[84] br[84] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_87 
+ bl[85] br[85] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_88 
+ bl[86] br[86] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_89 
+ bl[87] br[87] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_90 
+ bl[88] br[88] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_91 
+ bl[89] br[89] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_92 
+ bl[90] br[90] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_93 
+ bl[91] br[91] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_94 
+ bl[92] br[92] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_95 
+ bl[93] br[93] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_96 
+ bl[94] br[94] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_97 
+ bl[95] br[95] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_98 
+ bl[96] br[96] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_99 
+ bl[97] br[97] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_100 
+ bl[98] br[98] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_101 
+ bl[99] br[99] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_102 
+ bl[100] br[100] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_103 
+ bl[101] br[101] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_104 
+ bl[102] br[102] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_105 
+ bl[103] br[103] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_106 
+ bl[104] br[104] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_107 
+ bl[105] br[105] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_108 
+ bl[106] br[106] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_109 
+ bl[107] br[107] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_110 
+ bl[108] br[108] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_111 
+ bl[109] br[109] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_112 
+ bl[110] br[110] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_113 
+ bl[111] br[111] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_114 
+ bl[112] br[112] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_115 
+ bl[113] br[113] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_116 
+ bl[114] br[114] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_117 
+ bl[115] br[115] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_118 
+ bl[116] br[116] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_119 
+ bl[117] br[117] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_120 
+ bl[118] br[118] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_121 
+ bl[119] br[119] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_122 
+ bl[120] br[120] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_123 
+ bl[121] br[121] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_124 
+ bl[122] br[122] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_125 
+ bl[123] br[123] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_126 
+ bl[124] br[124] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_127 
+ bl[125] br[125] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_128 
+ bl[126] br[126] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_129 
+ bl[127] br[127] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_130 
+ bl[128] br[128] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_131 
+ bl[129] br[129] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_132 
+ bl[130] br[130] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_133 
+ bl[131] br[131] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_134 
+ bl[132] br[132] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_135 
+ bl[133] br[133] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_136 
+ bl[134] br[134] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_137 
+ bl[135] br[135] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_138 
+ bl[136] br[136] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_139 
+ bl[137] br[137] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_140 
+ bl[138] br[138] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_141 
+ bl[139] br[139] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_142 
+ bl[140] br[140] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_143 
+ bl[141] br[141] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_144 
+ bl[142] br[142] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_145 
+ bl[143] br[143] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_146 
+ bl[144] br[144] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_147 
+ bl[145] br[145] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_148 
+ bl[146] br[146] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_149 
+ bl[147] br[147] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_150 
+ bl[148] br[148] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_151 
+ bl[149] br[149] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_152 
+ bl[150] br[150] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_153 
+ bl[151] br[151] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_154 
+ bl[152] br[152] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_155 
+ bl[153] br[153] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_156 
+ bl[154] br[154] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_157 
+ bl[155] br[155] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_158 
+ bl[156] br[156] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_159 
+ bl[157] br[157] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_160 
+ bl[158] br[158] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_161 
+ bl[159] br[159] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_162 
+ bl[160] br[160] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_163 
+ bl[161] br[161] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_164 
+ bl[162] br[162] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_165 
+ bl[163] br[163] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_166 
+ bl[164] br[164] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_167 
+ bl[165] br[165] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_168 
+ bl[166] br[166] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_169 
+ bl[167] br[167] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_170 
+ bl[168] br[168] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_171 
+ bl[169] br[169] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_172 
+ bl[170] br[170] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_173 
+ bl[171] br[171] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_174 
+ bl[172] br[172] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_175 
+ bl[173] br[173] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_176 
+ bl[174] br[174] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_177 
+ bl[175] br[175] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_178 
+ bl[176] br[176] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_179 
+ bl[177] br[177] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_180 
+ bl[178] br[178] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_181 
+ bl[179] br[179] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_182 
+ bl[180] br[180] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_183 
+ bl[181] br[181] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_184 
+ bl[182] br[182] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_185 
+ bl[183] br[183] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_186 
+ bl[184] br[184] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_187 
+ bl[185] br[185] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_188 
+ bl[186] br[186] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_189 
+ bl[187] br[187] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_190 
+ bl[188] br[188] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_191 
+ bl[189] br[189] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_192 
+ bl[190] br[190] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_193 
+ bl[191] br[191] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_194 
+ bl[192] br[192] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_195 
+ bl[193] br[193] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_196 
+ bl[194] br[194] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_197 
+ bl[195] br[195] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_198 
+ bl[196] br[196] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_199 
+ bl[197] br[197] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_200 
+ bl[198] br[198] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_201 
+ bl[199] br[199] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_202 
+ bl[200] br[200] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_203 
+ bl[201] br[201] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_204 
+ bl[202] br[202] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_205 
+ bl[203] br[203] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_206 
+ bl[204] br[204] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_207 
+ bl[205] br[205] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_208 
+ bl[206] br[206] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_209 
+ bl[207] br[207] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_210 
+ bl[208] br[208] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_211 
+ bl[209] br[209] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_212 
+ bl[210] br[210] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_213 
+ bl[211] br[211] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_214 
+ bl[212] br[212] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_215 
+ bl[213] br[213] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_216 
+ bl[214] br[214] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_217 
+ bl[215] br[215] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_218 
+ bl[216] br[216] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_219 
+ bl[217] br[217] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_220 
+ bl[218] br[218] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_221 
+ bl[219] br[219] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_222 
+ bl[220] br[220] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_223 
+ bl[221] br[221] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_224 
+ bl[222] br[222] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_225 
+ bl[223] br[223] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_226 
+ bl[224] br[224] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_227 
+ bl[225] br[225] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_228 
+ bl[226] br[226] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_229 
+ bl[227] br[227] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_230 
+ bl[228] br[228] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_231 
+ bl[229] br[229] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_232 
+ bl[230] br[230] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_233 
+ bl[231] br[231] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_234 
+ bl[232] br[232] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_235 
+ bl[233] br[233] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_236 
+ bl[234] br[234] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_237 
+ bl[235] br[235] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_238 
+ bl[236] br[236] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_239 
+ bl[237] br[237] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_240 
+ bl[238] br[238] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_241 
+ bl[239] br[239] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_242 
+ bl[240] br[240] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_243 
+ bl[241] br[241] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_244 
+ bl[242] br[242] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_245 
+ bl[243] br[243] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_246 
+ bl[244] br[244] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_247 
+ bl[245] br[245] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_248 
+ bl[246] br[246] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_249 
+ bl[247] br[247] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_250 
+ bl[248] br[248] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_251 
+ bl[249] br[249] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_252 
+ bl[250] br[250] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_253 
+ bl[251] br[251] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_254 
+ bl[252] br[252] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_255 
+ bl[253] br[253] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_256 
+ bl[254] br[254] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_257 
+ bl[255] br[255] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_258 
+ vdd vdd vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_259 
+ vdd vdd vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_0 
+ vdd vdd vss vdd vpb vnb wl[33] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_35_1 
+ rbl rbr vss vdd vpb vnb wl[33] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_35_2 
+ bl[0] br[0] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_3 
+ bl[1] br[1] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_4 
+ bl[2] br[2] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_5 
+ bl[3] br[3] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_6 
+ bl[4] br[4] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_7 
+ bl[5] br[5] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_8 
+ bl[6] br[6] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_9 
+ bl[7] br[7] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_10 
+ bl[8] br[8] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_11 
+ bl[9] br[9] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_12 
+ bl[10] br[10] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_13 
+ bl[11] br[11] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_14 
+ bl[12] br[12] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_15 
+ bl[13] br[13] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_16 
+ bl[14] br[14] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_17 
+ bl[15] br[15] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_18 
+ bl[16] br[16] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_19 
+ bl[17] br[17] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_20 
+ bl[18] br[18] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_21 
+ bl[19] br[19] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_22 
+ bl[20] br[20] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_23 
+ bl[21] br[21] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_24 
+ bl[22] br[22] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_25 
+ bl[23] br[23] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_26 
+ bl[24] br[24] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_27 
+ bl[25] br[25] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_28 
+ bl[26] br[26] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_29 
+ bl[27] br[27] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_30 
+ bl[28] br[28] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_31 
+ bl[29] br[29] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_32 
+ bl[30] br[30] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_33 
+ bl[31] br[31] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_34 
+ bl[32] br[32] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_35 
+ bl[33] br[33] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_36 
+ bl[34] br[34] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_37 
+ bl[35] br[35] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_38 
+ bl[36] br[36] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_39 
+ bl[37] br[37] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_40 
+ bl[38] br[38] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_41 
+ bl[39] br[39] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_42 
+ bl[40] br[40] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_43 
+ bl[41] br[41] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_44 
+ bl[42] br[42] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_45 
+ bl[43] br[43] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_46 
+ bl[44] br[44] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_47 
+ bl[45] br[45] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_48 
+ bl[46] br[46] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_49 
+ bl[47] br[47] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_50 
+ bl[48] br[48] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_51 
+ bl[49] br[49] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_52 
+ bl[50] br[50] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_53 
+ bl[51] br[51] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_54 
+ bl[52] br[52] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_55 
+ bl[53] br[53] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_56 
+ bl[54] br[54] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_57 
+ bl[55] br[55] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_58 
+ bl[56] br[56] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_59 
+ bl[57] br[57] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_60 
+ bl[58] br[58] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_61 
+ bl[59] br[59] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_62 
+ bl[60] br[60] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_63 
+ bl[61] br[61] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_64 
+ bl[62] br[62] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_65 
+ bl[63] br[63] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_66 
+ bl[64] br[64] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_67 
+ bl[65] br[65] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_68 
+ bl[66] br[66] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_69 
+ bl[67] br[67] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_70 
+ bl[68] br[68] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_71 
+ bl[69] br[69] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_72 
+ bl[70] br[70] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_73 
+ bl[71] br[71] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_74 
+ bl[72] br[72] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_75 
+ bl[73] br[73] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_76 
+ bl[74] br[74] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_77 
+ bl[75] br[75] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_78 
+ bl[76] br[76] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_79 
+ bl[77] br[77] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_80 
+ bl[78] br[78] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_81 
+ bl[79] br[79] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_82 
+ bl[80] br[80] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_83 
+ bl[81] br[81] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_84 
+ bl[82] br[82] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_85 
+ bl[83] br[83] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_86 
+ bl[84] br[84] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_87 
+ bl[85] br[85] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_88 
+ bl[86] br[86] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_89 
+ bl[87] br[87] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_90 
+ bl[88] br[88] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_91 
+ bl[89] br[89] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_92 
+ bl[90] br[90] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_93 
+ bl[91] br[91] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_94 
+ bl[92] br[92] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_95 
+ bl[93] br[93] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_96 
+ bl[94] br[94] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_97 
+ bl[95] br[95] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_98 
+ bl[96] br[96] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_99 
+ bl[97] br[97] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_100 
+ bl[98] br[98] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_101 
+ bl[99] br[99] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_102 
+ bl[100] br[100] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_103 
+ bl[101] br[101] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_104 
+ bl[102] br[102] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_105 
+ bl[103] br[103] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_106 
+ bl[104] br[104] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_107 
+ bl[105] br[105] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_108 
+ bl[106] br[106] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_109 
+ bl[107] br[107] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_110 
+ bl[108] br[108] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_111 
+ bl[109] br[109] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_112 
+ bl[110] br[110] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_113 
+ bl[111] br[111] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_114 
+ bl[112] br[112] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_115 
+ bl[113] br[113] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_116 
+ bl[114] br[114] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_117 
+ bl[115] br[115] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_118 
+ bl[116] br[116] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_119 
+ bl[117] br[117] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_120 
+ bl[118] br[118] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_121 
+ bl[119] br[119] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_122 
+ bl[120] br[120] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_123 
+ bl[121] br[121] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_124 
+ bl[122] br[122] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_125 
+ bl[123] br[123] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_126 
+ bl[124] br[124] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_127 
+ bl[125] br[125] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_128 
+ bl[126] br[126] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_129 
+ bl[127] br[127] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_130 
+ bl[128] br[128] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_131 
+ bl[129] br[129] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_132 
+ bl[130] br[130] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_133 
+ bl[131] br[131] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_134 
+ bl[132] br[132] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_135 
+ bl[133] br[133] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_136 
+ bl[134] br[134] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_137 
+ bl[135] br[135] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_138 
+ bl[136] br[136] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_139 
+ bl[137] br[137] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_140 
+ bl[138] br[138] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_141 
+ bl[139] br[139] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_142 
+ bl[140] br[140] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_143 
+ bl[141] br[141] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_144 
+ bl[142] br[142] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_145 
+ bl[143] br[143] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_146 
+ bl[144] br[144] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_147 
+ bl[145] br[145] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_148 
+ bl[146] br[146] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_149 
+ bl[147] br[147] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_150 
+ bl[148] br[148] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_151 
+ bl[149] br[149] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_152 
+ bl[150] br[150] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_153 
+ bl[151] br[151] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_154 
+ bl[152] br[152] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_155 
+ bl[153] br[153] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_156 
+ bl[154] br[154] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_157 
+ bl[155] br[155] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_158 
+ bl[156] br[156] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_159 
+ bl[157] br[157] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_160 
+ bl[158] br[158] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_161 
+ bl[159] br[159] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_162 
+ bl[160] br[160] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_163 
+ bl[161] br[161] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_164 
+ bl[162] br[162] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_165 
+ bl[163] br[163] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_166 
+ bl[164] br[164] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_167 
+ bl[165] br[165] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_168 
+ bl[166] br[166] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_169 
+ bl[167] br[167] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_170 
+ bl[168] br[168] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_171 
+ bl[169] br[169] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_172 
+ bl[170] br[170] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_173 
+ bl[171] br[171] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_174 
+ bl[172] br[172] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_175 
+ bl[173] br[173] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_176 
+ bl[174] br[174] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_177 
+ bl[175] br[175] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_178 
+ bl[176] br[176] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_179 
+ bl[177] br[177] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_180 
+ bl[178] br[178] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_181 
+ bl[179] br[179] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_182 
+ bl[180] br[180] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_183 
+ bl[181] br[181] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_184 
+ bl[182] br[182] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_185 
+ bl[183] br[183] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_186 
+ bl[184] br[184] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_187 
+ bl[185] br[185] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_188 
+ bl[186] br[186] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_189 
+ bl[187] br[187] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_190 
+ bl[188] br[188] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_191 
+ bl[189] br[189] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_192 
+ bl[190] br[190] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_193 
+ bl[191] br[191] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_194 
+ bl[192] br[192] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_195 
+ bl[193] br[193] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_196 
+ bl[194] br[194] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_197 
+ bl[195] br[195] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_198 
+ bl[196] br[196] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_199 
+ bl[197] br[197] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_200 
+ bl[198] br[198] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_201 
+ bl[199] br[199] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_202 
+ bl[200] br[200] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_203 
+ bl[201] br[201] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_204 
+ bl[202] br[202] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_205 
+ bl[203] br[203] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_206 
+ bl[204] br[204] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_207 
+ bl[205] br[205] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_208 
+ bl[206] br[206] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_209 
+ bl[207] br[207] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_210 
+ bl[208] br[208] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_211 
+ bl[209] br[209] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_212 
+ bl[210] br[210] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_213 
+ bl[211] br[211] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_214 
+ bl[212] br[212] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_215 
+ bl[213] br[213] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_216 
+ bl[214] br[214] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_217 
+ bl[215] br[215] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_218 
+ bl[216] br[216] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_219 
+ bl[217] br[217] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_220 
+ bl[218] br[218] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_221 
+ bl[219] br[219] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_222 
+ bl[220] br[220] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_223 
+ bl[221] br[221] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_224 
+ bl[222] br[222] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_225 
+ bl[223] br[223] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_226 
+ bl[224] br[224] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_227 
+ bl[225] br[225] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_228 
+ bl[226] br[226] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_229 
+ bl[227] br[227] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_230 
+ bl[228] br[228] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_231 
+ bl[229] br[229] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_232 
+ bl[230] br[230] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_233 
+ bl[231] br[231] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_234 
+ bl[232] br[232] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_235 
+ bl[233] br[233] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_236 
+ bl[234] br[234] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_237 
+ bl[235] br[235] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_238 
+ bl[236] br[236] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_239 
+ bl[237] br[237] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_240 
+ bl[238] br[238] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_241 
+ bl[239] br[239] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_242 
+ bl[240] br[240] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_243 
+ bl[241] br[241] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_244 
+ bl[242] br[242] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_245 
+ bl[243] br[243] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_246 
+ bl[244] br[244] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_247 
+ bl[245] br[245] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_248 
+ bl[246] br[246] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_249 
+ bl[247] br[247] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_250 
+ bl[248] br[248] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_251 
+ bl[249] br[249] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_252 
+ bl[250] br[250] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_253 
+ bl[251] br[251] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_254 
+ bl[252] br[252] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_255 
+ bl[253] br[253] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_256 
+ bl[254] br[254] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_257 
+ bl[255] br[255] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_258 
+ vdd vdd vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_259 
+ vdd vdd vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_0 
+ vdd vdd vss vdd vpb vnb wl[34] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_36_1 
+ rbl rbr vss vdd vpb vnb wl[34] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_36_2 
+ bl[0] br[0] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_3 
+ bl[1] br[1] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_4 
+ bl[2] br[2] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_5 
+ bl[3] br[3] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_6 
+ bl[4] br[4] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_7 
+ bl[5] br[5] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_8 
+ bl[6] br[6] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_9 
+ bl[7] br[7] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_10 
+ bl[8] br[8] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_11 
+ bl[9] br[9] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_12 
+ bl[10] br[10] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_13 
+ bl[11] br[11] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_14 
+ bl[12] br[12] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_15 
+ bl[13] br[13] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_16 
+ bl[14] br[14] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_17 
+ bl[15] br[15] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_18 
+ bl[16] br[16] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_19 
+ bl[17] br[17] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_20 
+ bl[18] br[18] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_21 
+ bl[19] br[19] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_22 
+ bl[20] br[20] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_23 
+ bl[21] br[21] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_24 
+ bl[22] br[22] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_25 
+ bl[23] br[23] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_26 
+ bl[24] br[24] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_27 
+ bl[25] br[25] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_28 
+ bl[26] br[26] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_29 
+ bl[27] br[27] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_30 
+ bl[28] br[28] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_31 
+ bl[29] br[29] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_32 
+ bl[30] br[30] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_33 
+ bl[31] br[31] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_34 
+ bl[32] br[32] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_35 
+ bl[33] br[33] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_36 
+ bl[34] br[34] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_37 
+ bl[35] br[35] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_38 
+ bl[36] br[36] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_39 
+ bl[37] br[37] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_40 
+ bl[38] br[38] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_41 
+ bl[39] br[39] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_42 
+ bl[40] br[40] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_43 
+ bl[41] br[41] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_44 
+ bl[42] br[42] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_45 
+ bl[43] br[43] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_46 
+ bl[44] br[44] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_47 
+ bl[45] br[45] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_48 
+ bl[46] br[46] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_49 
+ bl[47] br[47] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_50 
+ bl[48] br[48] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_51 
+ bl[49] br[49] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_52 
+ bl[50] br[50] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_53 
+ bl[51] br[51] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_54 
+ bl[52] br[52] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_55 
+ bl[53] br[53] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_56 
+ bl[54] br[54] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_57 
+ bl[55] br[55] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_58 
+ bl[56] br[56] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_59 
+ bl[57] br[57] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_60 
+ bl[58] br[58] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_61 
+ bl[59] br[59] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_62 
+ bl[60] br[60] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_63 
+ bl[61] br[61] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_64 
+ bl[62] br[62] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_65 
+ bl[63] br[63] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_66 
+ bl[64] br[64] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_67 
+ bl[65] br[65] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_68 
+ bl[66] br[66] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_69 
+ bl[67] br[67] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_70 
+ bl[68] br[68] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_71 
+ bl[69] br[69] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_72 
+ bl[70] br[70] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_73 
+ bl[71] br[71] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_74 
+ bl[72] br[72] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_75 
+ bl[73] br[73] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_76 
+ bl[74] br[74] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_77 
+ bl[75] br[75] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_78 
+ bl[76] br[76] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_79 
+ bl[77] br[77] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_80 
+ bl[78] br[78] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_81 
+ bl[79] br[79] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_82 
+ bl[80] br[80] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_83 
+ bl[81] br[81] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_84 
+ bl[82] br[82] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_85 
+ bl[83] br[83] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_86 
+ bl[84] br[84] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_87 
+ bl[85] br[85] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_88 
+ bl[86] br[86] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_89 
+ bl[87] br[87] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_90 
+ bl[88] br[88] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_91 
+ bl[89] br[89] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_92 
+ bl[90] br[90] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_93 
+ bl[91] br[91] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_94 
+ bl[92] br[92] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_95 
+ bl[93] br[93] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_96 
+ bl[94] br[94] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_97 
+ bl[95] br[95] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_98 
+ bl[96] br[96] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_99 
+ bl[97] br[97] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_100 
+ bl[98] br[98] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_101 
+ bl[99] br[99] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_102 
+ bl[100] br[100] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_103 
+ bl[101] br[101] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_104 
+ bl[102] br[102] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_105 
+ bl[103] br[103] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_106 
+ bl[104] br[104] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_107 
+ bl[105] br[105] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_108 
+ bl[106] br[106] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_109 
+ bl[107] br[107] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_110 
+ bl[108] br[108] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_111 
+ bl[109] br[109] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_112 
+ bl[110] br[110] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_113 
+ bl[111] br[111] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_114 
+ bl[112] br[112] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_115 
+ bl[113] br[113] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_116 
+ bl[114] br[114] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_117 
+ bl[115] br[115] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_118 
+ bl[116] br[116] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_119 
+ bl[117] br[117] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_120 
+ bl[118] br[118] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_121 
+ bl[119] br[119] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_122 
+ bl[120] br[120] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_123 
+ bl[121] br[121] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_124 
+ bl[122] br[122] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_125 
+ bl[123] br[123] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_126 
+ bl[124] br[124] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_127 
+ bl[125] br[125] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_128 
+ bl[126] br[126] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_129 
+ bl[127] br[127] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_130 
+ bl[128] br[128] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_131 
+ bl[129] br[129] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_132 
+ bl[130] br[130] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_133 
+ bl[131] br[131] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_134 
+ bl[132] br[132] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_135 
+ bl[133] br[133] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_136 
+ bl[134] br[134] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_137 
+ bl[135] br[135] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_138 
+ bl[136] br[136] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_139 
+ bl[137] br[137] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_140 
+ bl[138] br[138] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_141 
+ bl[139] br[139] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_142 
+ bl[140] br[140] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_143 
+ bl[141] br[141] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_144 
+ bl[142] br[142] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_145 
+ bl[143] br[143] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_146 
+ bl[144] br[144] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_147 
+ bl[145] br[145] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_148 
+ bl[146] br[146] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_149 
+ bl[147] br[147] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_150 
+ bl[148] br[148] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_151 
+ bl[149] br[149] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_152 
+ bl[150] br[150] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_153 
+ bl[151] br[151] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_154 
+ bl[152] br[152] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_155 
+ bl[153] br[153] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_156 
+ bl[154] br[154] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_157 
+ bl[155] br[155] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_158 
+ bl[156] br[156] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_159 
+ bl[157] br[157] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_160 
+ bl[158] br[158] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_161 
+ bl[159] br[159] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_162 
+ bl[160] br[160] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_163 
+ bl[161] br[161] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_164 
+ bl[162] br[162] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_165 
+ bl[163] br[163] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_166 
+ bl[164] br[164] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_167 
+ bl[165] br[165] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_168 
+ bl[166] br[166] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_169 
+ bl[167] br[167] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_170 
+ bl[168] br[168] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_171 
+ bl[169] br[169] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_172 
+ bl[170] br[170] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_173 
+ bl[171] br[171] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_174 
+ bl[172] br[172] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_175 
+ bl[173] br[173] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_176 
+ bl[174] br[174] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_177 
+ bl[175] br[175] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_178 
+ bl[176] br[176] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_179 
+ bl[177] br[177] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_180 
+ bl[178] br[178] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_181 
+ bl[179] br[179] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_182 
+ bl[180] br[180] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_183 
+ bl[181] br[181] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_184 
+ bl[182] br[182] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_185 
+ bl[183] br[183] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_186 
+ bl[184] br[184] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_187 
+ bl[185] br[185] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_188 
+ bl[186] br[186] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_189 
+ bl[187] br[187] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_190 
+ bl[188] br[188] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_191 
+ bl[189] br[189] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_192 
+ bl[190] br[190] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_193 
+ bl[191] br[191] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_194 
+ bl[192] br[192] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_195 
+ bl[193] br[193] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_196 
+ bl[194] br[194] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_197 
+ bl[195] br[195] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_198 
+ bl[196] br[196] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_199 
+ bl[197] br[197] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_200 
+ bl[198] br[198] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_201 
+ bl[199] br[199] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_202 
+ bl[200] br[200] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_203 
+ bl[201] br[201] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_204 
+ bl[202] br[202] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_205 
+ bl[203] br[203] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_206 
+ bl[204] br[204] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_207 
+ bl[205] br[205] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_208 
+ bl[206] br[206] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_209 
+ bl[207] br[207] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_210 
+ bl[208] br[208] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_211 
+ bl[209] br[209] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_212 
+ bl[210] br[210] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_213 
+ bl[211] br[211] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_214 
+ bl[212] br[212] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_215 
+ bl[213] br[213] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_216 
+ bl[214] br[214] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_217 
+ bl[215] br[215] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_218 
+ bl[216] br[216] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_219 
+ bl[217] br[217] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_220 
+ bl[218] br[218] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_221 
+ bl[219] br[219] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_222 
+ bl[220] br[220] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_223 
+ bl[221] br[221] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_224 
+ bl[222] br[222] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_225 
+ bl[223] br[223] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_226 
+ bl[224] br[224] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_227 
+ bl[225] br[225] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_228 
+ bl[226] br[226] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_229 
+ bl[227] br[227] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_230 
+ bl[228] br[228] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_231 
+ bl[229] br[229] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_232 
+ bl[230] br[230] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_233 
+ bl[231] br[231] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_234 
+ bl[232] br[232] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_235 
+ bl[233] br[233] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_236 
+ bl[234] br[234] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_237 
+ bl[235] br[235] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_238 
+ bl[236] br[236] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_239 
+ bl[237] br[237] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_240 
+ bl[238] br[238] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_241 
+ bl[239] br[239] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_242 
+ bl[240] br[240] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_243 
+ bl[241] br[241] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_244 
+ bl[242] br[242] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_245 
+ bl[243] br[243] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_246 
+ bl[244] br[244] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_247 
+ bl[245] br[245] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_248 
+ bl[246] br[246] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_249 
+ bl[247] br[247] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_250 
+ bl[248] br[248] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_251 
+ bl[249] br[249] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_252 
+ bl[250] br[250] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_253 
+ bl[251] br[251] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_254 
+ bl[252] br[252] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_255 
+ bl[253] br[253] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_256 
+ bl[254] br[254] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_257 
+ bl[255] br[255] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_258 
+ vdd vdd vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_259 
+ vdd vdd vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_0 
+ vdd vdd vss vdd vpb vnb wl[35] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_37_1 
+ rbl rbr vss vdd vpb vnb wl[35] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_37_2 
+ bl[0] br[0] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_3 
+ bl[1] br[1] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_4 
+ bl[2] br[2] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_5 
+ bl[3] br[3] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_6 
+ bl[4] br[4] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_7 
+ bl[5] br[5] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_8 
+ bl[6] br[6] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_9 
+ bl[7] br[7] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_10 
+ bl[8] br[8] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_11 
+ bl[9] br[9] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_12 
+ bl[10] br[10] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_13 
+ bl[11] br[11] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_14 
+ bl[12] br[12] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_15 
+ bl[13] br[13] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_16 
+ bl[14] br[14] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_17 
+ bl[15] br[15] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_18 
+ bl[16] br[16] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_19 
+ bl[17] br[17] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_20 
+ bl[18] br[18] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_21 
+ bl[19] br[19] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_22 
+ bl[20] br[20] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_23 
+ bl[21] br[21] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_24 
+ bl[22] br[22] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_25 
+ bl[23] br[23] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_26 
+ bl[24] br[24] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_27 
+ bl[25] br[25] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_28 
+ bl[26] br[26] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_29 
+ bl[27] br[27] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_30 
+ bl[28] br[28] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_31 
+ bl[29] br[29] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_32 
+ bl[30] br[30] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_33 
+ bl[31] br[31] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_34 
+ bl[32] br[32] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_35 
+ bl[33] br[33] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_36 
+ bl[34] br[34] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_37 
+ bl[35] br[35] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_38 
+ bl[36] br[36] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_39 
+ bl[37] br[37] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_40 
+ bl[38] br[38] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_41 
+ bl[39] br[39] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_42 
+ bl[40] br[40] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_43 
+ bl[41] br[41] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_44 
+ bl[42] br[42] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_45 
+ bl[43] br[43] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_46 
+ bl[44] br[44] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_47 
+ bl[45] br[45] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_48 
+ bl[46] br[46] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_49 
+ bl[47] br[47] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_50 
+ bl[48] br[48] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_51 
+ bl[49] br[49] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_52 
+ bl[50] br[50] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_53 
+ bl[51] br[51] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_54 
+ bl[52] br[52] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_55 
+ bl[53] br[53] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_56 
+ bl[54] br[54] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_57 
+ bl[55] br[55] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_58 
+ bl[56] br[56] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_59 
+ bl[57] br[57] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_60 
+ bl[58] br[58] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_61 
+ bl[59] br[59] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_62 
+ bl[60] br[60] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_63 
+ bl[61] br[61] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_64 
+ bl[62] br[62] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_65 
+ bl[63] br[63] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_66 
+ bl[64] br[64] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_67 
+ bl[65] br[65] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_68 
+ bl[66] br[66] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_69 
+ bl[67] br[67] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_70 
+ bl[68] br[68] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_71 
+ bl[69] br[69] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_72 
+ bl[70] br[70] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_73 
+ bl[71] br[71] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_74 
+ bl[72] br[72] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_75 
+ bl[73] br[73] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_76 
+ bl[74] br[74] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_77 
+ bl[75] br[75] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_78 
+ bl[76] br[76] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_79 
+ bl[77] br[77] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_80 
+ bl[78] br[78] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_81 
+ bl[79] br[79] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_82 
+ bl[80] br[80] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_83 
+ bl[81] br[81] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_84 
+ bl[82] br[82] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_85 
+ bl[83] br[83] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_86 
+ bl[84] br[84] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_87 
+ bl[85] br[85] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_88 
+ bl[86] br[86] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_89 
+ bl[87] br[87] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_90 
+ bl[88] br[88] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_91 
+ bl[89] br[89] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_92 
+ bl[90] br[90] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_93 
+ bl[91] br[91] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_94 
+ bl[92] br[92] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_95 
+ bl[93] br[93] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_96 
+ bl[94] br[94] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_97 
+ bl[95] br[95] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_98 
+ bl[96] br[96] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_99 
+ bl[97] br[97] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_100 
+ bl[98] br[98] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_101 
+ bl[99] br[99] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_102 
+ bl[100] br[100] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_103 
+ bl[101] br[101] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_104 
+ bl[102] br[102] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_105 
+ bl[103] br[103] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_106 
+ bl[104] br[104] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_107 
+ bl[105] br[105] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_108 
+ bl[106] br[106] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_109 
+ bl[107] br[107] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_110 
+ bl[108] br[108] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_111 
+ bl[109] br[109] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_112 
+ bl[110] br[110] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_113 
+ bl[111] br[111] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_114 
+ bl[112] br[112] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_115 
+ bl[113] br[113] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_116 
+ bl[114] br[114] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_117 
+ bl[115] br[115] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_118 
+ bl[116] br[116] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_119 
+ bl[117] br[117] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_120 
+ bl[118] br[118] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_121 
+ bl[119] br[119] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_122 
+ bl[120] br[120] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_123 
+ bl[121] br[121] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_124 
+ bl[122] br[122] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_125 
+ bl[123] br[123] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_126 
+ bl[124] br[124] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_127 
+ bl[125] br[125] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_128 
+ bl[126] br[126] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_129 
+ bl[127] br[127] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_130 
+ bl[128] br[128] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_131 
+ bl[129] br[129] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_132 
+ bl[130] br[130] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_133 
+ bl[131] br[131] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_134 
+ bl[132] br[132] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_135 
+ bl[133] br[133] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_136 
+ bl[134] br[134] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_137 
+ bl[135] br[135] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_138 
+ bl[136] br[136] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_139 
+ bl[137] br[137] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_140 
+ bl[138] br[138] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_141 
+ bl[139] br[139] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_142 
+ bl[140] br[140] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_143 
+ bl[141] br[141] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_144 
+ bl[142] br[142] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_145 
+ bl[143] br[143] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_146 
+ bl[144] br[144] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_147 
+ bl[145] br[145] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_148 
+ bl[146] br[146] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_149 
+ bl[147] br[147] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_150 
+ bl[148] br[148] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_151 
+ bl[149] br[149] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_152 
+ bl[150] br[150] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_153 
+ bl[151] br[151] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_154 
+ bl[152] br[152] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_155 
+ bl[153] br[153] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_156 
+ bl[154] br[154] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_157 
+ bl[155] br[155] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_158 
+ bl[156] br[156] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_159 
+ bl[157] br[157] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_160 
+ bl[158] br[158] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_161 
+ bl[159] br[159] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_162 
+ bl[160] br[160] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_163 
+ bl[161] br[161] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_164 
+ bl[162] br[162] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_165 
+ bl[163] br[163] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_166 
+ bl[164] br[164] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_167 
+ bl[165] br[165] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_168 
+ bl[166] br[166] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_169 
+ bl[167] br[167] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_170 
+ bl[168] br[168] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_171 
+ bl[169] br[169] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_172 
+ bl[170] br[170] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_173 
+ bl[171] br[171] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_174 
+ bl[172] br[172] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_175 
+ bl[173] br[173] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_176 
+ bl[174] br[174] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_177 
+ bl[175] br[175] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_178 
+ bl[176] br[176] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_179 
+ bl[177] br[177] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_180 
+ bl[178] br[178] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_181 
+ bl[179] br[179] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_182 
+ bl[180] br[180] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_183 
+ bl[181] br[181] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_184 
+ bl[182] br[182] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_185 
+ bl[183] br[183] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_186 
+ bl[184] br[184] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_187 
+ bl[185] br[185] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_188 
+ bl[186] br[186] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_189 
+ bl[187] br[187] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_190 
+ bl[188] br[188] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_191 
+ bl[189] br[189] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_192 
+ bl[190] br[190] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_193 
+ bl[191] br[191] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_194 
+ bl[192] br[192] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_195 
+ bl[193] br[193] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_196 
+ bl[194] br[194] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_197 
+ bl[195] br[195] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_198 
+ bl[196] br[196] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_199 
+ bl[197] br[197] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_200 
+ bl[198] br[198] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_201 
+ bl[199] br[199] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_202 
+ bl[200] br[200] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_203 
+ bl[201] br[201] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_204 
+ bl[202] br[202] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_205 
+ bl[203] br[203] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_206 
+ bl[204] br[204] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_207 
+ bl[205] br[205] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_208 
+ bl[206] br[206] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_209 
+ bl[207] br[207] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_210 
+ bl[208] br[208] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_211 
+ bl[209] br[209] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_212 
+ bl[210] br[210] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_213 
+ bl[211] br[211] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_214 
+ bl[212] br[212] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_215 
+ bl[213] br[213] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_216 
+ bl[214] br[214] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_217 
+ bl[215] br[215] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_218 
+ bl[216] br[216] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_219 
+ bl[217] br[217] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_220 
+ bl[218] br[218] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_221 
+ bl[219] br[219] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_222 
+ bl[220] br[220] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_223 
+ bl[221] br[221] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_224 
+ bl[222] br[222] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_225 
+ bl[223] br[223] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_226 
+ bl[224] br[224] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_227 
+ bl[225] br[225] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_228 
+ bl[226] br[226] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_229 
+ bl[227] br[227] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_230 
+ bl[228] br[228] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_231 
+ bl[229] br[229] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_232 
+ bl[230] br[230] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_233 
+ bl[231] br[231] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_234 
+ bl[232] br[232] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_235 
+ bl[233] br[233] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_236 
+ bl[234] br[234] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_237 
+ bl[235] br[235] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_238 
+ bl[236] br[236] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_239 
+ bl[237] br[237] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_240 
+ bl[238] br[238] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_241 
+ bl[239] br[239] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_242 
+ bl[240] br[240] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_243 
+ bl[241] br[241] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_244 
+ bl[242] br[242] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_245 
+ bl[243] br[243] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_246 
+ bl[244] br[244] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_247 
+ bl[245] br[245] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_248 
+ bl[246] br[246] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_249 
+ bl[247] br[247] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_250 
+ bl[248] br[248] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_251 
+ bl[249] br[249] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_252 
+ bl[250] br[250] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_253 
+ bl[251] br[251] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_254 
+ bl[252] br[252] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_255 
+ bl[253] br[253] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_256 
+ bl[254] br[254] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_257 
+ bl[255] br[255] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_258 
+ vdd vdd vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_259 
+ vdd vdd vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_0 
+ vdd vdd vss vdd vpb vnb wl[36] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_38_1 
+ rbl rbr vss vdd vpb vnb wl[36] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_38_2 
+ bl[0] br[0] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_3 
+ bl[1] br[1] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_4 
+ bl[2] br[2] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_5 
+ bl[3] br[3] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_6 
+ bl[4] br[4] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_7 
+ bl[5] br[5] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_8 
+ bl[6] br[6] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_9 
+ bl[7] br[7] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_10 
+ bl[8] br[8] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_11 
+ bl[9] br[9] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_12 
+ bl[10] br[10] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_13 
+ bl[11] br[11] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_14 
+ bl[12] br[12] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_15 
+ bl[13] br[13] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_16 
+ bl[14] br[14] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_17 
+ bl[15] br[15] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_18 
+ bl[16] br[16] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_19 
+ bl[17] br[17] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_20 
+ bl[18] br[18] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_21 
+ bl[19] br[19] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_22 
+ bl[20] br[20] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_23 
+ bl[21] br[21] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_24 
+ bl[22] br[22] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_25 
+ bl[23] br[23] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_26 
+ bl[24] br[24] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_27 
+ bl[25] br[25] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_28 
+ bl[26] br[26] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_29 
+ bl[27] br[27] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_30 
+ bl[28] br[28] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_31 
+ bl[29] br[29] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_32 
+ bl[30] br[30] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_33 
+ bl[31] br[31] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_34 
+ bl[32] br[32] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_35 
+ bl[33] br[33] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_36 
+ bl[34] br[34] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_37 
+ bl[35] br[35] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_38 
+ bl[36] br[36] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_39 
+ bl[37] br[37] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_40 
+ bl[38] br[38] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_41 
+ bl[39] br[39] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_42 
+ bl[40] br[40] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_43 
+ bl[41] br[41] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_44 
+ bl[42] br[42] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_45 
+ bl[43] br[43] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_46 
+ bl[44] br[44] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_47 
+ bl[45] br[45] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_48 
+ bl[46] br[46] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_49 
+ bl[47] br[47] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_50 
+ bl[48] br[48] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_51 
+ bl[49] br[49] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_52 
+ bl[50] br[50] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_53 
+ bl[51] br[51] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_54 
+ bl[52] br[52] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_55 
+ bl[53] br[53] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_56 
+ bl[54] br[54] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_57 
+ bl[55] br[55] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_58 
+ bl[56] br[56] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_59 
+ bl[57] br[57] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_60 
+ bl[58] br[58] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_61 
+ bl[59] br[59] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_62 
+ bl[60] br[60] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_63 
+ bl[61] br[61] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_64 
+ bl[62] br[62] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_65 
+ bl[63] br[63] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_66 
+ bl[64] br[64] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_67 
+ bl[65] br[65] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_68 
+ bl[66] br[66] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_69 
+ bl[67] br[67] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_70 
+ bl[68] br[68] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_71 
+ bl[69] br[69] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_72 
+ bl[70] br[70] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_73 
+ bl[71] br[71] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_74 
+ bl[72] br[72] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_75 
+ bl[73] br[73] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_76 
+ bl[74] br[74] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_77 
+ bl[75] br[75] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_78 
+ bl[76] br[76] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_79 
+ bl[77] br[77] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_80 
+ bl[78] br[78] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_81 
+ bl[79] br[79] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_82 
+ bl[80] br[80] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_83 
+ bl[81] br[81] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_84 
+ bl[82] br[82] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_85 
+ bl[83] br[83] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_86 
+ bl[84] br[84] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_87 
+ bl[85] br[85] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_88 
+ bl[86] br[86] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_89 
+ bl[87] br[87] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_90 
+ bl[88] br[88] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_91 
+ bl[89] br[89] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_92 
+ bl[90] br[90] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_93 
+ bl[91] br[91] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_94 
+ bl[92] br[92] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_95 
+ bl[93] br[93] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_96 
+ bl[94] br[94] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_97 
+ bl[95] br[95] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_98 
+ bl[96] br[96] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_99 
+ bl[97] br[97] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_100 
+ bl[98] br[98] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_101 
+ bl[99] br[99] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_102 
+ bl[100] br[100] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_103 
+ bl[101] br[101] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_104 
+ bl[102] br[102] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_105 
+ bl[103] br[103] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_106 
+ bl[104] br[104] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_107 
+ bl[105] br[105] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_108 
+ bl[106] br[106] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_109 
+ bl[107] br[107] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_110 
+ bl[108] br[108] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_111 
+ bl[109] br[109] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_112 
+ bl[110] br[110] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_113 
+ bl[111] br[111] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_114 
+ bl[112] br[112] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_115 
+ bl[113] br[113] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_116 
+ bl[114] br[114] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_117 
+ bl[115] br[115] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_118 
+ bl[116] br[116] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_119 
+ bl[117] br[117] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_120 
+ bl[118] br[118] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_121 
+ bl[119] br[119] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_122 
+ bl[120] br[120] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_123 
+ bl[121] br[121] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_124 
+ bl[122] br[122] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_125 
+ bl[123] br[123] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_126 
+ bl[124] br[124] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_127 
+ bl[125] br[125] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_128 
+ bl[126] br[126] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_129 
+ bl[127] br[127] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_130 
+ bl[128] br[128] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_131 
+ bl[129] br[129] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_132 
+ bl[130] br[130] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_133 
+ bl[131] br[131] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_134 
+ bl[132] br[132] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_135 
+ bl[133] br[133] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_136 
+ bl[134] br[134] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_137 
+ bl[135] br[135] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_138 
+ bl[136] br[136] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_139 
+ bl[137] br[137] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_140 
+ bl[138] br[138] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_141 
+ bl[139] br[139] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_142 
+ bl[140] br[140] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_143 
+ bl[141] br[141] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_144 
+ bl[142] br[142] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_145 
+ bl[143] br[143] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_146 
+ bl[144] br[144] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_147 
+ bl[145] br[145] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_148 
+ bl[146] br[146] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_149 
+ bl[147] br[147] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_150 
+ bl[148] br[148] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_151 
+ bl[149] br[149] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_152 
+ bl[150] br[150] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_153 
+ bl[151] br[151] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_154 
+ bl[152] br[152] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_155 
+ bl[153] br[153] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_156 
+ bl[154] br[154] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_157 
+ bl[155] br[155] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_158 
+ bl[156] br[156] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_159 
+ bl[157] br[157] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_160 
+ bl[158] br[158] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_161 
+ bl[159] br[159] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_162 
+ bl[160] br[160] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_163 
+ bl[161] br[161] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_164 
+ bl[162] br[162] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_165 
+ bl[163] br[163] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_166 
+ bl[164] br[164] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_167 
+ bl[165] br[165] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_168 
+ bl[166] br[166] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_169 
+ bl[167] br[167] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_170 
+ bl[168] br[168] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_171 
+ bl[169] br[169] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_172 
+ bl[170] br[170] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_173 
+ bl[171] br[171] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_174 
+ bl[172] br[172] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_175 
+ bl[173] br[173] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_176 
+ bl[174] br[174] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_177 
+ bl[175] br[175] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_178 
+ bl[176] br[176] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_179 
+ bl[177] br[177] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_180 
+ bl[178] br[178] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_181 
+ bl[179] br[179] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_182 
+ bl[180] br[180] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_183 
+ bl[181] br[181] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_184 
+ bl[182] br[182] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_185 
+ bl[183] br[183] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_186 
+ bl[184] br[184] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_187 
+ bl[185] br[185] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_188 
+ bl[186] br[186] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_189 
+ bl[187] br[187] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_190 
+ bl[188] br[188] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_191 
+ bl[189] br[189] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_192 
+ bl[190] br[190] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_193 
+ bl[191] br[191] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_194 
+ bl[192] br[192] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_195 
+ bl[193] br[193] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_196 
+ bl[194] br[194] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_197 
+ bl[195] br[195] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_198 
+ bl[196] br[196] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_199 
+ bl[197] br[197] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_200 
+ bl[198] br[198] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_201 
+ bl[199] br[199] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_202 
+ bl[200] br[200] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_203 
+ bl[201] br[201] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_204 
+ bl[202] br[202] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_205 
+ bl[203] br[203] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_206 
+ bl[204] br[204] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_207 
+ bl[205] br[205] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_208 
+ bl[206] br[206] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_209 
+ bl[207] br[207] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_210 
+ bl[208] br[208] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_211 
+ bl[209] br[209] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_212 
+ bl[210] br[210] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_213 
+ bl[211] br[211] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_214 
+ bl[212] br[212] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_215 
+ bl[213] br[213] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_216 
+ bl[214] br[214] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_217 
+ bl[215] br[215] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_218 
+ bl[216] br[216] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_219 
+ bl[217] br[217] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_220 
+ bl[218] br[218] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_221 
+ bl[219] br[219] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_222 
+ bl[220] br[220] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_223 
+ bl[221] br[221] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_224 
+ bl[222] br[222] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_225 
+ bl[223] br[223] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_226 
+ bl[224] br[224] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_227 
+ bl[225] br[225] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_228 
+ bl[226] br[226] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_229 
+ bl[227] br[227] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_230 
+ bl[228] br[228] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_231 
+ bl[229] br[229] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_232 
+ bl[230] br[230] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_233 
+ bl[231] br[231] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_234 
+ bl[232] br[232] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_235 
+ bl[233] br[233] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_236 
+ bl[234] br[234] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_237 
+ bl[235] br[235] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_238 
+ bl[236] br[236] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_239 
+ bl[237] br[237] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_240 
+ bl[238] br[238] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_241 
+ bl[239] br[239] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_242 
+ bl[240] br[240] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_243 
+ bl[241] br[241] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_244 
+ bl[242] br[242] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_245 
+ bl[243] br[243] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_246 
+ bl[244] br[244] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_247 
+ bl[245] br[245] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_248 
+ bl[246] br[246] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_249 
+ bl[247] br[247] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_250 
+ bl[248] br[248] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_251 
+ bl[249] br[249] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_252 
+ bl[250] br[250] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_253 
+ bl[251] br[251] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_254 
+ bl[252] br[252] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_255 
+ bl[253] br[253] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_256 
+ bl[254] br[254] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_257 
+ bl[255] br[255] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_258 
+ vdd vdd vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_259 
+ vdd vdd vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_0 
+ vdd vdd vss vdd vpb vnb wl[37] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_39_1 
+ rbl rbr vss vdd vpb vnb wl[37] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_39_2 
+ bl[0] br[0] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_3 
+ bl[1] br[1] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_4 
+ bl[2] br[2] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_5 
+ bl[3] br[3] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_6 
+ bl[4] br[4] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_7 
+ bl[5] br[5] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_8 
+ bl[6] br[6] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_9 
+ bl[7] br[7] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_10 
+ bl[8] br[8] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_11 
+ bl[9] br[9] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_12 
+ bl[10] br[10] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_13 
+ bl[11] br[11] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_14 
+ bl[12] br[12] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_15 
+ bl[13] br[13] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_16 
+ bl[14] br[14] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_17 
+ bl[15] br[15] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_18 
+ bl[16] br[16] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_19 
+ bl[17] br[17] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_20 
+ bl[18] br[18] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_21 
+ bl[19] br[19] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_22 
+ bl[20] br[20] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_23 
+ bl[21] br[21] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_24 
+ bl[22] br[22] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_25 
+ bl[23] br[23] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_26 
+ bl[24] br[24] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_27 
+ bl[25] br[25] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_28 
+ bl[26] br[26] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_29 
+ bl[27] br[27] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_30 
+ bl[28] br[28] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_31 
+ bl[29] br[29] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_32 
+ bl[30] br[30] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_33 
+ bl[31] br[31] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_34 
+ bl[32] br[32] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_35 
+ bl[33] br[33] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_36 
+ bl[34] br[34] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_37 
+ bl[35] br[35] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_38 
+ bl[36] br[36] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_39 
+ bl[37] br[37] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_40 
+ bl[38] br[38] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_41 
+ bl[39] br[39] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_42 
+ bl[40] br[40] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_43 
+ bl[41] br[41] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_44 
+ bl[42] br[42] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_45 
+ bl[43] br[43] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_46 
+ bl[44] br[44] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_47 
+ bl[45] br[45] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_48 
+ bl[46] br[46] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_49 
+ bl[47] br[47] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_50 
+ bl[48] br[48] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_51 
+ bl[49] br[49] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_52 
+ bl[50] br[50] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_53 
+ bl[51] br[51] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_54 
+ bl[52] br[52] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_55 
+ bl[53] br[53] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_56 
+ bl[54] br[54] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_57 
+ bl[55] br[55] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_58 
+ bl[56] br[56] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_59 
+ bl[57] br[57] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_60 
+ bl[58] br[58] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_61 
+ bl[59] br[59] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_62 
+ bl[60] br[60] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_63 
+ bl[61] br[61] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_64 
+ bl[62] br[62] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_65 
+ bl[63] br[63] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_66 
+ bl[64] br[64] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_67 
+ bl[65] br[65] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_68 
+ bl[66] br[66] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_69 
+ bl[67] br[67] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_70 
+ bl[68] br[68] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_71 
+ bl[69] br[69] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_72 
+ bl[70] br[70] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_73 
+ bl[71] br[71] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_74 
+ bl[72] br[72] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_75 
+ bl[73] br[73] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_76 
+ bl[74] br[74] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_77 
+ bl[75] br[75] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_78 
+ bl[76] br[76] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_79 
+ bl[77] br[77] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_80 
+ bl[78] br[78] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_81 
+ bl[79] br[79] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_82 
+ bl[80] br[80] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_83 
+ bl[81] br[81] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_84 
+ bl[82] br[82] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_85 
+ bl[83] br[83] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_86 
+ bl[84] br[84] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_87 
+ bl[85] br[85] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_88 
+ bl[86] br[86] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_89 
+ bl[87] br[87] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_90 
+ bl[88] br[88] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_91 
+ bl[89] br[89] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_92 
+ bl[90] br[90] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_93 
+ bl[91] br[91] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_94 
+ bl[92] br[92] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_95 
+ bl[93] br[93] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_96 
+ bl[94] br[94] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_97 
+ bl[95] br[95] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_98 
+ bl[96] br[96] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_99 
+ bl[97] br[97] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_100 
+ bl[98] br[98] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_101 
+ bl[99] br[99] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_102 
+ bl[100] br[100] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_103 
+ bl[101] br[101] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_104 
+ bl[102] br[102] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_105 
+ bl[103] br[103] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_106 
+ bl[104] br[104] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_107 
+ bl[105] br[105] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_108 
+ bl[106] br[106] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_109 
+ bl[107] br[107] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_110 
+ bl[108] br[108] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_111 
+ bl[109] br[109] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_112 
+ bl[110] br[110] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_113 
+ bl[111] br[111] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_114 
+ bl[112] br[112] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_115 
+ bl[113] br[113] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_116 
+ bl[114] br[114] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_117 
+ bl[115] br[115] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_118 
+ bl[116] br[116] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_119 
+ bl[117] br[117] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_120 
+ bl[118] br[118] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_121 
+ bl[119] br[119] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_122 
+ bl[120] br[120] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_123 
+ bl[121] br[121] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_124 
+ bl[122] br[122] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_125 
+ bl[123] br[123] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_126 
+ bl[124] br[124] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_127 
+ bl[125] br[125] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_128 
+ bl[126] br[126] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_129 
+ bl[127] br[127] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_130 
+ bl[128] br[128] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_131 
+ bl[129] br[129] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_132 
+ bl[130] br[130] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_133 
+ bl[131] br[131] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_134 
+ bl[132] br[132] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_135 
+ bl[133] br[133] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_136 
+ bl[134] br[134] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_137 
+ bl[135] br[135] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_138 
+ bl[136] br[136] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_139 
+ bl[137] br[137] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_140 
+ bl[138] br[138] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_141 
+ bl[139] br[139] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_142 
+ bl[140] br[140] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_143 
+ bl[141] br[141] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_144 
+ bl[142] br[142] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_145 
+ bl[143] br[143] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_146 
+ bl[144] br[144] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_147 
+ bl[145] br[145] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_148 
+ bl[146] br[146] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_149 
+ bl[147] br[147] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_150 
+ bl[148] br[148] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_151 
+ bl[149] br[149] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_152 
+ bl[150] br[150] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_153 
+ bl[151] br[151] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_154 
+ bl[152] br[152] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_155 
+ bl[153] br[153] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_156 
+ bl[154] br[154] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_157 
+ bl[155] br[155] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_158 
+ bl[156] br[156] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_159 
+ bl[157] br[157] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_160 
+ bl[158] br[158] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_161 
+ bl[159] br[159] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_162 
+ bl[160] br[160] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_163 
+ bl[161] br[161] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_164 
+ bl[162] br[162] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_165 
+ bl[163] br[163] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_166 
+ bl[164] br[164] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_167 
+ bl[165] br[165] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_168 
+ bl[166] br[166] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_169 
+ bl[167] br[167] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_170 
+ bl[168] br[168] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_171 
+ bl[169] br[169] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_172 
+ bl[170] br[170] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_173 
+ bl[171] br[171] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_174 
+ bl[172] br[172] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_175 
+ bl[173] br[173] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_176 
+ bl[174] br[174] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_177 
+ bl[175] br[175] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_178 
+ bl[176] br[176] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_179 
+ bl[177] br[177] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_180 
+ bl[178] br[178] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_181 
+ bl[179] br[179] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_182 
+ bl[180] br[180] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_183 
+ bl[181] br[181] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_184 
+ bl[182] br[182] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_185 
+ bl[183] br[183] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_186 
+ bl[184] br[184] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_187 
+ bl[185] br[185] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_188 
+ bl[186] br[186] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_189 
+ bl[187] br[187] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_190 
+ bl[188] br[188] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_191 
+ bl[189] br[189] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_192 
+ bl[190] br[190] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_193 
+ bl[191] br[191] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_194 
+ bl[192] br[192] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_195 
+ bl[193] br[193] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_196 
+ bl[194] br[194] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_197 
+ bl[195] br[195] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_198 
+ bl[196] br[196] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_199 
+ bl[197] br[197] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_200 
+ bl[198] br[198] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_201 
+ bl[199] br[199] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_202 
+ bl[200] br[200] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_203 
+ bl[201] br[201] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_204 
+ bl[202] br[202] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_205 
+ bl[203] br[203] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_206 
+ bl[204] br[204] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_207 
+ bl[205] br[205] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_208 
+ bl[206] br[206] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_209 
+ bl[207] br[207] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_210 
+ bl[208] br[208] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_211 
+ bl[209] br[209] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_212 
+ bl[210] br[210] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_213 
+ bl[211] br[211] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_214 
+ bl[212] br[212] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_215 
+ bl[213] br[213] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_216 
+ bl[214] br[214] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_217 
+ bl[215] br[215] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_218 
+ bl[216] br[216] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_219 
+ bl[217] br[217] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_220 
+ bl[218] br[218] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_221 
+ bl[219] br[219] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_222 
+ bl[220] br[220] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_223 
+ bl[221] br[221] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_224 
+ bl[222] br[222] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_225 
+ bl[223] br[223] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_226 
+ bl[224] br[224] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_227 
+ bl[225] br[225] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_228 
+ bl[226] br[226] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_229 
+ bl[227] br[227] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_230 
+ bl[228] br[228] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_231 
+ bl[229] br[229] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_232 
+ bl[230] br[230] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_233 
+ bl[231] br[231] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_234 
+ bl[232] br[232] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_235 
+ bl[233] br[233] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_236 
+ bl[234] br[234] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_237 
+ bl[235] br[235] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_238 
+ bl[236] br[236] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_239 
+ bl[237] br[237] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_240 
+ bl[238] br[238] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_241 
+ bl[239] br[239] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_242 
+ bl[240] br[240] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_243 
+ bl[241] br[241] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_244 
+ bl[242] br[242] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_245 
+ bl[243] br[243] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_246 
+ bl[244] br[244] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_247 
+ bl[245] br[245] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_248 
+ bl[246] br[246] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_249 
+ bl[247] br[247] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_250 
+ bl[248] br[248] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_251 
+ bl[249] br[249] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_252 
+ bl[250] br[250] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_253 
+ bl[251] br[251] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_254 
+ bl[252] br[252] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_255 
+ bl[253] br[253] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_256 
+ bl[254] br[254] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_257 
+ bl[255] br[255] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_258 
+ vdd vdd vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_259 
+ vdd vdd vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_0 
+ vdd vdd vss vdd vpb vnb wl[38] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_40_1 
+ rbl rbr vss vdd vpb vnb wl[38] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_40_2 
+ bl[0] br[0] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_3 
+ bl[1] br[1] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_4 
+ bl[2] br[2] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_5 
+ bl[3] br[3] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_6 
+ bl[4] br[4] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_7 
+ bl[5] br[5] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_8 
+ bl[6] br[6] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_9 
+ bl[7] br[7] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_10 
+ bl[8] br[8] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_11 
+ bl[9] br[9] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_12 
+ bl[10] br[10] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_13 
+ bl[11] br[11] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_14 
+ bl[12] br[12] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_15 
+ bl[13] br[13] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_16 
+ bl[14] br[14] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_17 
+ bl[15] br[15] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_18 
+ bl[16] br[16] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_19 
+ bl[17] br[17] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_20 
+ bl[18] br[18] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_21 
+ bl[19] br[19] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_22 
+ bl[20] br[20] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_23 
+ bl[21] br[21] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_24 
+ bl[22] br[22] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_25 
+ bl[23] br[23] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_26 
+ bl[24] br[24] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_27 
+ bl[25] br[25] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_28 
+ bl[26] br[26] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_29 
+ bl[27] br[27] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_30 
+ bl[28] br[28] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_31 
+ bl[29] br[29] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_32 
+ bl[30] br[30] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_33 
+ bl[31] br[31] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_34 
+ bl[32] br[32] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_35 
+ bl[33] br[33] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_36 
+ bl[34] br[34] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_37 
+ bl[35] br[35] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_38 
+ bl[36] br[36] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_39 
+ bl[37] br[37] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_40 
+ bl[38] br[38] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_41 
+ bl[39] br[39] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_42 
+ bl[40] br[40] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_43 
+ bl[41] br[41] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_44 
+ bl[42] br[42] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_45 
+ bl[43] br[43] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_46 
+ bl[44] br[44] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_47 
+ bl[45] br[45] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_48 
+ bl[46] br[46] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_49 
+ bl[47] br[47] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_50 
+ bl[48] br[48] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_51 
+ bl[49] br[49] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_52 
+ bl[50] br[50] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_53 
+ bl[51] br[51] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_54 
+ bl[52] br[52] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_55 
+ bl[53] br[53] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_56 
+ bl[54] br[54] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_57 
+ bl[55] br[55] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_58 
+ bl[56] br[56] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_59 
+ bl[57] br[57] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_60 
+ bl[58] br[58] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_61 
+ bl[59] br[59] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_62 
+ bl[60] br[60] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_63 
+ bl[61] br[61] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_64 
+ bl[62] br[62] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_65 
+ bl[63] br[63] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_66 
+ bl[64] br[64] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_67 
+ bl[65] br[65] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_68 
+ bl[66] br[66] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_69 
+ bl[67] br[67] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_70 
+ bl[68] br[68] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_71 
+ bl[69] br[69] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_72 
+ bl[70] br[70] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_73 
+ bl[71] br[71] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_74 
+ bl[72] br[72] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_75 
+ bl[73] br[73] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_76 
+ bl[74] br[74] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_77 
+ bl[75] br[75] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_78 
+ bl[76] br[76] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_79 
+ bl[77] br[77] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_80 
+ bl[78] br[78] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_81 
+ bl[79] br[79] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_82 
+ bl[80] br[80] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_83 
+ bl[81] br[81] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_84 
+ bl[82] br[82] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_85 
+ bl[83] br[83] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_86 
+ bl[84] br[84] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_87 
+ bl[85] br[85] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_88 
+ bl[86] br[86] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_89 
+ bl[87] br[87] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_90 
+ bl[88] br[88] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_91 
+ bl[89] br[89] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_92 
+ bl[90] br[90] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_93 
+ bl[91] br[91] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_94 
+ bl[92] br[92] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_95 
+ bl[93] br[93] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_96 
+ bl[94] br[94] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_97 
+ bl[95] br[95] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_98 
+ bl[96] br[96] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_99 
+ bl[97] br[97] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_100 
+ bl[98] br[98] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_101 
+ bl[99] br[99] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_102 
+ bl[100] br[100] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_103 
+ bl[101] br[101] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_104 
+ bl[102] br[102] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_105 
+ bl[103] br[103] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_106 
+ bl[104] br[104] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_107 
+ bl[105] br[105] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_108 
+ bl[106] br[106] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_109 
+ bl[107] br[107] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_110 
+ bl[108] br[108] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_111 
+ bl[109] br[109] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_112 
+ bl[110] br[110] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_113 
+ bl[111] br[111] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_114 
+ bl[112] br[112] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_115 
+ bl[113] br[113] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_116 
+ bl[114] br[114] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_117 
+ bl[115] br[115] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_118 
+ bl[116] br[116] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_119 
+ bl[117] br[117] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_120 
+ bl[118] br[118] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_121 
+ bl[119] br[119] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_122 
+ bl[120] br[120] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_123 
+ bl[121] br[121] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_124 
+ bl[122] br[122] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_125 
+ bl[123] br[123] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_126 
+ bl[124] br[124] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_127 
+ bl[125] br[125] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_128 
+ bl[126] br[126] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_129 
+ bl[127] br[127] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_130 
+ bl[128] br[128] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_131 
+ bl[129] br[129] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_132 
+ bl[130] br[130] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_133 
+ bl[131] br[131] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_134 
+ bl[132] br[132] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_135 
+ bl[133] br[133] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_136 
+ bl[134] br[134] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_137 
+ bl[135] br[135] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_138 
+ bl[136] br[136] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_139 
+ bl[137] br[137] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_140 
+ bl[138] br[138] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_141 
+ bl[139] br[139] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_142 
+ bl[140] br[140] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_143 
+ bl[141] br[141] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_144 
+ bl[142] br[142] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_145 
+ bl[143] br[143] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_146 
+ bl[144] br[144] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_147 
+ bl[145] br[145] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_148 
+ bl[146] br[146] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_149 
+ bl[147] br[147] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_150 
+ bl[148] br[148] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_151 
+ bl[149] br[149] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_152 
+ bl[150] br[150] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_153 
+ bl[151] br[151] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_154 
+ bl[152] br[152] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_155 
+ bl[153] br[153] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_156 
+ bl[154] br[154] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_157 
+ bl[155] br[155] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_158 
+ bl[156] br[156] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_159 
+ bl[157] br[157] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_160 
+ bl[158] br[158] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_161 
+ bl[159] br[159] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_162 
+ bl[160] br[160] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_163 
+ bl[161] br[161] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_164 
+ bl[162] br[162] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_165 
+ bl[163] br[163] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_166 
+ bl[164] br[164] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_167 
+ bl[165] br[165] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_168 
+ bl[166] br[166] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_169 
+ bl[167] br[167] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_170 
+ bl[168] br[168] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_171 
+ bl[169] br[169] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_172 
+ bl[170] br[170] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_173 
+ bl[171] br[171] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_174 
+ bl[172] br[172] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_175 
+ bl[173] br[173] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_176 
+ bl[174] br[174] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_177 
+ bl[175] br[175] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_178 
+ bl[176] br[176] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_179 
+ bl[177] br[177] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_180 
+ bl[178] br[178] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_181 
+ bl[179] br[179] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_182 
+ bl[180] br[180] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_183 
+ bl[181] br[181] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_184 
+ bl[182] br[182] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_185 
+ bl[183] br[183] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_186 
+ bl[184] br[184] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_187 
+ bl[185] br[185] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_188 
+ bl[186] br[186] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_189 
+ bl[187] br[187] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_190 
+ bl[188] br[188] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_191 
+ bl[189] br[189] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_192 
+ bl[190] br[190] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_193 
+ bl[191] br[191] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_194 
+ bl[192] br[192] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_195 
+ bl[193] br[193] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_196 
+ bl[194] br[194] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_197 
+ bl[195] br[195] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_198 
+ bl[196] br[196] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_199 
+ bl[197] br[197] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_200 
+ bl[198] br[198] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_201 
+ bl[199] br[199] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_202 
+ bl[200] br[200] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_203 
+ bl[201] br[201] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_204 
+ bl[202] br[202] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_205 
+ bl[203] br[203] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_206 
+ bl[204] br[204] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_207 
+ bl[205] br[205] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_208 
+ bl[206] br[206] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_209 
+ bl[207] br[207] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_210 
+ bl[208] br[208] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_211 
+ bl[209] br[209] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_212 
+ bl[210] br[210] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_213 
+ bl[211] br[211] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_214 
+ bl[212] br[212] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_215 
+ bl[213] br[213] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_216 
+ bl[214] br[214] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_217 
+ bl[215] br[215] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_218 
+ bl[216] br[216] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_219 
+ bl[217] br[217] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_220 
+ bl[218] br[218] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_221 
+ bl[219] br[219] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_222 
+ bl[220] br[220] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_223 
+ bl[221] br[221] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_224 
+ bl[222] br[222] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_225 
+ bl[223] br[223] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_226 
+ bl[224] br[224] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_227 
+ bl[225] br[225] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_228 
+ bl[226] br[226] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_229 
+ bl[227] br[227] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_230 
+ bl[228] br[228] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_231 
+ bl[229] br[229] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_232 
+ bl[230] br[230] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_233 
+ bl[231] br[231] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_234 
+ bl[232] br[232] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_235 
+ bl[233] br[233] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_236 
+ bl[234] br[234] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_237 
+ bl[235] br[235] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_238 
+ bl[236] br[236] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_239 
+ bl[237] br[237] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_240 
+ bl[238] br[238] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_241 
+ bl[239] br[239] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_242 
+ bl[240] br[240] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_243 
+ bl[241] br[241] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_244 
+ bl[242] br[242] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_245 
+ bl[243] br[243] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_246 
+ bl[244] br[244] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_247 
+ bl[245] br[245] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_248 
+ bl[246] br[246] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_249 
+ bl[247] br[247] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_250 
+ bl[248] br[248] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_251 
+ bl[249] br[249] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_252 
+ bl[250] br[250] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_253 
+ bl[251] br[251] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_254 
+ bl[252] br[252] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_255 
+ bl[253] br[253] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_256 
+ bl[254] br[254] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_257 
+ bl[255] br[255] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_258 
+ vdd vdd vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_259 
+ vdd vdd vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_0 
+ vdd vdd vss vdd vpb vnb wl[39] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_41_1 
+ rbl rbr vss vdd vpb vnb wl[39] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_41_2 
+ bl[0] br[0] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_3 
+ bl[1] br[1] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_4 
+ bl[2] br[2] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_5 
+ bl[3] br[3] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_6 
+ bl[4] br[4] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_7 
+ bl[5] br[5] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_8 
+ bl[6] br[6] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_9 
+ bl[7] br[7] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_10 
+ bl[8] br[8] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_11 
+ bl[9] br[9] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_12 
+ bl[10] br[10] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_13 
+ bl[11] br[11] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_14 
+ bl[12] br[12] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_15 
+ bl[13] br[13] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_16 
+ bl[14] br[14] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_17 
+ bl[15] br[15] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_18 
+ bl[16] br[16] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_19 
+ bl[17] br[17] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_20 
+ bl[18] br[18] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_21 
+ bl[19] br[19] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_22 
+ bl[20] br[20] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_23 
+ bl[21] br[21] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_24 
+ bl[22] br[22] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_25 
+ bl[23] br[23] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_26 
+ bl[24] br[24] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_27 
+ bl[25] br[25] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_28 
+ bl[26] br[26] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_29 
+ bl[27] br[27] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_30 
+ bl[28] br[28] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_31 
+ bl[29] br[29] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_32 
+ bl[30] br[30] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_33 
+ bl[31] br[31] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_34 
+ bl[32] br[32] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_35 
+ bl[33] br[33] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_36 
+ bl[34] br[34] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_37 
+ bl[35] br[35] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_38 
+ bl[36] br[36] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_39 
+ bl[37] br[37] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_40 
+ bl[38] br[38] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_41 
+ bl[39] br[39] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_42 
+ bl[40] br[40] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_43 
+ bl[41] br[41] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_44 
+ bl[42] br[42] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_45 
+ bl[43] br[43] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_46 
+ bl[44] br[44] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_47 
+ bl[45] br[45] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_48 
+ bl[46] br[46] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_49 
+ bl[47] br[47] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_50 
+ bl[48] br[48] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_51 
+ bl[49] br[49] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_52 
+ bl[50] br[50] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_53 
+ bl[51] br[51] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_54 
+ bl[52] br[52] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_55 
+ bl[53] br[53] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_56 
+ bl[54] br[54] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_57 
+ bl[55] br[55] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_58 
+ bl[56] br[56] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_59 
+ bl[57] br[57] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_60 
+ bl[58] br[58] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_61 
+ bl[59] br[59] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_62 
+ bl[60] br[60] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_63 
+ bl[61] br[61] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_64 
+ bl[62] br[62] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_65 
+ bl[63] br[63] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_66 
+ bl[64] br[64] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_67 
+ bl[65] br[65] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_68 
+ bl[66] br[66] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_69 
+ bl[67] br[67] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_70 
+ bl[68] br[68] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_71 
+ bl[69] br[69] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_72 
+ bl[70] br[70] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_73 
+ bl[71] br[71] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_74 
+ bl[72] br[72] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_75 
+ bl[73] br[73] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_76 
+ bl[74] br[74] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_77 
+ bl[75] br[75] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_78 
+ bl[76] br[76] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_79 
+ bl[77] br[77] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_80 
+ bl[78] br[78] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_81 
+ bl[79] br[79] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_82 
+ bl[80] br[80] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_83 
+ bl[81] br[81] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_84 
+ bl[82] br[82] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_85 
+ bl[83] br[83] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_86 
+ bl[84] br[84] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_87 
+ bl[85] br[85] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_88 
+ bl[86] br[86] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_89 
+ bl[87] br[87] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_90 
+ bl[88] br[88] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_91 
+ bl[89] br[89] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_92 
+ bl[90] br[90] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_93 
+ bl[91] br[91] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_94 
+ bl[92] br[92] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_95 
+ bl[93] br[93] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_96 
+ bl[94] br[94] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_97 
+ bl[95] br[95] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_98 
+ bl[96] br[96] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_99 
+ bl[97] br[97] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_100 
+ bl[98] br[98] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_101 
+ bl[99] br[99] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_102 
+ bl[100] br[100] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_103 
+ bl[101] br[101] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_104 
+ bl[102] br[102] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_105 
+ bl[103] br[103] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_106 
+ bl[104] br[104] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_107 
+ bl[105] br[105] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_108 
+ bl[106] br[106] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_109 
+ bl[107] br[107] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_110 
+ bl[108] br[108] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_111 
+ bl[109] br[109] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_112 
+ bl[110] br[110] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_113 
+ bl[111] br[111] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_114 
+ bl[112] br[112] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_115 
+ bl[113] br[113] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_116 
+ bl[114] br[114] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_117 
+ bl[115] br[115] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_118 
+ bl[116] br[116] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_119 
+ bl[117] br[117] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_120 
+ bl[118] br[118] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_121 
+ bl[119] br[119] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_122 
+ bl[120] br[120] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_123 
+ bl[121] br[121] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_124 
+ bl[122] br[122] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_125 
+ bl[123] br[123] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_126 
+ bl[124] br[124] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_127 
+ bl[125] br[125] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_128 
+ bl[126] br[126] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_129 
+ bl[127] br[127] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_130 
+ bl[128] br[128] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_131 
+ bl[129] br[129] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_132 
+ bl[130] br[130] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_133 
+ bl[131] br[131] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_134 
+ bl[132] br[132] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_135 
+ bl[133] br[133] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_136 
+ bl[134] br[134] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_137 
+ bl[135] br[135] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_138 
+ bl[136] br[136] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_139 
+ bl[137] br[137] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_140 
+ bl[138] br[138] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_141 
+ bl[139] br[139] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_142 
+ bl[140] br[140] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_143 
+ bl[141] br[141] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_144 
+ bl[142] br[142] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_145 
+ bl[143] br[143] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_146 
+ bl[144] br[144] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_147 
+ bl[145] br[145] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_148 
+ bl[146] br[146] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_149 
+ bl[147] br[147] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_150 
+ bl[148] br[148] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_151 
+ bl[149] br[149] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_152 
+ bl[150] br[150] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_153 
+ bl[151] br[151] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_154 
+ bl[152] br[152] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_155 
+ bl[153] br[153] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_156 
+ bl[154] br[154] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_157 
+ bl[155] br[155] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_158 
+ bl[156] br[156] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_159 
+ bl[157] br[157] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_160 
+ bl[158] br[158] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_161 
+ bl[159] br[159] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_162 
+ bl[160] br[160] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_163 
+ bl[161] br[161] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_164 
+ bl[162] br[162] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_165 
+ bl[163] br[163] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_166 
+ bl[164] br[164] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_167 
+ bl[165] br[165] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_168 
+ bl[166] br[166] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_169 
+ bl[167] br[167] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_170 
+ bl[168] br[168] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_171 
+ bl[169] br[169] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_172 
+ bl[170] br[170] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_173 
+ bl[171] br[171] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_174 
+ bl[172] br[172] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_175 
+ bl[173] br[173] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_176 
+ bl[174] br[174] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_177 
+ bl[175] br[175] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_178 
+ bl[176] br[176] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_179 
+ bl[177] br[177] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_180 
+ bl[178] br[178] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_181 
+ bl[179] br[179] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_182 
+ bl[180] br[180] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_183 
+ bl[181] br[181] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_184 
+ bl[182] br[182] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_185 
+ bl[183] br[183] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_186 
+ bl[184] br[184] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_187 
+ bl[185] br[185] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_188 
+ bl[186] br[186] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_189 
+ bl[187] br[187] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_190 
+ bl[188] br[188] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_191 
+ bl[189] br[189] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_192 
+ bl[190] br[190] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_193 
+ bl[191] br[191] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_194 
+ bl[192] br[192] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_195 
+ bl[193] br[193] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_196 
+ bl[194] br[194] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_197 
+ bl[195] br[195] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_198 
+ bl[196] br[196] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_199 
+ bl[197] br[197] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_200 
+ bl[198] br[198] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_201 
+ bl[199] br[199] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_202 
+ bl[200] br[200] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_203 
+ bl[201] br[201] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_204 
+ bl[202] br[202] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_205 
+ bl[203] br[203] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_206 
+ bl[204] br[204] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_207 
+ bl[205] br[205] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_208 
+ bl[206] br[206] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_209 
+ bl[207] br[207] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_210 
+ bl[208] br[208] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_211 
+ bl[209] br[209] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_212 
+ bl[210] br[210] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_213 
+ bl[211] br[211] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_214 
+ bl[212] br[212] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_215 
+ bl[213] br[213] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_216 
+ bl[214] br[214] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_217 
+ bl[215] br[215] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_218 
+ bl[216] br[216] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_219 
+ bl[217] br[217] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_220 
+ bl[218] br[218] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_221 
+ bl[219] br[219] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_222 
+ bl[220] br[220] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_223 
+ bl[221] br[221] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_224 
+ bl[222] br[222] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_225 
+ bl[223] br[223] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_226 
+ bl[224] br[224] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_227 
+ bl[225] br[225] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_228 
+ bl[226] br[226] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_229 
+ bl[227] br[227] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_230 
+ bl[228] br[228] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_231 
+ bl[229] br[229] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_232 
+ bl[230] br[230] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_233 
+ bl[231] br[231] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_234 
+ bl[232] br[232] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_235 
+ bl[233] br[233] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_236 
+ bl[234] br[234] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_237 
+ bl[235] br[235] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_238 
+ bl[236] br[236] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_239 
+ bl[237] br[237] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_240 
+ bl[238] br[238] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_241 
+ bl[239] br[239] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_242 
+ bl[240] br[240] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_243 
+ bl[241] br[241] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_244 
+ bl[242] br[242] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_245 
+ bl[243] br[243] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_246 
+ bl[244] br[244] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_247 
+ bl[245] br[245] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_248 
+ bl[246] br[246] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_249 
+ bl[247] br[247] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_250 
+ bl[248] br[248] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_251 
+ bl[249] br[249] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_252 
+ bl[250] br[250] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_253 
+ bl[251] br[251] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_254 
+ bl[252] br[252] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_255 
+ bl[253] br[253] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_256 
+ bl[254] br[254] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_257 
+ bl[255] br[255] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_258 
+ vdd vdd vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_259 
+ vdd vdd vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_0 
+ vdd vdd vss vdd vpb vnb wl[40] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_42_1 
+ rbl rbr vss vdd vpb vnb wl[40] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_42_2 
+ bl[0] br[0] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_3 
+ bl[1] br[1] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_4 
+ bl[2] br[2] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_5 
+ bl[3] br[3] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_6 
+ bl[4] br[4] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_7 
+ bl[5] br[5] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_8 
+ bl[6] br[6] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_9 
+ bl[7] br[7] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_10 
+ bl[8] br[8] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_11 
+ bl[9] br[9] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_12 
+ bl[10] br[10] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_13 
+ bl[11] br[11] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_14 
+ bl[12] br[12] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_15 
+ bl[13] br[13] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_16 
+ bl[14] br[14] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_17 
+ bl[15] br[15] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_18 
+ bl[16] br[16] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_19 
+ bl[17] br[17] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_20 
+ bl[18] br[18] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_21 
+ bl[19] br[19] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_22 
+ bl[20] br[20] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_23 
+ bl[21] br[21] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_24 
+ bl[22] br[22] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_25 
+ bl[23] br[23] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_26 
+ bl[24] br[24] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_27 
+ bl[25] br[25] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_28 
+ bl[26] br[26] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_29 
+ bl[27] br[27] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_30 
+ bl[28] br[28] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_31 
+ bl[29] br[29] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_32 
+ bl[30] br[30] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_33 
+ bl[31] br[31] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_34 
+ bl[32] br[32] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_35 
+ bl[33] br[33] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_36 
+ bl[34] br[34] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_37 
+ bl[35] br[35] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_38 
+ bl[36] br[36] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_39 
+ bl[37] br[37] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_40 
+ bl[38] br[38] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_41 
+ bl[39] br[39] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_42 
+ bl[40] br[40] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_43 
+ bl[41] br[41] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_44 
+ bl[42] br[42] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_45 
+ bl[43] br[43] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_46 
+ bl[44] br[44] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_47 
+ bl[45] br[45] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_48 
+ bl[46] br[46] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_49 
+ bl[47] br[47] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_50 
+ bl[48] br[48] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_51 
+ bl[49] br[49] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_52 
+ bl[50] br[50] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_53 
+ bl[51] br[51] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_54 
+ bl[52] br[52] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_55 
+ bl[53] br[53] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_56 
+ bl[54] br[54] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_57 
+ bl[55] br[55] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_58 
+ bl[56] br[56] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_59 
+ bl[57] br[57] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_60 
+ bl[58] br[58] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_61 
+ bl[59] br[59] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_62 
+ bl[60] br[60] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_63 
+ bl[61] br[61] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_64 
+ bl[62] br[62] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_65 
+ bl[63] br[63] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_66 
+ bl[64] br[64] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_67 
+ bl[65] br[65] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_68 
+ bl[66] br[66] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_69 
+ bl[67] br[67] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_70 
+ bl[68] br[68] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_71 
+ bl[69] br[69] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_72 
+ bl[70] br[70] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_73 
+ bl[71] br[71] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_74 
+ bl[72] br[72] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_75 
+ bl[73] br[73] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_76 
+ bl[74] br[74] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_77 
+ bl[75] br[75] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_78 
+ bl[76] br[76] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_79 
+ bl[77] br[77] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_80 
+ bl[78] br[78] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_81 
+ bl[79] br[79] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_82 
+ bl[80] br[80] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_83 
+ bl[81] br[81] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_84 
+ bl[82] br[82] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_85 
+ bl[83] br[83] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_86 
+ bl[84] br[84] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_87 
+ bl[85] br[85] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_88 
+ bl[86] br[86] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_89 
+ bl[87] br[87] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_90 
+ bl[88] br[88] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_91 
+ bl[89] br[89] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_92 
+ bl[90] br[90] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_93 
+ bl[91] br[91] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_94 
+ bl[92] br[92] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_95 
+ bl[93] br[93] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_96 
+ bl[94] br[94] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_97 
+ bl[95] br[95] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_98 
+ bl[96] br[96] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_99 
+ bl[97] br[97] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_100 
+ bl[98] br[98] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_101 
+ bl[99] br[99] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_102 
+ bl[100] br[100] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_103 
+ bl[101] br[101] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_104 
+ bl[102] br[102] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_105 
+ bl[103] br[103] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_106 
+ bl[104] br[104] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_107 
+ bl[105] br[105] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_108 
+ bl[106] br[106] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_109 
+ bl[107] br[107] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_110 
+ bl[108] br[108] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_111 
+ bl[109] br[109] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_112 
+ bl[110] br[110] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_113 
+ bl[111] br[111] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_114 
+ bl[112] br[112] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_115 
+ bl[113] br[113] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_116 
+ bl[114] br[114] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_117 
+ bl[115] br[115] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_118 
+ bl[116] br[116] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_119 
+ bl[117] br[117] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_120 
+ bl[118] br[118] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_121 
+ bl[119] br[119] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_122 
+ bl[120] br[120] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_123 
+ bl[121] br[121] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_124 
+ bl[122] br[122] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_125 
+ bl[123] br[123] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_126 
+ bl[124] br[124] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_127 
+ bl[125] br[125] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_128 
+ bl[126] br[126] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_129 
+ bl[127] br[127] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_130 
+ bl[128] br[128] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_131 
+ bl[129] br[129] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_132 
+ bl[130] br[130] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_133 
+ bl[131] br[131] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_134 
+ bl[132] br[132] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_135 
+ bl[133] br[133] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_136 
+ bl[134] br[134] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_137 
+ bl[135] br[135] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_138 
+ bl[136] br[136] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_139 
+ bl[137] br[137] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_140 
+ bl[138] br[138] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_141 
+ bl[139] br[139] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_142 
+ bl[140] br[140] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_143 
+ bl[141] br[141] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_144 
+ bl[142] br[142] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_145 
+ bl[143] br[143] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_146 
+ bl[144] br[144] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_147 
+ bl[145] br[145] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_148 
+ bl[146] br[146] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_149 
+ bl[147] br[147] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_150 
+ bl[148] br[148] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_151 
+ bl[149] br[149] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_152 
+ bl[150] br[150] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_153 
+ bl[151] br[151] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_154 
+ bl[152] br[152] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_155 
+ bl[153] br[153] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_156 
+ bl[154] br[154] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_157 
+ bl[155] br[155] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_158 
+ bl[156] br[156] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_159 
+ bl[157] br[157] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_160 
+ bl[158] br[158] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_161 
+ bl[159] br[159] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_162 
+ bl[160] br[160] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_163 
+ bl[161] br[161] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_164 
+ bl[162] br[162] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_165 
+ bl[163] br[163] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_166 
+ bl[164] br[164] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_167 
+ bl[165] br[165] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_168 
+ bl[166] br[166] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_169 
+ bl[167] br[167] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_170 
+ bl[168] br[168] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_171 
+ bl[169] br[169] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_172 
+ bl[170] br[170] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_173 
+ bl[171] br[171] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_174 
+ bl[172] br[172] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_175 
+ bl[173] br[173] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_176 
+ bl[174] br[174] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_177 
+ bl[175] br[175] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_178 
+ bl[176] br[176] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_179 
+ bl[177] br[177] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_180 
+ bl[178] br[178] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_181 
+ bl[179] br[179] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_182 
+ bl[180] br[180] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_183 
+ bl[181] br[181] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_184 
+ bl[182] br[182] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_185 
+ bl[183] br[183] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_186 
+ bl[184] br[184] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_187 
+ bl[185] br[185] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_188 
+ bl[186] br[186] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_189 
+ bl[187] br[187] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_190 
+ bl[188] br[188] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_191 
+ bl[189] br[189] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_192 
+ bl[190] br[190] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_193 
+ bl[191] br[191] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_194 
+ bl[192] br[192] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_195 
+ bl[193] br[193] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_196 
+ bl[194] br[194] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_197 
+ bl[195] br[195] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_198 
+ bl[196] br[196] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_199 
+ bl[197] br[197] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_200 
+ bl[198] br[198] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_201 
+ bl[199] br[199] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_202 
+ bl[200] br[200] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_203 
+ bl[201] br[201] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_204 
+ bl[202] br[202] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_205 
+ bl[203] br[203] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_206 
+ bl[204] br[204] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_207 
+ bl[205] br[205] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_208 
+ bl[206] br[206] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_209 
+ bl[207] br[207] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_210 
+ bl[208] br[208] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_211 
+ bl[209] br[209] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_212 
+ bl[210] br[210] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_213 
+ bl[211] br[211] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_214 
+ bl[212] br[212] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_215 
+ bl[213] br[213] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_216 
+ bl[214] br[214] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_217 
+ bl[215] br[215] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_218 
+ bl[216] br[216] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_219 
+ bl[217] br[217] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_220 
+ bl[218] br[218] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_221 
+ bl[219] br[219] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_222 
+ bl[220] br[220] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_223 
+ bl[221] br[221] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_224 
+ bl[222] br[222] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_225 
+ bl[223] br[223] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_226 
+ bl[224] br[224] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_227 
+ bl[225] br[225] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_228 
+ bl[226] br[226] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_229 
+ bl[227] br[227] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_230 
+ bl[228] br[228] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_231 
+ bl[229] br[229] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_232 
+ bl[230] br[230] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_233 
+ bl[231] br[231] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_234 
+ bl[232] br[232] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_235 
+ bl[233] br[233] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_236 
+ bl[234] br[234] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_237 
+ bl[235] br[235] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_238 
+ bl[236] br[236] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_239 
+ bl[237] br[237] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_240 
+ bl[238] br[238] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_241 
+ bl[239] br[239] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_242 
+ bl[240] br[240] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_243 
+ bl[241] br[241] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_244 
+ bl[242] br[242] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_245 
+ bl[243] br[243] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_246 
+ bl[244] br[244] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_247 
+ bl[245] br[245] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_248 
+ bl[246] br[246] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_249 
+ bl[247] br[247] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_250 
+ bl[248] br[248] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_251 
+ bl[249] br[249] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_252 
+ bl[250] br[250] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_253 
+ bl[251] br[251] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_254 
+ bl[252] br[252] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_255 
+ bl[253] br[253] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_256 
+ bl[254] br[254] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_257 
+ bl[255] br[255] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_258 
+ vdd vdd vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_259 
+ vdd vdd vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_0 
+ vdd vdd vss vdd vpb vnb wl[41] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_43_1 
+ rbl rbr vss vdd vpb vnb wl[41] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_43_2 
+ bl[0] br[0] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_3 
+ bl[1] br[1] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_4 
+ bl[2] br[2] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_5 
+ bl[3] br[3] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_6 
+ bl[4] br[4] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_7 
+ bl[5] br[5] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_8 
+ bl[6] br[6] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_9 
+ bl[7] br[7] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_10 
+ bl[8] br[8] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_11 
+ bl[9] br[9] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_12 
+ bl[10] br[10] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_13 
+ bl[11] br[11] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_14 
+ bl[12] br[12] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_15 
+ bl[13] br[13] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_16 
+ bl[14] br[14] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_17 
+ bl[15] br[15] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_18 
+ bl[16] br[16] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_19 
+ bl[17] br[17] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_20 
+ bl[18] br[18] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_21 
+ bl[19] br[19] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_22 
+ bl[20] br[20] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_23 
+ bl[21] br[21] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_24 
+ bl[22] br[22] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_25 
+ bl[23] br[23] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_26 
+ bl[24] br[24] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_27 
+ bl[25] br[25] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_28 
+ bl[26] br[26] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_29 
+ bl[27] br[27] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_30 
+ bl[28] br[28] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_31 
+ bl[29] br[29] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_32 
+ bl[30] br[30] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_33 
+ bl[31] br[31] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_34 
+ bl[32] br[32] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_35 
+ bl[33] br[33] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_36 
+ bl[34] br[34] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_37 
+ bl[35] br[35] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_38 
+ bl[36] br[36] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_39 
+ bl[37] br[37] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_40 
+ bl[38] br[38] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_41 
+ bl[39] br[39] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_42 
+ bl[40] br[40] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_43 
+ bl[41] br[41] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_44 
+ bl[42] br[42] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_45 
+ bl[43] br[43] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_46 
+ bl[44] br[44] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_47 
+ bl[45] br[45] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_48 
+ bl[46] br[46] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_49 
+ bl[47] br[47] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_50 
+ bl[48] br[48] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_51 
+ bl[49] br[49] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_52 
+ bl[50] br[50] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_53 
+ bl[51] br[51] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_54 
+ bl[52] br[52] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_55 
+ bl[53] br[53] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_56 
+ bl[54] br[54] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_57 
+ bl[55] br[55] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_58 
+ bl[56] br[56] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_59 
+ bl[57] br[57] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_60 
+ bl[58] br[58] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_61 
+ bl[59] br[59] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_62 
+ bl[60] br[60] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_63 
+ bl[61] br[61] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_64 
+ bl[62] br[62] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_65 
+ bl[63] br[63] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_66 
+ bl[64] br[64] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_67 
+ bl[65] br[65] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_68 
+ bl[66] br[66] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_69 
+ bl[67] br[67] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_70 
+ bl[68] br[68] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_71 
+ bl[69] br[69] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_72 
+ bl[70] br[70] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_73 
+ bl[71] br[71] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_74 
+ bl[72] br[72] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_75 
+ bl[73] br[73] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_76 
+ bl[74] br[74] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_77 
+ bl[75] br[75] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_78 
+ bl[76] br[76] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_79 
+ bl[77] br[77] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_80 
+ bl[78] br[78] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_81 
+ bl[79] br[79] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_82 
+ bl[80] br[80] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_83 
+ bl[81] br[81] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_84 
+ bl[82] br[82] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_85 
+ bl[83] br[83] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_86 
+ bl[84] br[84] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_87 
+ bl[85] br[85] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_88 
+ bl[86] br[86] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_89 
+ bl[87] br[87] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_90 
+ bl[88] br[88] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_91 
+ bl[89] br[89] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_92 
+ bl[90] br[90] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_93 
+ bl[91] br[91] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_94 
+ bl[92] br[92] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_95 
+ bl[93] br[93] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_96 
+ bl[94] br[94] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_97 
+ bl[95] br[95] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_98 
+ bl[96] br[96] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_99 
+ bl[97] br[97] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_100 
+ bl[98] br[98] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_101 
+ bl[99] br[99] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_102 
+ bl[100] br[100] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_103 
+ bl[101] br[101] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_104 
+ bl[102] br[102] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_105 
+ bl[103] br[103] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_106 
+ bl[104] br[104] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_107 
+ bl[105] br[105] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_108 
+ bl[106] br[106] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_109 
+ bl[107] br[107] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_110 
+ bl[108] br[108] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_111 
+ bl[109] br[109] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_112 
+ bl[110] br[110] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_113 
+ bl[111] br[111] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_114 
+ bl[112] br[112] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_115 
+ bl[113] br[113] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_116 
+ bl[114] br[114] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_117 
+ bl[115] br[115] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_118 
+ bl[116] br[116] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_119 
+ bl[117] br[117] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_120 
+ bl[118] br[118] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_121 
+ bl[119] br[119] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_122 
+ bl[120] br[120] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_123 
+ bl[121] br[121] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_124 
+ bl[122] br[122] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_125 
+ bl[123] br[123] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_126 
+ bl[124] br[124] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_127 
+ bl[125] br[125] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_128 
+ bl[126] br[126] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_129 
+ bl[127] br[127] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_130 
+ bl[128] br[128] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_131 
+ bl[129] br[129] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_132 
+ bl[130] br[130] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_133 
+ bl[131] br[131] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_134 
+ bl[132] br[132] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_135 
+ bl[133] br[133] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_136 
+ bl[134] br[134] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_137 
+ bl[135] br[135] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_138 
+ bl[136] br[136] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_139 
+ bl[137] br[137] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_140 
+ bl[138] br[138] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_141 
+ bl[139] br[139] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_142 
+ bl[140] br[140] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_143 
+ bl[141] br[141] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_144 
+ bl[142] br[142] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_145 
+ bl[143] br[143] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_146 
+ bl[144] br[144] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_147 
+ bl[145] br[145] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_148 
+ bl[146] br[146] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_149 
+ bl[147] br[147] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_150 
+ bl[148] br[148] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_151 
+ bl[149] br[149] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_152 
+ bl[150] br[150] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_153 
+ bl[151] br[151] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_154 
+ bl[152] br[152] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_155 
+ bl[153] br[153] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_156 
+ bl[154] br[154] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_157 
+ bl[155] br[155] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_158 
+ bl[156] br[156] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_159 
+ bl[157] br[157] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_160 
+ bl[158] br[158] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_161 
+ bl[159] br[159] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_162 
+ bl[160] br[160] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_163 
+ bl[161] br[161] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_164 
+ bl[162] br[162] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_165 
+ bl[163] br[163] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_166 
+ bl[164] br[164] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_167 
+ bl[165] br[165] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_168 
+ bl[166] br[166] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_169 
+ bl[167] br[167] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_170 
+ bl[168] br[168] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_171 
+ bl[169] br[169] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_172 
+ bl[170] br[170] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_173 
+ bl[171] br[171] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_174 
+ bl[172] br[172] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_175 
+ bl[173] br[173] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_176 
+ bl[174] br[174] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_177 
+ bl[175] br[175] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_178 
+ bl[176] br[176] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_179 
+ bl[177] br[177] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_180 
+ bl[178] br[178] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_181 
+ bl[179] br[179] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_182 
+ bl[180] br[180] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_183 
+ bl[181] br[181] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_184 
+ bl[182] br[182] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_185 
+ bl[183] br[183] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_186 
+ bl[184] br[184] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_187 
+ bl[185] br[185] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_188 
+ bl[186] br[186] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_189 
+ bl[187] br[187] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_190 
+ bl[188] br[188] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_191 
+ bl[189] br[189] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_192 
+ bl[190] br[190] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_193 
+ bl[191] br[191] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_194 
+ bl[192] br[192] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_195 
+ bl[193] br[193] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_196 
+ bl[194] br[194] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_197 
+ bl[195] br[195] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_198 
+ bl[196] br[196] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_199 
+ bl[197] br[197] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_200 
+ bl[198] br[198] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_201 
+ bl[199] br[199] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_202 
+ bl[200] br[200] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_203 
+ bl[201] br[201] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_204 
+ bl[202] br[202] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_205 
+ bl[203] br[203] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_206 
+ bl[204] br[204] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_207 
+ bl[205] br[205] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_208 
+ bl[206] br[206] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_209 
+ bl[207] br[207] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_210 
+ bl[208] br[208] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_211 
+ bl[209] br[209] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_212 
+ bl[210] br[210] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_213 
+ bl[211] br[211] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_214 
+ bl[212] br[212] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_215 
+ bl[213] br[213] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_216 
+ bl[214] br[214] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_217 
+ bl[215] br[215] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_218 
+ bl[216] br[216] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_219 
+ bl[217] br[217] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_220 
+ bl[218] br[218] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_221 
+ bl[219] br[219] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_222 
+ bl[220] br[220] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_223 
+ bl[221] br[221] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_224 
+ bl[222] br[222] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_225 
+ bl[223] br[223] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_226 
+ bl[224] br[224] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_227 
+ bl[225] br[225] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_228 
+ bl[226] br[226] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_229 
+ bl[227] br[227] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_230 
+ bl[228] br[228] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_231 
+ bl[229] br[229] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_232 
+ bl[230] br[230] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_233 
+ bl[231] br[231] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_234 
+ bl[232] br[232] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_235 
+ bl[233] br[233] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_236 
+ bl[234] br[234] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_237 
+ bl[235] br[235] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_238 
+ bl[236] br[236] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_239 
+ bl[237] br[237] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_240 
+ bl[238] br[238] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_241 
+ bl[239] br[239] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_242 
+ bl[240] br[240] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_243 
+ bl[241] br[241] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_244 
+ bl[242] br[242] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_245 
+ bl[243] br[243] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_246 
+ bl[244] br[244] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_247 
+ bl[245] br[245] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_248 
+ bl[246] br[246] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_249 
+ bl[247] br[247] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_250 
+ bl[248] br[248] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_251 
+ bl[249] br[249] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_252 
+ bl[250] br[250] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_253 
+ bl[251] br[251] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_254 
+ bl[252] br[252] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_255 
+ bl[253] br[253] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_256 
+ bl[254] br[254] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_257 
+ bl[255] br[255] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_258 
+ vdd vdd vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_259 
+ vdd vdd vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_0 
+ vdd vdd vss vdd vpb vnb wl[42] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_44_1 
+ rbl rbr vss vdd vpb vnb wl[42] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_44_2 
+ bl[0] br[0] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_3 
+ bl[1] br[1] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_4 
+ bl[2] br[2] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_5 
+ bl[3] br[3] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_6 
+ bl[4] br[4] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_7 
+ bl[5] br[5] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_8 
+ bl[6] br[6] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_9 
+ bl[7] br[7] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_10 
+ bl[8] br[8] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_11 
+ bl[9] br[9] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_12 
+ bl[10] br[10] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_13 
+ bl[11] br[11] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_14 
+ bl[12] br[12] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_15 
+ bl[13] br[13] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_16 
+ bl[14] br[14] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_17 
+ bl[15] br[15] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_18 
+ bl[16] br[16] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_19 
+ bl[17] br[17] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_20 
+ bl[18] br[18] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_21 
+ bl[19] br[19] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_22 
+ bl[20] br[20] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_23 
+ bl[21] br[21] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_24 
+ bl[22] br[22] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_25 
+ bl[23] br[23] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_26 
+ bl[24] br[24] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_27 
+ bl[25] br[25] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_28 
+ bl[26] br[26] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_29 
+ bl[27] br[27] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_30 
+ bl[28] br[28] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_31 
+ bl[29] br[29] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_32 
+ bl[30] br[30] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_33 
+ bl[31] br[31] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_34 
+ bl[32] br[32] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_35 
+ bl[33] br[33] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_36 
+ bl[34] br[34] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_37 
+ bl[35] br[35] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_38 
+ bl[36] br[36] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_39 
+ bl[37] br[37] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_40 
+ bl[38] br[38] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_41 
+ bl[39] br[39] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_42 
+ bl[40] br[40] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_43 
+ bl[41] br[41] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_44 
+ bl[42] br[42] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_45 
+ bl[43] br[43] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_46 
+ bl[44] br[44] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_47 
+ bl[45] br[45] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_48 
+ bl[46] br[46] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_49 
+ bl[47] br[47] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_50 
+ bl[48] br[48] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_51 
+ bl[49] br[49] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_52 
+ bl[50] br[50] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_53 
+ bl[51] br[51] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_54 
+ bl[52] br[52] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_55 
+ bl[53] br[53] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_56 
+ bl[54] br[54] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_57 
+ bl[55] br[55] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_58 
+ bl[56] br[56] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_59 
+ bl[57] br[57] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_60 
+ bl[58] br[58] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_61 
+ bl[59] br[59] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_62 
+ bl[60] br[60] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_63 
+ bl[61] br[61] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_64 
+ bl[62] br[62] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_65 
+ bl[63] br[63] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_66 
+ bl[64] br[64] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_67 
+ bl[65] br[65] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_68 
+ bl[66] br[66] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_69 
+ bl[67] br[67] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_70 
+ bl[68] br[68] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_71 
+ bl[69] br[69] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_72 
+ bl[70] br[70] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_73 
+ bl[71] br[71] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_74 
+ bl[72] br[72] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_75 
+ bl[73] br[73] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_76 
+ bl[74] br[74] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_77 
+ bl[75] br[75] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_78 
+ bl[76] br[76] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_79 
+ bl[77] br[77] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_80 
+ bl[78] br[78] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_81 
+ bl[79] br[79] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_82 
+ bl[80] br[80] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_83 
+ bl[81] br[81] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_84 
+ bl[82] br[82] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_85 
+ bl[83] br[83] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_86 
+ bl[84] br[84] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_87 
+ bl[85] br[85] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_88 
+ bl[86] br[86] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_89 
+ bl[87] br[87] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_90 
+ bl[88] br[88] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_91 
+ bl[89] br[89] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_92 
+ bl[90] br[90] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_93 
+ bl[91] br[91] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_94 
+ bl[92] br[92] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_95 
+ bl[93] br[93] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_96 
+ bl[94] br[94] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_97 
+ bl[95] br[95] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_98 
+ bl[96] br[96] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_99 
+ bl[97] br[97] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_100 
+ bl[98] br[98] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_101 
+ bl[99] br[99] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_102 
+ bl[100] br[100] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_103 
+ bl[101] br[101] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_104 
+ bl[102] br[102] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_105 
+ bl[103] br[103] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_106 
+ bl[104] br[104] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_107 
+ bl[105] br[105] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_108 
+ bl[106] br[106] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_109 
+ bl[107] br[107] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_110 
+ bl[108] br[108] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_111 
+ bl[109] br[109] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_112 
+ bl[110] br[110] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_113 
+ bl[111] br[111] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_114 
+ bl[112] br[112] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_115 
+ bl[113] br[113] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_116 
+ bl[114] br[114] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_117 
+ bl[115] br[115] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_118 
+ bl[116] br[116] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_119 
+ bl[117] br[117] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_120 
+ bl[118] br[118] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_121 
+ bl[119] br[119] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_122 
+ bl[120] br[120] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_123 
+ bl[121] br[121] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_124 
+ bl[122] br[122] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_125 
+ bl[123] br[123] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_126 
+ bl[124] br[124] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_127 
+ bl[125] br[125] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_128 
+ bl[126] br[126] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_129 
+ bl[127] br[127] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_130 
+ bl[128] br[128] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_131 
+ bl[129] br[129] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_132 
+ bl[130] br[130] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_133 
+ bl[131] br[131] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_134 
+ bl[132] br[132] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_135 
+ bl[133] br[133] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_136 
+ bl[134] br[134] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_137 
+ bl[135] br[135] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_138 
+ bl[136] br[136] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_139 
+ bl[137] br[137] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_140 
+ bl[138] br[138] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_141 
+ bl[139] br[139] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_142 
+ bl[140] br[140] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_143 
+ bl[141] br[141] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_144 
+ bl[142] br[142] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_145 
+ bl[143] br[143] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_146 
+ bl[144] br[144] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_147 
+ bl[145] br[145] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_148 
+ bl[146] br[146] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_149 
+ bl[147] br[147] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_150 
+ bl[148] br[148] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_151 
+ bl[149] br[149] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_152 
+ bl[150] br[150] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_153 
+ bl[151] br[151] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_154 
+ bl[152] br[152] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_155 
+ bl[153] br[153] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_156 
+ bl[154] br[154] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_157 
+ bl[155] br[155] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_158 
+ bl[156] br[156] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_159 
+ bl[157] br[157] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_160 
+ bl[158] br[158] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_161 
+ bl[159] br[159] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_162 
+ bl[160] br[160] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_163 
+ bl[161] br[161] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_164 
+ bl[162] br[162] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_165 
+ bl[163] br[163] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_166 
+ bl[164] br[164] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_167 
+ bl[165] br[165] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_168 
+ bl[166] br[166] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_169 
+ bl[167] br[167] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_170 
+ bl[168] br[168] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_171 
+ bl[169] br[169] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_172 
+ bl[170] br[170] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_173 
+ bl[171] br[171] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_174 
+ bl[172] br[172] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_175 
+ bl[173] br[173] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_176 
+ bl[174] br[174] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_177 
+ bl[175] br[175] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_178 
+ bl[176] br[176] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_179 
+ bl[177] br[177] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_180 
+ bl[178] br[178] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_181 
+ bl[179] br[179] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_182 
+ bl[180] br[180] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_183 
+ bl[181] br[181] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_184 
+ bl[182] br[182] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_185 
+ bl[183] br[183] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_186 
+ bl[184] br[184] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_187 
+ bl[185] br[185] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_188 
+ bl[186] br[186] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_189 
+ bl[187] br[187] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_190 
+ bl[188] br[188] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_191 
+ bl[189] br[189] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_192 
+ bl[190] br[190] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_193 
+ bl[191] br[191] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_194 
+ bl[192] br[192] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_195 
+ bl[193] br[193] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_196 
+ bl[194] br[194] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_197 
+ bl[195] br[195] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_198 
+ bl[196] br[196] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_199 
+ bl[197] br[197] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_200 
+ bl[198] br[198] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_201 
+ bl[199] br[199] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_202 
+ bl[200] br[200] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_203 
+ bl[201] br[201] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_204 
+ bl[202] br[202] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_205 
+ bl[203] br[203] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_206 
+ bl[204] br[204] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_207 
+ bl[205] br[205] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_208 
+ bl[206] br[206] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_209 
+ bl[207] br[207] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_210 
+ bl[208] br[208] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_211 
+ bl[209] br[209] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_212 
+ bl[210] br[210] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_213 
+ bl[211] br[211] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_214 
+ bl[212] br[212] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_215 
+ bl[213] br[213] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_216 
+ bl[214] br[214] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_217 
+ bl[215] br[215] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_218 
+ bl[216] br[216] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_219 
+ bl[217] br[217] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_220 
+ bl[218] br[218] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_221 
+ bl[219] br[219] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_222 
+ bl[220] br[220] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_223 
+ bl[221] br[221] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_224 
+ bl[222] br[222] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_225 
+ bl[223] br[223] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_226 
+ bl[224] br[224] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_227 
+ bl[225] br[225] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_228 
+ bl[226] br[226] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_229 
+ bl[227] br[227] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_230 
+ bl[228] br[228] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_231 
+ bl[229] br[229] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_232 
+ bl[230] br[230] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_233 
+ bl[231] br[231] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_234 
+ bl[232] br[232] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_235 
+ bl[233] br[233] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_236 
+ bl[234] br[234] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_237 
+ bl[235] br[235] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_238 
+ bl[236] br[236] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_239 
+ bl[237] br[237] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_240 
+ bl[238] br[238] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_241 
+ bl[239] br[239] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_242 
+ bl[240] br[240] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_243 
+ bl[241] br[241] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_244 
+ bl[242] br[242] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_245 
+ bl[243] br[243] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_246 
+ bl[244] br[244] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_247 
+ bl[245] br[245] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_248 
+ bl[246] br[246] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_249 
+ bl[247] br[247] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_250 
+ bl[248] br[248] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_251 
+ bl[249] br[249] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_252 
+ bl[250] br[250] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_253 
+ bl[251] br[251] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_254 
+ bl[252] br[252] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_255 
+ bl[253] br[253] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_256 
+ bl[254] br[254] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_257 
+ bl[255] br[255] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_258 
+ vdd vdd vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_259 
+ vdd vdd vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_0 
+ vdd vdd vss vdd vpb vnb wl[43] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_45_1 
+ rbl rbr vss vdd vpb vnb wl[43] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_45_2 
+ bl[0] br[0] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_3 
+ bl[1] br[1] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_4 
+ bl[2] br[2] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_5 
+ bl[3] br[3] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_6 
+ bl[4] br[4] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_7 
+ bl[5] br[5] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_8 
+ bl[6] br[6] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_9 
+ bl[7] br[7] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_10 
+ bl[8] br[8] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_11 
+ bl[9] br[9] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_12 
+ bl[10] br[10] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_13 
+ bl[11] br[11] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_14 
+ bl[12] br[12] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_15 
+ bl[13] br[13] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_16 
+ bl[14] br[14] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_17 
+ bl[15] br[15] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_18 
+ bl[16] br[16] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_19 
+ bl[17] br[17] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_20 
+ bl[18] br[18] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_21 
+ bl[19] br[19] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_22 
+ bl[20] br[20] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_23 
+ bl[21] br[21] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_24 
+ bl[22] br[22] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_25 
+ bl[23] br[23] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_26 
+ bl[24] br[24] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_27 
+ bl[25] br[25] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_28 
+ bl[26] br[26] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_29 
+ bl[27] br[27] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_30 
+ bl[28] br[28] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_31 
+ bl[29] br[29] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_32 
+ bl[30] br[30] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_33 
+ bl[31] br[31] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_34 
+ bl[32] br[32] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_35 
+ bl[33] br[33] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_36 
+ bl[34] br[34] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_37 
+ bl[35] br[35] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_38 
+ bl[36] br[36] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_39 
+ bl[37] br[37] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_40 
+ bl[38] br[38] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_41 
+ bl[39] br[39] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_42 
+ bl[40] br[40] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_43 
+ bl[41] br[41] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_44 
+ bl[42] br[42] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_45 
+ bl[43] br[43] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_46 
+ bl[44] br[44] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_47 
+ bl[45] br[45] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_48 
+ bl[46] br[46] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_49 
+ bl[47] br[47] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_50 
+ bl[48] br[48] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_51 
+ bl[49] br[49] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_52 
+ bl[50] br[50] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_53 
+ bl[51] br[51] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_54 
+ bl[52] br[52] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_55 
+ bl[53] br[53] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_56 
+ bl[54] br[54] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_57 
+ bl[55] br[55] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_58 
+ bl[56] br[56] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_59 
+ bl[57] br[57] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_60 
+ bl[58] br[58] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_61 
+ bl[59] br[59] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_62 
+ bl[60] br[60] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_63 
+ bl[61] br[61] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_64 
+ bl[62] br[62] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_65 
+ bl[63] br[63] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_66 
+ bl[64] br[64] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_67 
+ bl[65] br[65] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_68 
+ bl[66] br[66] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_69 
+ bl[67] br[67] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_70 
+ bl[68] br[68] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_71 
+ bl[69] br[69] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_72 
+ bl[70] br[70] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_73 
+ bl[71] br[71] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_74 
+ bl[72] br[72] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_75 
+ bl[73] br[73] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_76 
+ bl[74] br[74] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_77 
+ bl[75] br[75] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_78 
+ bl[76] br[76] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_79 
+ bl[77] br[77] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_80 
+ bl[78] br[78] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_81 
+ bl[79] br[79] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_82 
+ bl[80] br[80] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_83 
+ bl[81] br[81] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_84 
+ bl[82] br[82] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_85 
+ bl[83] br[83] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_86 
+ bl[84] br[84] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_87 
+ bl[85] br[85] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_88 
+ bl[86] br[86] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_89 
+ bl[87] br[87] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_90 
+ bl[88] br[88] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_91 
+ bl[89] br[89] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_92 
+ bl[90] br[90] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_93 
+ bl[91] br[91] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_94 
+ bl[92] br[92] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_95 
+ bl[93] br[93] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_96 
+ bl[94] br[94] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_97 
+ bl[95] br[95] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_98 
+ bl[96] br[96] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_99 
+ bl[97] br[97] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_100 
+ bl[98] br[98] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_101 
+ bl[99] br[99] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_102 
+ bl[100] br[100] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_103 
+ bl[101] br[101] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_104 
+ bl[102] br[102] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_105 
+ bl[103] br[103] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_106 
+ bl[104] br[104] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_107 
+ bl[105] br[105] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_108 
+ bl[106] br[106] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_109 
+ bl[107] br[107] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_110 
+ bl[108] br[108] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_111 
+ bl[109] br[109] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_112 
+ bl[110] br[110] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_113 
+ bl[111] br[111] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_114 
+ bl[112] br[112] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_115 
+ bl[113] br[113] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_116 
+ bl[114] br[114] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_117 
+ bl[115] br[115] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_118 
+ bl[116] br[116] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_119 
+ bl[117] br[117] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_120 
+ bl[118] br[118] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_121 
+ bl[119] br[119] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_122 
+ bl[120] br[120] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_123 
+ bl[121] br[121] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_124 
+ bl[122] br[122] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_125 
+ bl[123] br[123] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_126 
+ bl[124] br[124] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_127 
+ bl[125] br[125] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_128 
+ bl[126] br[126] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_129 
+ bl[127] br[127] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_130 
+ bl[128] br[128] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_131 
+ bl[129] br[129] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_132 
+ bl[130] br[130] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_133 
+ bl[131] br[131] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_134 
+ bl[132] br[132] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_135 
+ bl[133] br[133] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_136 
+ bl[134] br[134] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_137 
+ bl[135] br[135] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_138 
+ bl[136] br[136] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_139 
+ bl[137] br[137] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_140 
+ bl[138] br[138] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_141 
+ bl[139] br[139] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_142 
+ bl[140] br[140] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_143 
+ bl[141] br[141] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_144 
+ bl[142] br[142] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_145 
+ bl[143] br[143] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_146 
+ bl[144] br[144] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_147 
+ bl[145] br[145] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_148 
+ bl[146] br[146] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_149 
+ bl[147] br[147] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_150 
+ bl[148] br[148] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_151 
+ bl[149] br[149] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_152 
+ bl[150] br[150] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_153 
+ bl[151] br[151] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_154 
+ bl[152] br[152] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_155 
+ bl[153] br[153] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_156 
+ bl[154] br[154] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_157 
+ bl[155] br[155] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_158 
+ bl[156] br[156] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_159 
+ bl[157] br[157] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_160 
+ bl[158] br[158] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_161 
+ bl[159] br[159] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_162 
+ bl[160] br[160] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_163 
+ bl[161] br[161] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_164 
+ bl[162] br[162] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_165 
+ bl[163] br[163] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_166 
+ bl[164] br[164] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_167 
+ bl[165] br[165] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_168 
+ bl[166] br[166] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_169 
+ bl[167] br[167] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_170 
+ bl[168] br[168] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_171 
+ bl[169] br[169] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_172 
+ bl[170] br[170] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_173 
+ bl[171] br[171] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_174 
+ bl[172] br[172] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_175 
+ bl[173] br[173] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_176 
+ bl[174] br[174] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_177 
+ bl[175] br[175] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_178 
+ bl[176] br[176] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_179 
+ bl[177] br[177] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_180 
+ bl[178] br[178] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_181 
+ bl[179] br[179] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_182 
+ bl[180] br[180] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_183 
+ bl[181] br[181] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_184 
+ bl[182] br[182] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_185 
+ bl[183] br[183] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_186 
+ bl[184] br[184] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_187 
+ bl[185] br[185] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_188 
+ bl[186] br[186] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_189 
+ bl[187] br[187] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_190 
+ bl[188] br[188] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_191 
+ bl[189] br[189] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_192 
+ bl[190] br[190] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_193 
+ bl[191] br[191] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_194 
+ bl[192] br[192] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_195 
+ bl[193] br[193] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_196 
+ bl[194] br[194] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_197 
+ bl[195] br[195] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_198 
+ bl[196] br[196] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_199 
+ bl[197] br[197] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_200 
+ bl[198] br[198] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_201 
+ bl[199] br[199] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_202 
+ bl[200] br[200] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_203 
+ bl[201] br[201] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_204 
+ bl[202] br[202] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_205 
+ bl[203] br[203] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_206 
+ bl[204] br[204] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_207 
+ bl[205] br[205] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_208 
+ bl[206] br[206] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_209 
+ bl[207] br[207] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_210 
+ bl[208] br[208] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_211 
+ bl[209] br[209] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_212 
+ bl[210] br[210] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_213 
+ bl[211] br[211] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_214 
+ bl[212] br[212] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_215 
+ bl[213] br[213] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_216 
+ bl[214] br[214] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_217 
+ bl[215] br[215] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_218 
+ bl[216] br[216] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_219 
+ bl[217] br[217] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_220 
+ bl[218] br[218] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_221 
+ bl[219] br[219] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_222 
+ bl[220] br[220] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_223 
+ bl[221] br[221] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_224 
+ bl[222] br[222] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_225 
+ bl[223] br[223] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_226 
+ bl[224] br[224] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_227 
+ bl[225] br[225] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_228 
+ bl[226] br[226] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_229 
+ bl[227] br[227] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_230 
+ bl[228] br[228] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_231 
+ bl[229] br[229] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_232 
+ bl[230] br[230] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_233 
+ bl[231] br[231] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_234 
+ bl[232] br[232] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_235 
+ bl[233] br[233] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_236 
+ bl[234] br[234] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_237 
+ bl[235] br[235] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_238 
+ bl[236] br[236] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_239 
+ bl[237] br[237] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_240 
+ bl[238] br[238] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_241 
+ bl[239] br[239] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_242 
+ bl[240] br[240] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_243 
+ bl[241] br[241] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_244 
+ bl[242] br[242] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_245 
+ bl[243] br[243] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_246 
+ bl[244] br[244] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_247 
+ bl[245] br[245] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_248 
+ bl[246] br[246] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_249 
+ bl[247] br[247] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_250 
+ bl[248] br[248] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_251 
+ bl[249] br[249] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_252 
+ bl[250] br[250] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_253 
+ bl[251] br[251] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_254 
+ bl[252] br[252] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_255 
+ bl[253] br[253] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_256 
+ bl[254] br[254] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_257 
+ bl[255] br[255] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_258 
+ vdd vdd vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_259 
+ vdd vdd vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_0 
+ vdd vdd vss vdd vpb vnb wl[44] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_46_1 
+ rbl rbr vss vdd vpb vnb wl[44] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_46_2 
+ bl[0] br[0] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_3 
+ bl[1] br[1] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_4 
+ bl[2] br[2] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_5 
+ bl[3] br[3] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_6 
+ bl[4] br[4] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_7 
+ bl[5] br[5] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_8 
+ bl[6] br[6] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_9 
+ bl[7] br[7] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_10 
+ bl[8] br[8] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_11 
+ bl[9] br[9] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_12 
+ bl[10] br[10] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_13 
+ bl[11] br[11] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_14 
+ bl[12] br[12] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_15 
+ bl[13] br[13] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_16 
+ bl[14] br[14] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_17 
+ bl[15] br[15] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_18 
+ bl[16] br[16] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_19 
+ bl[17] br[17] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_20 
+ bl[18] br[18] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_21 
+ bl[19] br[19] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_22 
+ bl[20] br[20] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_23 
+ bl[21] br[21] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_24 
+ bl[22] br[22] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_25 
+ bl[23] br[23] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_26 
+ bl[24] br[24] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_27 
+ bl[25] br[25] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_28 
+ bl[26] br[26] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_29 
+ bl[27] br[27] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_30 
+ bl[28] br[28] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_31 
+ bl[29] br[29] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_32 
+ bl[30] br[30] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_33 
+ bl[31] br[31] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_34 
+ bl[32] br[32] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_35 
+ bl[33] br[33] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_36 
+ bl[34] br[34] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_37 
+ bl[35] br[35] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_38 
+ bl[36] br[36] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_39 
+ bl[37] br[37] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_40 
+ bl[38] br[38] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_41 
+ bl[39] br[39] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_42 
+ bl[40] br[40] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_43 
+ bl[41] br[41] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_44 
+ bl[42] br[42] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_45 
+ bl[43] br[43] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_46 
+ bl[44] br[44] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_47 
+ bl[45] br[45] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_48 
+ bl[46] br[46] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_49 
+ bl[47] br[47] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_50 
+ bl[48] br[48] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_51 
+ bl[49] br[49] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_52 
+ bl[50] br[50] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_53 
+ bl[51] br[51] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_54 
+ bl[52] br[52] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_55 
+ bl[53] br[53] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_56 
+ bl[54] br[54] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_57 
+ bl[55] br[55] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_58 
+ bl[56] br[56] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_59 
+ bl[57] br[57] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_60 
+ bl[58] br[58] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_61 
+ bl[59] br[59] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_62 
+ bl[60] br[60] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_63 
+ bl[61] br[61] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_64 
+ bl[62] br[62] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_65 
+ bl[63] br[63] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_66 
+ bl[64] br[64] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_67 
+ bl[65] br[65] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_68 
+ bl[66] br[66] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_69 
+ bl[67] br[67] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_70 
+ bl[68] br[68] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_71 
+ bl[69] br[69] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_72 
+ bl[70] br[70] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_73 
+ bl[71] br[71] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_74 
+ bl[72] br[72] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_75 
+ bl[73] br[73] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_76 
+ bl[74] br[74] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_77 
+ bl[75] br[75] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_78 
+ bl[76] br[76] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_79 
+ bl[77] br[77] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_80 
+ bl[78] br[78] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_81 
+ bl[79] br[79] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_82 
+ bl[80] br[80] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_83 
+ bl[81] br[81] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_84 
+ bl[82] br[82] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_85 
+ bl[83] br[83] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_86 
+ bl[84] br[84] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_87 
+ bl[85] br[85] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_88 
+ bl[86] br[86] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_89 
+ bl[87] br[87] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_90 
+ bl[88] br[88] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_91 
+ bl[89] br[89] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_92 
+ bl[90] br[90] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_93 
+ bl[91] br[91] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_94 
+ bl[92] br[92] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_95 
+ bl[93] br[93] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_96 
+ bl[94] br[94] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_97 
+ bl[95] br[95] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_98 
+ bl[96] br[96] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_99 
+ bl[97] br[97] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_100 
+ bl[98] br[98] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_101 
+ bl[99] br[99] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_102 
+ bl[100] br[100] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_103 
+ bl[101] br[101] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_104 
+ bl[102] br[102] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_105 
+ bl[103] br[103] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_106 
+ bl[104] br[104] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_107 
+ bl[105] br[105] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_108 
+ bl[106] br[106] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_109 
+ bl[107] br[107] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_110 
+ bl[108] br[108] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_111 
+ bl[109] br[109] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_112 
+ bl[110] br[110] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_113 
+ bl[111] br[111] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_114 
+ bl[112] br[112] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_115 
+ bl[113] br[113] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_116 
+ bl[114] br[114] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_117 
+ bl[115] br[115] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_118 
+ bl[116] br[116] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_119 
+ bl[117] br[117] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_120 
+ bl[118] br[118] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_121 
+ bl[119] br[119] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_122 
+ bl[120] br[120] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_123 
+ bl[121] br[121] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_124 
+ bl[122] br[122] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_125 
+ bl[123] br[123] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_126 
+ bl[124] br[124] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_127 
+ bl[125] br[125] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_128 
+ bl[126] br[126] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_129 
+ bl[127] br[127] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_130 
+ bl[128] br[128] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_131 
+ bl[129] br[129] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_132 
+ bl[130] br[130] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_133 
+ bl[131] br[131] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_134 
+ bl[132] br[132] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_135 
+ bl[133] br[133] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_136 
+ bl[134] br[134] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_137 
+ bl[135] br[135] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_138 
+ bl[136] br[136] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_139 
+ bl[137] br[137] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_140 
+ bl[138] br[138] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_141 
+ bl[139] br[139] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_142 
+ bl[140] br[140] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_143 
+ bl[141] br[141] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_144 
+ bl[142] br[142] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_145 
+ bl[143] br[143] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_146 
+ bl[144] br[144] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_147 
+ bl[145] br[145] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_148 
+ bl[146] br[146] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_149 
+ bl[147] br[147] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_150 
+ bl[148] br[148] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_151 
+ bl[149] br[149] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_152 
+ bl[150] br[150] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_153 
+ bl[151] br[151] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_154 
+ bl[152] br[152] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_155 
+ bl[153] br[153] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_156 
+ bl[154] br[154] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_157 
+ bl[155] br[155] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_158 
+ bl[156] br[156] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_159 
+ bl[157] br[157] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_160 
+ bl[158] br[158] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_161 
+ bl[159] br[159] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_162 
+ bl[160] br[160] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_163 
+ bl[161] br[161] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_164 
+ bl[162] br[162] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_165 
+ bl[163] br[163] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_166 
+ bl[164] br[164] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_167 
+ bl[165] br[165] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_168 
+ bl[166] br[166] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_169 
+ bl[167] br[167] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_170 
+ bl[168] br[168] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_171 
+ bl[169] br[169] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_172 
+ bl[170] br[170] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_173 
+ bl[171] br[171] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_174 
+ bl[172] br[172] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_175 
+ bl[173] br[173] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_176 
+ bl[174] br[174] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_177 
+ bl[175] br[175] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_178 
+ bl[176] br[176] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_179 
+ bl[177] br[177] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_180 
+ bl[178] br[178] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_181 
+ bl[179] br[179] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_182 
+ bl[180] br[180] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_183 
+ bl[181] br[181] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_184 
+ bl[182] br[182] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_185 
+ bl[183] br[183] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_186 
+ bl[184] br[184] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_187 
+ bl[185] br[185] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_188 
+ bl[186] br[186] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_189 
+ bl[187] br[187] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_190 
+ bl[188] br[188] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_191 
+ bl[189] br[189] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_192 
+ bl[190] br[190] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_193 
+ bl[191] br[191] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_194 
+ bl[192] br[192] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_195 
+ bl[193] br[193] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_196 
+ bl[194] br[194] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_197 
+ bl[195] br[195] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_198 
+ bl[196] br[196] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_199 
+ bl[197] br[197] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_200 
+ bl[198] br[198] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_201 
+ bl[199] br[199] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_202 
+ bl[200] br[200] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_203 
+ bl[201] br[201] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_204 
+ bl[202] br[202] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_205 
+ bl[203] br[203] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_206 
+ bl[204] br[204] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_207 
+ bl[205] br[205] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_208 
+ bl[206] br[206] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_209 
+ bl[207] br[207] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_210 
+ bl[208] br[208] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_211 
+ bl[209] br[209] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_212 
+ bl[210] br[210] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_213 
+ bl[211] br[211] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_214 
+ bl[212] br[212] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_215 
+ bl[213] br[213] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_216 
+ bl[214] br[214] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_217 
+ bl[215] br[215] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_218 
+ bl[216] br[216] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_219 
+ bl[217] br[217] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_220 
+ bl[218] br[218] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_221 
+ bl[219] br[219] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_222 
+ bl[220] br[220] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_223 
+ bl[221] br[221] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_224 
+ bl[222] br[222] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_225 
+ bl[223] br[223] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_226 
+ bl[224] br[224] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_227 
+ bl[225] br[225] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_228 
+ bl[226] br[226] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_229 
+ bl[227] br[227] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_230 
+ bl[228] br[228] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_231 
+ bl[229] br[229] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_232 
+ bl[230] br[230] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_233 
+ bl[231] br[231] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_234 
+ bl[232] br[232] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_235 
+ bl[233] br[233] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_236 
+ bl[234] br[234] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_237 
+ bl[235] br[235] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_238 
+ bl[236] br[236] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_239 
+ bl[237] br[237] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_240 
+ bl[238] br[238] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_241 
+ bl[239] br[239] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_242 
+ bl[240] br[240] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_243 
+ bl[241] br[241] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_244 
+ bl[242] br[242] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_245 
+ bl[243] br[243] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_246 
+ bl[244] br[244] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_247 
+ bl[245] br[245] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_248 
+ bl[246] br[246] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_249 
+ bl[247] br[247] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_250 
+ bl[248] br[248] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_251 
+ bl[249] br[249] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_252 
+ bl[250] br[250] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_253 
+ bl[251] br[251] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_254 
+ bl[252] br[252] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_255 
+ bl[253] br[253] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_256 
+ bl[254] br[254] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_257 
+ bl[255] br[255] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_258 
+ vdd vdd vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_259 
+ vdd vdd vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_0 
+ vdd vdd vss vdd vpb vnb wl[45] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_47_1 
+ rbl rbr vss vdd vpb vnb wl[45] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_47_2 
+ bl[0] br[0] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_3 
+ bl[1] br[1] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_4 
+ bl[2] br[2] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_5 
+ bl[3] br[3] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_6 
+ bl[4] br[4] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_7 
+ bl[5] br[5] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_8 
+ bl[6] br[6] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_9 
+ bl[7] br[7] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_10 
+ bl[8] br[8] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_11 
+ bl[9] br[9] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_12 
+ bl[10] br[10] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_13 
+ bl[11] br[11] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_14 
+ bl[12] br[12] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_15 
+ bl[13] br[13] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_16 
+ bl[14] br[14] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_17 
+ bl[15] br[15] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_18 
+ bl[16] br[16] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_19 
+ bl[17] br[17] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_20 
+ bl[18] br[18] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_21 
+ bl[19] br[19] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_22 
+ bl[20] br[20] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_23 
+ bl[21] br[21] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_24 
+ bl[22] br[22] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_25 
+ bl[23] br[23] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_26 
+ bl[24] br[24] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_27 
+ bl[25] br[25] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_28 
+ bl[26] br[26] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_29 
+ bl[27] br[27] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_30 
+ bl[28] br[28] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_31 
+ bl[29] br[29] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_32 
+ bl[30] br[30] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_33 
+ bl[31] br[31] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_34 
+ bl[32] br[32] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_35 
+ bl[33] br[33] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_36 
+ bl[34] br[34] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_37 
+ bl[35] br[35] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_38 
+ bl[36] br[36] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_39 
+ bl[37] br[37] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_40 
+ bl[38] br[38] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_41 
+ bl[39] br[39] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_42 
+ bl[40] br[40] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_43 
+ bl[41] br[41] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_44 
+ bl[42] br[42] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_45 
+ bl[43] br[43] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_46 
+ bl[44] br[44] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_47 
+ bl[45] br[45] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_48 
+ bl[46] br[46] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_49 
+ bl[47] br[47] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_50 
+ bl[48] br[48] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_51 
+ bl[49] br[49] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_52 
+ bl[50] br[50] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_53 
+ bl[51] br[51] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_54 
+ bl[52] br[52] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_55 
+ bl[53] br[53] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_56 
+ bl[54] br[54] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_57 
+ bl[55] br[55] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_58 
+ bl[56] br[56] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_59 
+ bl[57] br[57] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_60 
+ bl[58] br[58] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_61 
+ bl[59] br[59] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_62 
+ bl[60] br[60] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_63 
+ bl[61] br[61] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_64 
+ bl[62] br[62] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_65 
+ bl[63] br[63] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_66 
+ bl[64] br[64] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_67 
+ bl[65] br[65] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_68 
+ bl[66] br[66] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_69 
+ bl[67] br[67] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_70 
+ bl[68] br[68] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_71 
+ bl[69] br[69] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_72 
+ bl[70] br[70] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_73 
+ bl[71] br[71] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_74 
+ bl[72] br[72] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_75 
+ bl[73] br[73] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_76 
+ bl[74] br[74] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_77 
+ bl[75] br[75] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_78 
+ bl[76] br[76] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_79 
+ bl[77] br[77] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_80 
+ bl[78] br[78] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_81 
+ bl[79] br[79] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_82 
+ bl[80] br[80] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_83 
+ bl[81] br[81] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_84 
+ bl[82] br[82] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_85 
+ bl[83] br[83] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_86 
+ bl[84] br[84] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_87 
+ bl[85] br[85] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_88 
+ bl[86] br[86] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_89 
+ bl[87] br[87] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_90 
+ bl[88] br[88] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_91 
+ bl[89] br[89] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_92 
+ bl[90] br[90] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_93 
+ bl[91] br[91] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_94 
+ bl[92] br[92] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_95 
+ bl[93] br[93] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_96 
+ bl[94] br[94] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_97 
+ bl[95] br[95] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_98 
+ bl[96] br[96] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_99 
+ bl[97] br[97] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_100 
+ bl[98] br[98] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_101 
+ bl[99] br[99] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_102 
+ bl[100] br[100] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_103 
+ bl[101] br[101] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_104 
+ bl[102] br[102] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_105 
+ bl[103] br[103] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_106 
+ bl[104] br[104] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_107 
+ bl[105] br[105] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_108 
+ bl[106] br[106] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_109 
+ bl[107] br[107] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_110 
+ bl[108] br[108] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_111 
+ bl[109] br[109] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_112 
+ bl[110] br[110] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_113 
+ bl[111] br[111] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_114 
+ bl[112] br[112] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_115 
+ bl[113] br[113] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_116 
+ bl[114] br[114] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_117 
+ bl[115] br[115] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_118 
+ bl[116] br[116] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_119 
+ bl[117] br[117] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_120 
+ bl[118] br[118] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_121 
+ bl[119] br[119] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_122 
+ bl[120] br[120] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_123 
+ bl[121] br[121] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_124 
+ bl[122] br[122] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_125 
+ bl[123] br[123] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_126 
+ bl[124] br[124] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_127 
+ bl[125] br[125] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_128 
+ bl[126] br[126] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_129 
+ bl[127] br[127] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_130 
+ bl[128] br[128] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_131 
+ bl[129] br[129] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_132 
+ bl[130] br[130] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_133 
+ bl[131] br[131] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_134 
+ bl[132] br[132] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_135 
+ bl[133] br[133] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_136 
+ bl[134] br[134] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_137 
+ bl[135] br[135] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_138 
+ bl[136] br[136] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_139 
+ bl[137] br[137] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_140 
+ bl[138] br[138] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_141 
+ bl[139] br[139] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_142 
+ bl[140] br[140] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_143 
+ bl[141] br[141] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_144 
+ bl[142] br[142] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_145 
+ bl[143] br[143] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_146 
+ bl[144] br[144] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_147 
+ bl[145] br[145] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_148 
+ bl[146] br[146] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_149 
+ bl[147] br[147] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_150 
+ bl[148] br[148] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_151 
+ bl[149] br[149] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_152 
+ bl[150] br[150] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_153 
+ bl[151] br[151] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_154 
+ bl[152] br[152] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_155 
+ bl[153] br[153] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_156 
+ bl[154] br[154] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_157 
+ bl[155] br[155] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_158 
+ bl[156] br[156] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_159 
+ bl[157] br[157] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_160 
+ bl[158] br[158] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_161 
+ bl[159] br[159] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_162 
+ bl[160] br[160] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_163 
+ bl[161] br[161] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_164 
+ bl[162] br[162] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_165 
+ bl[163] br[163] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_166 
+ bl[164] br[164] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_167 
+ bl[165] br[165] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_168 
+ bl[166] br[166] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_169 
+ bl[167] br[167] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_170 
+ bl[168] br[168] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_171 
+ bl[169] br[169] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_172 
+ bl[170] br[170] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_173 
+ bl[171] br[171] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_174 
+ bl[172] br[172] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_175 
+ bl[173] br[173] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_176 
+ bl[174] br[174] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_177 
+ bl[175] br[175] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_178 
+ bl[176] br[176] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_179 
+ bl[177] br[177] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_180 
+ bl[178] br[178] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_181 
+ bl[179] br[179] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_182 
+ bl[180] br[180] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_183 
+ bl[181] br[181] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_184 
+ bl[182] br[182] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_185 
+ bl[183] br[183] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_186 
+ bl[184] br[184] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_187 
+ bl[185] br[185] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_188 
+ bl[186] br[186] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_189 
+ bl[187] br[187] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_190 
+ bl[188] br[188] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_191 
+ bl[189] br[189] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_192 
+ bl[190] br[190] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_193 
+ bl[191] br[191] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_194 
+ bl[192] br[192] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_195 
+ bl[193] br[193] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_196 
+ bl[194] br[194] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_197 
+ bl[195] br[195] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_198 
+ bl[196] br[196] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_199 
+ bl[197] br[197] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_200 
+ bl[198] br[198] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_201 
+ bl[199] br[199] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_202 
+ bl[200] br[200] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_203 
+ bl[201] br[201] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_204 
+ bl[202] br[202] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_205 
+ bl[203] br[203] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_206 
+ bl[204] br[204] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_207 
+ bl[205] br[205] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_208 
+ bl[206] br[206] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_209 
+ bl[207] br[207] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_210 
+ bl[208] br[208] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_211 
+ bl[209] br[209] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_212 
+ bl[210] br[210] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_213 
+ bl[211] br[211] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_214 
+ bl[212] br[212] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_215 
+ bl[213] br[213] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_216 
+ bl[214] br[214] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_217 
+ bl[215] br[215] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_218 
+ bl[216] br[216] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_219 
+ bl[217] br[217] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_220 
+ bl[218] br[218] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_221 
+ bl[219] br[219] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_222 
+ bl[220] br[220] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_223 
+ bl[221] br[221] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_224 
+ bl[222] br[222] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_225 
+ bl[223] br[223] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_226 
+ bl[224] br[224] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_227 
+ bl[225] br[225] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_228 
+ bl[226] br[226] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_229 
+ bl[227] br[227] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_230 
+ bl[228] br[228] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_231 
+ bl[229] br[229] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_232 
+ bl[230] br[230] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_233 
+ bl[231] br[231] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_234 
+ bl[232] br[232] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_235 
+ bl[233] br[233] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_236 
+ bl[234] br[234] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_237 
+ bl[235] br[235] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_238 
+ bl[236] br[236] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_239 
+ bl[237] br[237] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_240 
+ bl[238] br[238] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_241 
+ bl[239] br[239] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_242 
+ bl[240] br[240] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_243 
+ bl[241] br[241] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_244 
+ bl[242] br[242] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_245 
+ bl[243] br[243] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_246 
+ bl[244] br[244] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_247 
+ bl[245] br[245] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_248 
+ bl[246] br[246] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_249 
+ bl[247] br[247] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_250 
+ bl[248] br[248] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_251 
+ bl[249] br[249] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_252 
+ bl[250] br[250] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_253 
+ bl[251] br[251] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_254 
+ bl[252] br[252] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_255 
+ bl[253] br[253] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_256 
+ bl[254] br[254] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_257 
+ bl[255] br[255] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_258 
+ vdd vdd vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_259 
+ vdd vdd vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_0 
+ vdd vdd vss vdd vpb vnb wl[46] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_48_1 
+ rbl rbr vss vdd vpb vnb wl[46] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_48_2 
+ bl[0] br[0] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_3 
+ bl[1] br[1] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_4 
+ bl[2] br[2] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_5 
+ bl[3] br[3] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_6 
+ bl[4] br[4] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_7 
+ bl[5] br[5] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_8 
+ bl[6] br[6] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_9 
+ bl[7] br[7] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_10 
+ bl[8] br[8] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_11 
+ bl[9] br[9] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_12 
+ bl[10] br[10] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_13 
+ bl[11] br[11] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_14 
+ bl[12] br[12] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_15 
+ bl[13] br[13] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_16 
+ bl[14] br[14] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_17 
+ bl[15] br[15] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_18 
+ bl[16] br[16] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_19 
+ bl[17] br[17] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_20 
+ bl[18] br[18] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_21 
+ bl[19] br[19] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_22 
+ bl[20] br[20] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_23 
+ bl[21] br[21] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_24 
+ bl[22] br[22] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_25 
+ bl[23] br[23] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_26 
+ bl[24] br[24] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_27 
+ bl[25] br[25] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_28 
+ bl[26] br[26] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_29 
+ bl[27] br[27] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_30 
+ bl[28] br[28] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_31 
+ bl[29] br[29] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_32 
+ bl[30] br[30] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_33 
+ bl[31] br[31] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_34 
+ bl[32] br[32] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_35 
+ bl[33] br[33] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_36 
+ bl[34] br[34] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_37 
+ bl[35] br[35] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_38 
+ bl[36] br[36] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_39 
+ bl[37] br[37] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_40 
+ bl[38] br[38] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_41 
+ bl[39] br[39] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_42 
+ bl[40] br[40] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_43 
+ bl[41] br[41] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_44 
+ bl[42] br[42] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_45 
+ bl[43] br[43] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_46 
+ bl[44] br[44] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_47 
+ bl[45] br[45] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_48 
+ bl[46] br[46] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_49 
+ bl[47] br[47] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_50 
+ bl[48] br[48] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_51 
+ bl[49] br[49] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_52 
+ bl[50] br[50] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_53 
+ bl[51] br[51] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_54 
+ bl[52] br[52] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_55 
+ bl[53] br[53] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_56 
+ bl[54] br[54] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_57 
+ bl[55] br[55] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_58 
+ bl[56] br[56] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_59 
+ bl[57] br[57] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_60 
+ bl[58] br[58] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_61 
+ bl[59] br[59] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_62 
+ bl[60] br[60] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_63 
+ bl[61] br[61] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_64 
+ bl[62] br[62] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_65 
+ bl[63] br[63] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_66 
+ bl[64] br[64] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_67 
+ bl[65] br[65] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_68 
+ bl[66] br[66] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_69 
+ bl[67] br[67] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_70 
+ bl[68] br[68] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_71 
+ bl[69] br[69] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_72 
+ bl[70] br[70] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_73 
+ bl[71] br[71] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_74 
+ bl[72] br[72] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_75 
+ bl[73] br[73] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_76 
+ bl[74] br[74] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_77 
+ bl[75] br[75] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_78 
+ bl[76] br[76] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_79 
+ bl[77] br[77] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_80 
+ bl[78] br[78] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_81 
+ bl[79] br[79] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_82 
+ bl[80] br[80] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_83 
+ bl[81] br[81] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_84 
+ bl[82] br[82] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_85 
+ bl[83] br[83] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_86 
+ bl[84] br[84] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_87 
+ bl[85] br[85] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_88 
+ bl[86] br[86] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_89 
+ bl[87] br[87] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_90 
+ bl[88] br[88] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_91 
+ bl[89] br[89] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_92 
+ bl[90] br[90] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_93 
+ bl[91] br[91] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_94 
+ bl[92] br[92] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_95 
+ bl[93] br[93] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_96 
+ bl[94] br[94] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_97 
+ bl[95] br[95] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_98 
+ bl[96] br[96] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_99 
+ bl[97] br[97] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_100 
+ bl[98] br[98] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_101 
+ bl[99] br[99] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_102 
+ bl[100] br[100] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_103 
+ bl[101] br[101] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_104 
+ bl[102] br[102] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_105 
+ bl[103] br[103] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_106 
+ bl[104] br[104] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_107 
+ bl[105] br[105] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_108 
+ bl[106] br[106] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_109 
+ bl[107] br[107] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_110 
+ bl[108] br[108] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_111 
+ bl[109] br[109] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_112 
+ bl[110] br[110] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_113 
+ bl[111] br[111] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_114 
+ bl[112] br[112] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_115 
+ bl[113] br[113] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_116 
+ bl[114] br[114] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_117 
+ bl[115] br[115] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_118 
+ bl[116] br[116] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_119 
+ bl[117] br[117] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_120 
+ bl[118] br[118] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_121 
+ bl[119] br[119] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_122 
+ bl[120] br[120] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_123 
+ bl[121] br[121] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_124 
+ bl[122] br[122] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_125 
+ bl[123] br[123] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_126 
+ bl[124] br[124] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_127 
+ bl[125] br[125] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_128 
+ bl[126] br[126] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_129 
+ bl[127] br[127] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_130 
+ bl[128] br[128] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_131 
+ bl[129] br[129] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_132 
+ bl[130] br[130] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_133 
+ bl[131] br[131] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_134 
+ bl[132] br[132] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_135 
+ bl[133] br[133] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_136 
+ bl[134] br[134] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_137 
+ bl[135] br[135] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_138 
+ bl[136] br[136] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_139 
+ bl[137] br[137] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_140 
+ bl[138] br[138] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_141 
+ bl[139] br[139] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_142 
+ bl[140] br[140] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_143 
+ bl[141] br[141] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_144 
+ bl[142] br[142] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_145 
+ bl[143] br[143] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_146 
+ bl[144] br[144] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_147 
+ bl[145] br[145] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_148 
+ bl[146] br[146] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_149 
+ bl[147] br[147] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_150 
+ bl[148] br[148] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_151 
+ bl[149] br[149] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_152 
+ bl[150] br[150] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_153 
+ bl[151] br[151] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_154 
+ bl[152] br[152] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_155 
+ bl[153] br[153] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_156 
+ bl[154] br[154] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_157 
+ bl[155] br[155] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_158 
+ bl[156] br[156] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_159 
+ bl[157] br[157] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_160 
+ bl[158] br[158] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_161 
+ bl[159] br[159] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_162 
+ bl[160] br[160] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_163 
+ bl[161] br[161] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_164 
+ bl[162] br[162] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_165 
+ bl[163] br[163] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_166 
+ bl[164] br[164] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_167 
+ bl[165] br[165] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_168 
+ bl[166] br[166] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_169 
+ bl[167] br[167] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_170 
+ bl[168] br[168] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_171 
+ bl[169] br[169] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_172 
+ bl[170] br[170] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_173 
+ bl[171] br[171] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_174 
+ bl[172] br[172] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_175 
+ bl[173] br[173] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_176 
+ bl[174] br[174] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_177 
+ bl[175] br[175] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_178 
+ bl[176] br[176] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_179 
+ bl[177] br[177] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_180 
+ bl[178] br[178] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_181 
+ bl[179] br[179] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_182 
+ bl[180] br[180] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_183 
+ bl[181] br[181] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_184 
+ bl[182] br[182] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_185 
+ bl[183] br[183] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_186 
+ bl[184] br[184] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_187 
+ bl[185] br[185] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_188 
+ bl[186] br[186] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_189 
+ bl[187] br[187] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_190 
+ bl[188] br[188] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_191 
+ bl[189] br[189] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_192 
+ bl[190] br[190] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_193 
+ bl[191] br[191] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_194 
+ bl[192] br[192] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_195 
+ bl[193] br[193] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_196 
+ bl[194] br[194] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_197 
+ bl[195] br[195] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_198 
+ bl[196] br[196] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_199 
+ bl[197] br[197] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_200 
+ bl[198] br[198] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_201 
+ bl[199] br[199] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_202 
+ bl[200] br[200] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_203 
+ bl[201] br[201] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_204 
+ bl[202] br[202] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_205 
+ bl[203] br[203] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_206 
+ bl[204] br[204] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_207 
+ bl[205] br[205] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_208 
+ bl[206] br[206] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_209 
+ bl[207] br[207] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_210 
+ bl[208] br[208] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_211 
+ bl[209] br[209] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_212 
+ bl[210] br[210] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_213 
+ bl[211] br[211] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_214 
+ bl[212] br[212] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_215 
+ bl[213] br[213] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_216 
+ bl[214] br[214] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_217 
+ bl[215] br[215] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_218 
+ bl[216] br[216] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_219 
+ bl[217] br[217] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_220 
+ bl[218] br[218] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_221 
+ bl[219] br[219] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_222 
+ bl[220] br[220] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_223 
+ bl[221] br[221] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_224 
+ bl[222] br[222] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_225 
+ bl[223] br[223] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_226 
+ bl[224] br[224] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_227 
+ bl[225] br[225] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_228 
+ bl[226] br[226] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_229 
+ bl[227] br[227] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_230 
+ bl[228] br[228] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_231 
+ bl[229] br[229] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_232 
+ bl[230] br[230] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_233 
+ bl[231] br[231] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_234 
+ bl[232] br[232] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_235 
+ bl[233] br[233] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_236 
+ bl[234] br[234] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_237 
+ bl[235] br[235] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_238 
+ bl[236] br[236] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_239 
+ bl[237] br[237] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_240 
+ bl[238] br[238] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_241 
+ bl[239] br[239] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_242 
+ bl[240] br[240] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_243 
+ bl[241] br[241] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_244 
+ bl[242] br[242] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_245 
+ bl[243] br[243] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_246 
+ bl[244] br[244] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_247 
+ bl[245] br[245] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_248 
+ bl[246] br[246] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_249 
+ bl[247] br[247] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_250 
+ bl[248] br[248] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_251 
+ bl[249] br[249] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_252 
+ bl[250] br[250] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_253 
+ bl[251] br[251] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_254 
+ bl[252] br[252] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_255 
+ bl[253] br[253] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_256 
+ bl[254] br[254] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_257 
+ bl[255] br[255] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_258 
+ vdd vdd vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_259 
+ vdd vdd vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_0 
+ vdd vdd vss vdd vpb vnb wl[47] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_49_1 
+ rbl rbr vss vdd vpb vnb wl[47] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_49_2 
+ bl[0] br[0] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_3 
+ bl[1] br[1] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_4 
+ bl[2] br[2] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_5 
+ bl[3] br[3] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_6 
+ bl[4] br[4] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_7 
+ bl[5] br[5] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_8 
+ bl[6] br[6] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_9 
+ bl[7] br[7] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_10 
+ bl[8] br[8] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_11 
+ bl[9] br[9] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_12 
+ bl[10] br[10] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_13 
+ bl[11] br[11] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_14 
+ bl[12] br[12] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_15 
+ bl[13] br[13] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_16 
+ bl[14] br[14] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_17 
+ bl[15] br[15] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_18 
+ bl[16] br[16] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_19 
+ bl[17] br[17] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_20 
+ bl[18] br[18] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_21 
+ bl[19] br[19] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_22 
+ bl[20] br[20] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_23 
+ bl[21] br[21] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_24 
+ bl[22] br[22] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_25 
+ bl[23] br[23] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_26 
+ bl[24] br[24] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_27 
+ bl[25] br[25] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_28 
+ bl[26] br[26] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_29 
+ bl[27] br[27] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_30 
+ bl[28] br[28] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_31 
+ bl[29] br[29] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_32 
+ bl[30] br[30] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_33 
+ bl[31] br[31] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_34 
+ bl[32] br[32] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_35 
+ bl[33] br[33] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_36 
+ bl[34] br[34] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_37 
+ bl[35] br[35] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_38 
+ bl[36] br[36] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_39 
+ bl[37] br[37] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_40 
+ bl[38] br[38] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_41 
+ bl[39] br[39] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_42 
+ bl[40] br[40] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_43 
+ bl[41] br[41] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_44 
+ bl[42] br[42] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_45 
+ bl[43] br[43] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_46 
+ bl[44] br[44] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_47 
+ bl[45] br[45] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_48 
+ bl[46] br[46] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_49 
+ bl[47] br[47] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_50 
+ bl[48] br[48] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_51 
+ bl[49] br[49] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_52 
+ bl[50] br[50] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_53 
+ bl[51] br[51] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_54 
+ bl[52] br[52] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_55 
+ bl[53] br[53] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_56 
+ bl[54] br[54] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_57 
+ bl[55] br[55] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_58 
+ bl[56] br[56] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_59 
+ bl[57] br[57] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_60 
+ bl[58] br[58] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_61 
+ bl[59] br[59] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_62 
+ bl[60] br[60] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_63 
+ bl[61] br[61] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_64 
+ bl[62] br[62] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_65 
+ bl[63] br[63] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_66 
+ bl[64] br[64] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_67 
+ bl[65] br[65] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_68 
+ bl[66] br[66] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_69 
+ bl[67] br[67] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_70 
+ bl[68] br[68] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_71 
+ bl[69] br[69] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_72 
+ bl[70] br[70] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_73 
+ bl[71] br[71] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_74 
+ bl[72] br[72] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_75 
+ bl[73] br[73] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_76 
+ bl[74] br[74] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_77 
+ bl[75] br[75] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_78 
+ bl[76] br[76] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_79 
+ bl[77] br[77] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_80 
+ bl[78] br[78] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_81 
+ bl[79] br[79] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_82 
+ bl[80] br[80] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_83 
+ bl[81] br[81] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_84 
+ bl[82] br[82] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_85 
+ bl[83] br[83] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_86 
+ bl[84] br[84] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_87 
+ bl[85] br[85] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_88 
+ bl[86] br[86] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_89 
+ bl[87] br[87] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_90 
+ bl[88] br[88] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_91 
+ bl[89] br[89] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_92 
+ bl[90] br[90] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_93 
+ bl[91] br[91] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_94 
+ bl[92] br[92] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_95 
+ bl[93] br[93] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_96 
+ bl[94] br[94] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_97 
+ bl[95] br[95] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_98 
+ bl[96] br[96] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_99 
+ bl[97] br[97] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_100 
+ bl[98] br[98] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_101 
+ bl[99] br[99] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_102 
+ bl[100] br[100] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_103 
+ bl[101] br[101] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_104 
+ bl[102] br[102] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_105 
+ bl[103] br[103] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_106 
+ bl[104] br[104] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_107 
+ bl[105] br[105] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_108 
+ bl[106] br[106] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_109 
+ bl[107] br[107] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_110 
+ bl[108] br[108] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_111 
+ bl[109] br[109] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_112 
+ bl[110] br[110] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_113 
+ bl[111] br[111] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_114 
+ bl[112] br[112] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_115 
+ bl[113] br[113] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_116 
+ bl[114] br[114] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_117 
+ bl[115] br[115] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_118 
+ bl[116] br[116] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_119 
+ bl[117] br[117] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_120 
+ bl[118] br[118] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_121 
+ bl[119] br[119] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_122 
+ bl[120] br[120] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_123 
+ bl[121] br[121] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_124 
+ bl[122] br[122] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_125 
+ bl[123] br[123] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_126 
+ bl[124] br[124] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_127 
+ bl[125] br[125] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_128 
+ bl[126] br[126] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_129 
+ bl[127] br[127] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_130 
+ bl[128] br[128] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_131 
+ bl[129] br[129] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_132 
+ bl[130] br[130] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_133 
+ bl[131] br[131] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_134 
+ bl[132] br[132] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_135 
+ bl[133] br[133] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_136 
+ bl[134] br[134] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_137 
+ bl[135] br[135] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_138 
+ bl[136] br[136] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_139 
+ bl[137] br[137] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_140 
+ bl[138] br[138] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_141 
+ bl[139] br[139] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_142 
+ bl[140] br[140] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_143 
+ bl[141] br[141] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_144 
+ bl[142] br[142] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_145 
+ bl[143] br[143] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_146 
+ bl[144] br[144] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_147 
+ bl[145] br[145] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_148 
+ bl[146] br[146] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_149 
+ bl[147] br[147] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_150 
+ bl[148] br[148] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_151 
+ bl[149] br[149] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_152 
+ bl[150] br[150] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_153 
+ bl[151] br[151] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_154 
+ bl[152] br[152] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_155 
+ bl[153] br[153] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_156 
+ bl[154] br[154] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_157 
+ bl[155] br[155] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_158 
+ bl[156] br[156] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_159 
+ bl[157] br[157] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_160 
+ bl[158] br[158] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_161 
+ bl[159] br[159] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_162 
+ bl[160] br[160] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_163 
+ bl[161] br[161] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_164 
+ bl[162] br[162] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_165 
+ bl[163] br[163] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_166 
+ bl[164] br[164] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_167 
+ bl[165] br[165] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_168 
+ bl[166] br[166] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_169 
+ bl[167] br[167] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_170 
+ bl[168] br[168] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_171 
+ bl[169] br[169] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_172 
+ bl[170] br[170] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_173 
+ bl[171] br[171] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_174 
+ bl[172] br[172] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_175 
+ bl[173] br[173] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_176 
+ bl[174] br[174] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_177 
+ bl[175] br[175] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_178 
+ bl[176] br[176] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_179 
+ bl[177] br[177] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_180 
+ bl[178] br[178] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_181 
+ bl[179] br[179] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_182 
+ bl[180] br[180] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_183 
+ bl[181] br[181] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_184 
+ bl[182] br[182] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_185 
+ bl[183] br[183] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_186 
+ bl[184] br[184] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_187 
+ bl[185] br[185] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_188 
+ bl[186] br[186] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_189 
+ bl[187] br[187] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_190 
+ bl[188] br[188] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_191 
+ bl[189] br[189] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_192 
+ bl[190] br[190] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_193 
+ bl[191] br[191] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_194 
+ bl[192] br[192] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_195 
+ bl[193] br[193] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_196 
+ bl[194] br[194] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_197 
+ bl[195] br[195] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_198 
+ bl[196] br[196] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_199 
+ bl[197] br[197] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_200 
+ bl[198] br[198] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_201 
+ bl[199] br[199] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_202 
+ bl[200] br[200] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_203 
+ bl[201] br[201] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_204 
+ bl[202] br[202] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_205 
+ bl[203] br[203] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_206 
+ bl[204] br[204] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_207 
+ bl[205] br[205] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_208 
+ bl[206] br[206] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_209 
+ bl[207] br[207] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_210 
+ bl[208] br[208] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_211 
+ bl[209] br[209] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_212 
+ bl[210] br[210] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_213 
+ bl[211] br[211] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_214 
+ bl[212] br[212] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_215 
+ bl[213] br[213] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_216 
+ bl[214] br[214] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_217 
+ bl[215] br[215] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_218 
+ bl[216] br[216] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_219 
+ bl[217] br[217] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_220 
+ bl[218] br[218] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_221 
+ bl[219] br[219] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_222 
+ bl[220] br[220] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_223 
+ bl[221] br[221] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_224 
+ bl[222] br[222] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_225 
+ bl[223] br[223] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_226 
+ bl[224] br[224] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_227 
+ bl[225] br[225] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_228 
+ bl[226] br[226] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_229 
+ bl[227] br[227] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_230 
+ bl[228] br[228] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_231 
+ bl[229] br[229] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_232 
+ bl[230] br[230] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_233 
+ bl[231] br[231] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_234 
+ bl[232] br[232] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_235 
+ bl[233] br[233] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_236 
+ bl[234] br[234] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_237 
+ bl[235] br[235] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_238 
+ bl[236] br[236] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_239 
+ bl[237] br[237] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_240 
+ bl[238] br[238] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_241 
+ bl[239] br[239] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_242 
+ bl[240] br[240] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_243 
+ bl[241] br[241] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_244 
+ bl[242] br[242] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_245 
+ bl[243] br[243] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_246 
+ bl[244] br[244] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_247 
+ bl[245] br[245] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_248 
+ bl[246] br[246] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_249 
+ bl[247] br[247] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_250 
+ bl[248] br[248] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_251 
+ bl[249] br[249] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_252 
+ bl[250] br[250] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_253 
+ bl[251] br[251] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_254 
+ bl[252] br[252] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_255 
+ bl[253] br[253] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_256 
+ bl[254] br[254] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_257 
+ bl[255] br[255] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_258 
+ vdd vdd vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_259 
+ vdd vdd vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_0 
+ vdd vdd vss vdd vpb vnb wl[48] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_50_1 
+ rbl rbr vss vdd vpb vnb wl[48] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_50_2 
+ bl[0] br[0] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_3 
+ bl[1] br[1] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_4 
+ bl[2] br[2] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_5 
+ bl[3] br[3] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_6 
+ bl[4] br[4] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_7 
+ bl[5] br[5] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_8 
+ bl[6] br[6] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_9 
+ bl[7] br[7] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_10 
+ bl[8] br[8] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_11 
+ bl[9] br[9] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_12 
+ bl[10] br[10] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_13 
+ bl[11] br[11] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_14 
+ bl[12] br[12] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_15 
+ bl[13] br[13] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_16 
+ bl[14] br[14] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_17 
+ bl[15] br[15] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_18 
+ bl[16] br[16] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_19 
+ bl[17] br[17] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_20 
+ bl[18] br[18] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_21 
+ bl[19] br[19] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_22 
+ bl[20] br[20] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_23 
+ bl[21] br[21] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_24 
+ bl[22] br[22] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_25 
+ bl[23] br[23] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_26 
+ bl[24] br[24] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_27 
+ bl[25] br[25] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_28 
+ bl[26] br[26] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_29 
+ bl[27] br[27] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_30 
+ bl[28] br[28] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_31 
+ bl[29] br[29] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_32 
+ bl[30] br[30] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_33 
+ bl[31] br[31] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_34 
+ bl[32] br[32] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_35 
+ bl[33] br[33] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_36 
+ bl[34] br[34] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_37 
+ bl[35] br[35] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_38 
+ bl[36] br[36] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_39 
+ bl[37] br[37] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_40 
+ bl[38] br[38] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_41 
+ bl[39] br[39] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_42 
+ bl[40] br[40] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_43 
+ bl[41] br[41] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_44 
+ bl[42] br[42] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_45 
+ bl[43] br[43] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_46 
+ bl[44] br[44] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_47 
+ bl[45] br[45] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_48 
+ bl[46] br[46] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_49 
+ bl[47] br[47] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_50 
+ bl[48] br[48] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_51 
+ bl[49] br[49] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_52 
+ bl[50] br[50] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_53 
+ bl[51] br[51] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_54 
+ bl[52] br[52] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_55 
+ bl[53] br[53] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_56 
+ bl[54] br[54] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_57 
+ bl[55] br[55] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_58 
+ bl[56] br[56] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_59 
+ bl[57] br[57] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_60 
+ bl[58] br[58] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_61 
+ bl[59] br[59] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_62 
+ bl[60] br[60] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_63 
+ bl[61] br[61] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_64 
+ bl[62] br[62] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_65 
+ bl[63] br[63] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_66 
+ bl[64] br[64] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_67 
+ bl[65] br[65] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_68 
+ bl[66] br[66] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_69 
+ bl[67] br[67] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_70 
+ bl[68] br[68] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_71 
+ bl[69] br[69] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_72 
+ bl[70] br[70] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_73 
+ bl[71] br[71] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_74 
+ bl[72] br[72] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_75 
+ bl[73] br[73] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_76 
+ bl[74] br[74] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_77 
+ bl[75] br[75] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_78 
+ bl[76] br[76] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_79 
+ bl[77] br[77] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_80 
+ bl[78] br[78] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_81 
+ bl[79] br[79] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_82 
+ bl[80] br[80] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_83 
+ bl[81] br[81] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_84 
+ bl[82] br[82] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_85 
+ bl[83] br[83] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_86 
+ bl[84] br[84] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_87 
+ bl[85] br[85] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_88 
+ bl[86] br[86] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_89 
+ bl[87] br[87] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_90 
+ bl[88] br[88] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_91 
+ bl[89] br[89] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_92 
+ bl[90] br[90] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_93 
+ bl[91] br[91] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_94 
+ bl[92] br[92] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_95 
+ bl[93] br[93] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_96 
+ bl[94] br[94] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_97 
+ bl[95] br[95] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_98 
+ bl[96] br[96] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_99 
+ bl[97] br[97] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_100 
+ bl[98] br[98] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_101 
+ bl[99] br[99] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_102 
+ bl[100] br[100] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_103 
+ bl[101] br[101] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_104 
+ bl[102] br[102] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_105 
+ bl[103] br[103] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_106 
+ bl[104] br[104] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_107 
+ bl[105] br[105] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_108 
+ bl[106] br[106] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_109 
+ bl[107] br[107] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_110 
+ bl[108] br[108] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_111 
+ bl[109] br[109] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_112 
+ bl[110] br[110] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_113 
+ bl[111] br[111] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_114 
+ bl[112] br[112] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_115 
+ bl[113] br[113] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_116 
+ bl[114] br[114] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_117 
+ bl[115] br[115] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_118 
+ bl[116] br[116] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_119 
+ bl[117] br[117] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_120 
+ bl[118] br[118] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_121 
+ bl[119] br[119] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_122 
+ bl[120] br[120] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_123 
+ bl[121] br[121] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_124 
+ bl[122] br[122] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_125 
+ bl[123] br[123] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_126 
+ bl[124] br[124] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_127 
+ bl[125] br[125] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_128 
+ bl[126] br[126] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_129 
+ bl[127] br[127] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_130 
+ bl[128] br[128] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_131 
+ bl[129] br[129] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_132 
+ bl[130] br[130] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_133 
+ bl[131] br[131] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_134 
+ bl[132] br[132] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_135 
+ bl[133] br[133] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_136 
+ bl[134] br[134] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_137 
+ bl[135] br[135] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_138 
+ bl[136] br[136] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_139 
+ bl[137] br[137] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_140 
+ bl[138] br[138] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_141 
+ bl[139] br[139] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_142 
+ bl[140] br[140] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_143 
+ bl[141] br[141] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_144 
+ bl[142] br[142] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_145 
+ bl[143] br[143] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_146 
+ bl[144] br[144] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_147 
+ bl[145] br[145] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_148 
+ bl[146] br[146] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_149 
+ bl[147] br[147] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_150 
+ bl[148] br[148] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_151 
+ bl[149] br[149] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_152 
+ bl[150] br[150] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_153 
+ bl[151] br[151] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_154 
+ bl[152] br[152] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_155 
+ bl[153] br[153] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_156 
+ bl[154] br[154] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_157 
+ bl[155] br[155] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_158 
+ bl[156] br[156] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_159 
+ bl[157] br[157] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_160 
+ bl[158] br[158] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_161 
+ bl[159] br[159] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_162 
+ bl[160] br[160] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_163 
+ bl[161] br[161] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_164 
+ bl[162] br[162] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_165 
+ bl[163] br[163] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_166 
+ bl[164] br[164] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_167 
+ bl[165] br[165] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_168 
+ bl[166] br[166] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_169 
+ bl[167] br[167] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_170 
+ bl[168] br[168] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_171 
+ bl[169] br[169] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_172 
+ bl[170] br[170] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_173 
+ bl[171] br[171] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_174 
+ bl[172] br[172] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_175 
+ bl[173] br[173] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_176 
+ bl[174] br[174] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_177 
+ bl[175] br[175] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_178 
+ bl[176] br[176] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_179 
+ bl[177] br[177] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_180 
+ bl[178] br[178] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_181 
+ bl[179] br[179] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_182 
+ bl[180] br[180] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_183 
+ bl[181] br[181] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_184 
+ bl[182] br[182] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_185 
+ bl[183] br[183] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_186 
+ bl[184] br[184] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_187 
+ bl[185] br[185] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_188 
+ bl[186] br[186] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_189 
+ bl[187] br[187] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_190 
+ bl[188] br[188] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_191 
+ bl[189] br[189] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_192 
+ bl[190] br[190] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_193 
+ bl[191] br[191] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_194 
+ bl[192] br[192] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_195 
+ bl[193] br[193] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_196 
+ bl[194] br[194] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_197 
+ bl[195] br[195] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_198 
+ bl[196] br[196] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_199 
+ bl[197] br[197] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_200 
+ bl[198] br[198] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_201 
+ bl[199] br[199] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_202 
+ bl[200] br[200] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_203 
+ bl[201] br[201] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_204 
+ bl[202] br[202] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_205 
+ bl[203] br[203] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_206 
+ bl[204] br[204] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_207 
+ bl[205] br[205] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_208 
+ bl[206] br[206] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_209 
+ bl[207] br[207] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_210 
+ bl[208] br[208] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_211 
+ bl[209] br[209] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_212 
+ bl[210] br[210] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_213 
+ bl[211] br[211] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_214 
+ bl[212] br[212] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_215 
+ bl[213] br[213] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_216 
+ bl[214] br[214] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_217 
+ bl[215] br[215] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_218 
+ bl[216] br[216] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_219 
+ bl[217] br[217] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_220 
+ bl[218] br[218] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_221 
+ bl[219] br[219] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_222 
+ bl[220] br[220] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_223 
+ bl[221] br[221] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_224 
+ bl[222] br[222] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_225 
+ bl[223] br[223] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_226 
+ bl[224] br[224] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_227 
+ bl[225] br[225] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_228 
+ bl[226] br[226] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_229 
+ bl[227] br[227] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_230 
+ bl[228] br[228] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_231 
+ bl[229] br[229] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_232 
+ bl[230] br[230] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_233 
+ bl[231] br[231] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_234 
+ bl[232] br[232] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_235 
+ bl[233] br[233] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_236 
+ bl[234] br[234] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_237 
+ bl[235] br[235] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_238 
+ bl[236] br[236] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_239 
+ bl[237] br[237] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_240 
+ bl[238] br[238] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_241 
+ bl[239] br[239] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_242 
+ bl[240] br[240] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_243 
+ bl[241] br[241] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_244 
+ bl[242] br[242] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_245 
+ bl[243] br[243] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_246 
+ bl[244] br[244] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_247 
+ bl[245] br[245] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_248 
+ bl[246] br[246] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_249 
+ bl[247] br[247] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_250 
+ bl[248] br[248] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_251 
+ bl[249] br[249] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_252 
+ bl[250] br[250] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_253 
+ bl[251] br[251] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_254 
+ bl[252] br[252] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_255 
+ bl[253] br[253] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_256 
+ bl[254] br[254] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_257 
+ bl[255] br[255] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_258 
+ vdd vdd vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_259 
+ vdd vdd vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_0 
+ vdd vdd vss vdd vpb vnb wl[49] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_51_1 
+ rbl rbr vss vdd vpb vnb wl[49] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_51_2 
+ bl[0] br[0] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_3 
+ bl[1] br[1] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_4 
+ bl[2] br[2] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_5 
+ bl[3] br[3] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_6 
+ bl[4] br[4] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_7 
+ bl[5] br[5] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_8 
+ bl[6] br[6] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_9 
+ bl[7] br[7] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_10 
+ bl[8] br[8] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_11 
+ bl[9] br[9] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_12 
+ bl[10] br[10] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_13 
+ bl[11] br[11] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_14 
+ bl[12] br[12] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_15 
+ bl[13] br[13] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_16 
+ bl[14] br[14] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_17 
+ bl[15] br[15] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_18 
+ bl[16] br[16] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_19 
+ bl[17] br[17] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_20 
+ bl[18] br[18] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_21 
+ bl[19] br[19] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_22 
+ bl[20] br[20] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_23 
+ bl[21] br[21] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_24 
+ bl[22] br[22] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_25 
+ bl[23] br[23] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_26 
+ bl[24] br[24] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_27 
+ bl[25] br[25] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_28 
+ bl[26] br[26] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_29 
+ bl[27] br[27] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_30 
+ bl[28] br[28] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_31 
+ bl[29] br[29] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_32 
+ bl[30] br[30] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_33 
+ bl[31] br[31] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_34 
+ bl[32] br[32] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_35 
+ bl[33] br[33] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_36 
+ bl[34] br[34] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_37 
+ bl[35] br[35] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_38 
+ bl[36] br[36] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_39 
+ bl[37] br[37] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_40 
+ bl[38] br[38] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_41 
+ bl[39] br[39] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_42 
+ bl[40] br[40] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_43 
+ bl[41] br[41] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_44 
+ bl[42] br[42] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_45 
+ bl[43] br[43] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_46 
+ bl[44] br[44] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_47 
+ bl[45] br[45] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_48 
+ bl[46] br[46] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_49 
+ bl[47] br[47] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_50 
+ bl[48] br[48] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_51 
+ bl[49] br[49] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_52 
+ bl[50] br[50] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_53 
+ bl[51] br[51] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_54 
+ bl[52] br[52] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_55 
+ bl[53] br[53] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_56 
+ bl[54] br[54] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_57 
+ bl[55] br[55] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_58 
+ bl[56] br[56] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_59 
+ bl[57] br[57] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_60 
+ bl[58] br[58] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_61 
+ bl[59] br[59] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_62 
+ bl[60] br[60] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_63 
+ bl[61] br[61] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_64 
+ bl[62] br[62] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_65 
+ bl[63] br[63] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_66 
+ bl[64] br[64] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_67 
+ bl[65] br[65] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_68 
+ bl[66] br[66] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_69 
+ bl[67] br[67] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_70 
+ bl[68] br[68] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_71 
+ bl[69] br[69] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_72 
+ bl[70] br[70] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_73 
+ bl[71] br[71] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_74 
+ bl[72] br[72] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_75 
+ bl[73] br[73] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_76 
+ bl[74] br[74] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_77 
+ bl[75] br[75] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_78 
+ bl[76] br[76] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_79 
+ bl[77] br[77] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_80 
+ bl[78] br[78] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_81 
+ bl[79] br[79] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_82 
+ bl[80] br[80] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_83 
+ bl[81] br[81] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_84 
+ bl[82] br[82] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_85 
+ bl[83] br[83] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_86 
+ bl[84] br[84] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_87 
+ bl[85] br[85] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_88 
+ bl[86] br[86] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_89 
+ bl[87] br[87] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_90 
+ bl[88] br[88] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_91 
+ bl[89] br[89] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_92 
+ bl[90] br[90] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_93 
+ bl[91] br[91] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_94 
+ bl[92] br[92] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_95 
+ bl[93] br[93] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_96 
+ bl[94] br[94] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_97 
+ bl[95] br[95] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_98 
+ bl[96] br[96] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_99 
+ bl[97] br[97] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_100 
+ bl[98] br[98] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_101 
+ bl[99] br[99] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_102 
+ bl[100] br[100] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_103 
+ bl[101] br[101] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_104 
+ bl[102] br[102] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_105 
+ bl[103] br[103] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_106 
+ bl[104] br[104] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_107 
+ bl[105] br[105] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_108 
+ bl[106] br[106] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_109 
+ bl[107] br[107] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_110 
+ bl[108] br[108] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_111 
+ bl[109] br[109] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_112 
+ bl[110] br[110] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_113 
+ bl[111] br[111] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_114 
+ bl[112] br[112] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_115 
+ bl[113] br[113] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_116 
+ bl[114] br[114] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_117 
+ bl[115] br[115] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_118 
+ bl[116] br[116] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_119 
+ bl[117] br[117] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_120 
+ bl[118] br[118] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_121 
+ bl[119] br[119] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_122 
+ bl[120] br[120] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_123 
+ bl[121] br[121] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_124 
+ bl[122] br[122] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_125 
+ bl[123] br[123] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_126 
+ bl[124] br[124] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_127 
+ bl[125] br[125] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_128 
+ bl[126] br[126] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_129 
+ bl[127] br[127] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_130 
+ bl[128] br[128] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_131 
+ bl[129] br[129] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_132 
+ bl[130] br[130] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_133 
+ bl[131] br[131] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_134 
+ bl[132] br[132] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_135 
+ bl[133] br[133] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_136 
+ bl[134] br[134] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_137 
+ bl[135] br[135] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_138 
+ bl[136] br[136] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_139 
+ bl[137] br[137] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_140 
+ bl[138] br[138] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_141 
+ bl[139] br[139] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_142 
+ bl[140] br[140] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_143 
+ bl[141] br[141] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_144 
+ bl[142] br[142] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_145 
+ bl[143] br[143] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_146 
+ bl[144] br[144] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_147 
+ bl[145] br[145] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_148 
+ bl[146] br[146] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_149 
+ bl[147] br[147] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_150 
+ bl[148] br[148] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_151 
+ bl[149] br[149] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_152 
+ bl[150] br[150] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_153 
+ bl[151] br[151] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_154 
+ bl[152] br[152] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_155 
+ bl[153] br[153] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_156 
+ bl[154] br[154] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_157 
+ bl[155] br[155] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_158 
+ bl[156] br[156] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_159 
+ bl[157] br[157] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_160 
+ bl[158] br[158] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_161 
+ bl[159] br[159] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_162 
+ bl[160] br[160] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_163 
+ bl[161] br[161] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_164 
+ bl[162] br[162] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_165 
+ bl[163] br[163] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_166 
+ bl[164] br[164] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_167 
+ bl[165] br[165] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_168 
+ bl[166] br[166] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_169 
+ bl[167] br[167] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_170 
+ bl[168] br[168] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_171 
+ bl[169] br[169] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_172 
+ bl[170] br[170] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_173 
+ bl[171] br[171] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_174 
+ bl[172] br[172] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_175 
+ bl[173] br[173] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_176 
+ bl[174] br[174] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_177 
+ bl[175] br[175] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_178 
+ bl[176] br[176] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_179 
+ bl[177] br[177] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_180 
+ bl[178] br[178] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_181 
+ bl[179] br[179] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_182 
+ bl[180] br[180] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_183 
+ bl[181] br[181] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_184 
+ bl[182] br[182] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_185 
+ bl[183] br[183] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_186 
+ bl[184] br[184] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_187 
+ bl[185] br[185] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_188 
+ bl[186] br[186] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_189 
+ bl[187] br[187] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_190 
+ bl[188] br[188] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_191 
+ bl[189] br[189] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_192 
+ bl[190] br[190] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_193 
+ bl[191] br[191] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_194 
+ bl[192] br[192] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_195 
+ bl[193] br[193] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_196 
+ bl[194] br[194] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_197 
+ bl[195] br[195] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_198 
+ bl[196] br[196] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_199 
+ bl[197] br[197] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_200 
+ bl[198] br[198] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_201 
+ bl[199] br[199] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_202 
+ bl[200] br[200] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_203 
+ bl[201] br[201] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_204 
+ bl[202] br[202] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_205 
+ bl[203] br[203] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_206 
+ bl[204] br[204] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_207 
+ bl[205] br[205] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_208 
+ bl[206] br[206] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_209 
+ bl[207] br[207] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_210 
+ bl[208] br[208] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_211 
+ bl[209] br[209] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_212 
+ bl[210] br[210] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_213 
+ bl[211] br[211] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_214 
+ bl[212] br[212] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_215 
+ bl[213] br[213] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_216 
+ bl[214] br[214] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_217 
+ bl[215] br[215] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_218 
+ bl[216] br[216] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_219 
+ bl[217] br[217] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_220 
+ bl[218] br[218] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_221 
+ bl[219] br[219] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_222 
+ bl[220] br[220] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_223 
+ bl[221] br[221] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_224 
+ bl[222] br[222] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_225 
+ bl[223] br[223] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_226 
+ bl[224] br[224] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_227 
+ bl[225] br[225] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_228 
+ bl[226] br[226] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_229 
+ bl[227] br[227] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_230 
+ bl[228] br[228] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_231 
+ bl[229] br[229] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_232 
+ bl[230] br[230] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_233 
+ bl[231] br[231] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_234 
+ bl[232] br[232] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_235 
+ bl[233] br[233] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_236 
+ bl[234] br[234] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_237 
+ bl[235] br[235] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_238 
+ bl[236] br[236] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_239 
+ bl[237] br[237] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_240 
+ bl[238] br[238] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_241 
+ bl[239] br[239] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_242 
+ bl[240] br[240] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_243 
+ bl[241] br[241] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_244 
+ bl[242] br[242] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_245 
+ bl[243] br[243] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_246 
+ bl[244] br[244] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_247 
+ bl[245] br[245] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_248 
+ bl[246] br[246] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_249 
+ bl[247] br[247] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_250 
+ bl[248] br[248] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_251 
+ bl[249] br[249] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_252 
+ bl[250] br[250] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_253 
+ bl[251] br[251] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_254 
+ bl[252] br[252] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_255 
+ bl[253] br[253] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_256 
+ bl[254] br[254] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_257 
+ bl[255] br[255] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_258 
+ vdd vdd vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_259 
+ vdd vdd vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_0 
+ vdd vdd vss vdd vpb vnb wl[50] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_52_1 
+ rbl rbr vss vdd vpb vnb wl[50] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_52_2 
+ bl[0] br[0] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_3 
+ bl[1] br[1] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_4 
+ bl[2] br[2] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_5 
+ bl[3] br[3] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_6 
+ bl[4] br[4] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_7 
+ bl[5] br[5] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_8 
+ bl[6] br[6] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_9 
+ bl[7] br[7] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_10 
+ bl[8] br[8] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_11 
+ bl[9] br[9] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_12 
+ bl[10] br[10] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_13 
+ bl[11] br[11] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_14 
+ bl[12] br[12] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_15 
+ bl[13] br[13] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_16 
+ bl[14] br[14] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_17 
+ bl[15] br[15] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_18 
+ bl[16] br[16] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_19 
+ bl[17] br[17] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_20 
+ bl[18] br[18] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_21 
+ bl[19] br[19] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_22 
+ bl[20] br[20] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_23 
+ bl[21] br[21] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_24 
+ bl[22] br[22] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_25 
+ bl[23] br[23] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_26 
+ bl[24] br[24] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_27 
+ bl[25] br[25] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_28 
+ bl[26] br[26] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_29 
+ bl[27] br[27] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_30 
+ bl[28] br[28] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_31 
+ bl[29] br[29] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_32 
+ bl[30] br[30] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_33 
+ bl[31] br[31] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_34 
+ bl[32] br[32] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_35 
+ bl[33] br[33] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_36 
+ bl[34] br[34] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_37 
+ bl[35] br[35] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_38 
+ bl[36] br[36] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_39 
+ bl[37] br[37] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_40 
+ bl[38] br[38] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_41 
+ bl[39] br[39] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_42 
+ bl[40] br[40] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_43 
+ bl[41] br[41] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_44 
+ bl[42] br[42] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_45 
+ bl[43] br[43] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_46 
+ bl[44] br[44] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_47 
+ bl[45] br[45] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_48 
+ bl[46] br[46] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_49 
+ bl[47] br[47] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_50 
+ bl[48] br[48] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_51 
+ bl[49] br[49] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_52 
+ bl[50] br[50] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_53 
+ bl[51] br[51] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_54 
+ bl[52] br[52] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_55 
+ bl[53] br[53] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_56 
+ bl[54] br[54] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_57 
+ bl[55] br[55] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_58 
+ bl[56] br[56] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_59 
+ bl[57] br[57] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_60 
+ bl[58] br[58] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_61 
+ bl[59] br[59] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_62 
+ bl[60] br[60] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_63 
+ bl[61] br[61] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_64 
+ bl[62] br[62] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_65 
+ bl[63] br[63] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_66 
+ bl[64] br[64] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_67 
+ bl[65] br[65] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_68 
+ bl[66] br[66] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_69 
+ bl[67] br[67] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_70 
+ bl[68] br[68] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_71 
+ bl[69] br[69] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_72 
+ bl[70] br[70] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_73 
+ bl[71] br[71] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_74 
+ bl[72] br[72] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_75 
+ bl[73] br[73] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_76 
+ bl[74] br[74] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_77 
+ bl[75] br[75] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_78 
+ bl[76] br[76] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_79 
+ bl[77] br[77] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_80 
+ bl[78] br[78] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_81 
+ bl[79] br[79] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_82 
+ bl[80] br[80] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_83 
+ bl[81] br[81] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_84 
+ bl[82] br[82] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_85 
+ bl[83] br[83] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_86 
+ bl[84] br[84] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_87 
+ bl[85] br[85] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_88 
+ bl[86] br[86] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_89 
+ bl[87] br[87] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_90 
+ bl[88] br[88] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_91 
+ bl[89] br[89] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_92 
+ bl[90] br[90] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_93 
+ bl[91] br[91] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_94 
+ bl[92] br[92] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_95 
+ bl[93] br[93] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_96 
+ bl[94] br[94] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_97 
+ bl[95] br[95] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_98 
+ bl[96] br[96] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_99 
+ bl[97] br[97] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_100 
+ bl[98] br[98] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_101 
+ bl[99] br[99] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_102 
+ bl[100] br[100] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_103 
+ bl[101] br[101] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_104 
+ bl[102] br[102] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_105 
+ bl[103] br[103] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_106 
+ bl[104] br[104] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_107 
+ bl[105] br[105] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_108 
+ bl[106] br[106] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_109 
+ bl[107] br[107] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_110 
+ bl[108] br[108] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_111 
+ bl[109] br[109] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_112 
+ bl[110] br[110] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_113 
+ bl[111] br[111] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_114 
+ bl[112] br[112] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_115 
+ bl[113] br[113] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_116 
+ bl[114] br[114] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_117 
+ bl[115] br[115] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_118 
+ bl[116] br[116] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_119 
+ bl[117] br[117] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_120 
+ bl[118] br[118] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_121 
+ bl[119] br[119] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_122 
+ bl[120] br[120] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_123 
+ bl[121] br[121] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_124 
+ bl[122] br[122] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_125 
+ bl[123] br[123] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_126 
+ bl[124] br[124] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_127 
+ bl[125] br[125] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_128 
+ bl[126] br[126] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_129 
+ bl[127] br[127] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_130 
+ bl[128] br[128] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_131 
+ bl[129] br[129] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_132 
+ bl[130] br[130] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_133 
+ bl[131] br[131] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_134 
+ bl[132] br[132] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_135 
+ bl[133] br[133] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_136 
+ bl[134] br[134] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_137 
+ bl[135] br[135] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_138 
+ bl[136] br[136] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_139 
+ bl[137] br[137] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_140 
+ bl[138] br[138] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_141 
+ bl[139] br[139] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_142 
+ bl[140] br[140] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_143 
+ bl[141] br[141] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_144 
+ bl[142] br[142] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_145 
+ bl[143] br[143] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_146 
+ bl[144] br[144] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_147 
+ bl[145] br[145] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_148 
+ bl[146] br[146] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_149 
+ bl[147] br[147] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_150 
+ bl[148] br[148] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_151 
+ bl[149] br[149] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_152 
+ bl[150] br[150] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_153 
+ bl[151] br[151] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_154 
+ bl[152] br[152] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_155 
+ bl[153] br[153] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_156 
+ bl[154] br[154] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_157 
+ bl[155] br[155] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_158 
+ bl[156] br[156] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_159 
+ bl[157] br[157] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_160 
+ bl[158] br[158] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_161 
+ bl[159] br[159] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_162 
+ bl[160] br[160] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_163 
+ bl[161] br[161] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_164 
+ bl[162] br[162] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_165 
+ bl[163] br[163] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_166 
+ bl[164] br[164] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_167 
+ bl[165] br[165] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_168 
+ bl[166] br[166] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_169 
+ bl[167] br[167] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_170 
+ bl[168] br[168] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_171 
+ bl[169] br[169] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_172 
+ bl[170] br[170] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_173 
+ bl[171] br[171] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_174 
+ bl[172] br[172] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_175 
+ bl[173] br[173] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_176 
+ bl[174] br[174] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_177 
+ bl[175] br[175] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_178 
+ bl[176] br[176] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_179 
+ bl[177] br[177] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_180 
+ bl[178] br[178] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_181 
+ bl[179] br[179] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_182 
+ bl[180] br[180] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_183 
+ bl[181] br[181] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_184 
+ bl[182] br[182] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_185 
+ bl[183] br[183] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_186 
+ bl[184] br[184] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_187 
+ bl[185] br[185] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_188 
+ bl[186] br[186] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_189 
+ bl[187] br[187] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_190 
+ bl[188] br[188] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_191 
+ bl[189] br[189] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_192 
+ bl[190] br[190] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_193 
+ bl[191] br[191] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_194 
+ bl[192] br[192] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_195 
+ bl[193] br[193] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_196 
+ bl[194] br[194] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_197 
+ bl[195] br[195] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_198 
+ bl[196] br[196] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_199 
+ bl[197] br[197] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_200 
+ bl[198] br[198] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_201 
+ bl[199] br[199] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_202 
+ bl[200] br[200] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_203 
+ bl[201] br[201] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_204 
+ bl[202] br[202] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_205 
+ bl[203] br[203] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_206 
+ bl[204] br[204] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_207 
+ bl[205] br[205] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_208 
+ bl[206] br[206] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_209 
+ bl[207] br[207] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_210 
+ bl[208] br[208] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_211 
+ bl[209] br[209] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_212 
+ bl[210] br[210] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_213 
+ bl[211] br[211] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_214 
+ bl[212] br[212] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_215 
+ bl[213] br[213] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_216 
+ bl[214] br[214] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_217 
+ bl[215] br[215] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_218 
+ bl[216] br[216] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_219 
+ bl[217] br[217] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_220 
+ bl[218] br[218] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_221 
+ bl[219] br[219] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_222 
+ bl[220] br[220] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_223 
+ bl[221] br[221] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_224 
+ bl[222] br[222] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_225 
+ bl[223] br[223] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_226 
+ bl[224] br[224] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_227 
+ bl[225] br[225] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_228 
+ bl[226] br[226] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_229 
+ bl[227] br[227] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_230 
+ bl[228] br[228] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_231 
+ bl[229] br[229] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_232 
+ bl[230] br[230] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_233 
+ bl[231] br[231] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_234 
+ bl[232] br[232] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_235 
+ bl[233] br[233] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_236 
+ bl[234] br[234] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_237 
+ bl[235] br[235] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_238 
+ bl[236] br[236] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_239 
+ bl[237] br[237] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_240 
+ bl[238] br[238] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_241 
+ bl[239] br[239] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_242 
+ bl[240] br[240] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_243 
+ bl[241] br[241] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_244 
+ bl[242] br[242] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_245 
+ bl[243] br[243] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_246 
+ bl[244] br[244] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_247 
+ bl[245] br[245] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_248 
+ bl[246] br[246] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_249 
+ bl[247] br[247] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_250 
+ bl[248] br[248] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_251 
+ bl[249] br[249] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_252 
+ bl[250] br[250] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_253 
+ bl[251] br[251] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_254 
+ bl[252] br[252] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_255 
+ bl[253] br[253] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_256 
+ bl[254] br[254] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_257 
+ bl[255] br[255] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_258 
+ vdd vdd vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_259 
+ vdd vdd vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_0 
+ vdd vdd vss vdd vpb vnb wl[51] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_53_1 
+ rbl rbr vss vdd vpb vnb wl[51] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_53_2 
+ bl[0] br[0] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_3 
+ bl[1] br[1] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_4 
+ bl[2] br[2] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_5 
+ bl[3] br[3] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_6 
+ bl[4] br[4] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_7 
+ bl[5] br[5] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_8 
+ bl[6] br[6] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_9 
+ bl[7] br[7] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_10 
+ bl[8] br[8] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_11 
+ bl[9] br[9] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_12 
+ bl[10] br[10] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_13 
+ bl[11] br[11] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_14 
+ bl[12] br[12] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_15 
+ bl[13] br[13] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_16 
+ bl[14] br[14] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_17 
+ bl[15] br[15] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_18 
+ bl[16] br[16] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_19 
+ bl[17] br[17] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_20 
+ bl[18] br[18] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_21 
+ bl[19] br[19] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_22 
+ bl[20] br[20] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_23 
+ bl[21] br[21] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_24 
+ bl[22] br[22] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_25 
+ bl[23] br[23] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_26 
+ bl[24] br[24] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_27 
+ bl[25] br[25] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_28 
+ bl[26] br[26] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_29 
+ bl[27] br[27] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_30 
+ bl[28] br[28] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_31 
+ bl[29] br[29] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_32 
+ bl[30] br[30] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_33 
+ bl[31] br[31] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_34 
+ bl[32] br[32] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_35 
+ bl[33] br[33] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_36 
+ bl[34] br[34] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_37 
+ bl[35] br[35] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_38 
+ bl[36] br[36] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_39 
+ bl[37] br[37] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_40 
+ bl[38] br[38] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_41 
+ bl[39] br[39] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_42 
+ bl[40] br[40] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_43 
+ bl[41] br[41] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_44 
+ bl[42] br[42] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_45 
+ bl[43] br[43] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_46 
+ bl[44] br[44] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_47 
+ bl[45] br[45] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_48 
+ bl[46] br[46] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_49 
+ bl[47] br[47] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_50 
+ bl[48] br[48] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_51 
+ bl[49] br[49] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_52 
+ bl[50] br[50] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_53 
+ bl[51] br[51] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_54 
+ bl[52] br[52] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_55 
+ bl[53] br[53] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_56 
+ bl[54] br[54] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_57 
+ bl[55] br[55] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_58 
+ bl[56] br[56] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_59 
+ bl[57] br[57] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_60 
+ bl[58] br[58] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_61 
+ bl[59] br[59] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_62 
+ bl[60] br[60] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_63 
+ bl[61] br[61] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_64 
+ bl[62] br[62] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_65 
+ bl[63] br[63] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_66 
+ bl[64] br[64] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_67 
+ bl[65] br[65] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_68 
+ bl[66] br[66] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_69 
+ bl[67] br[67] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_70 
+ bl[68] br[68] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_71 
+ bl[69] br[69] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_72 
+ bl[70] br[70] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_73 
+ bl[71] br[71] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_74 
+ bl[72] br[72] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_75 
+ bl[73] br[73] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_76 
+ bl[74] br[74] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_77 
+ bl[75] br[75] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_78 
+ bl[76] br[76] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_79 
+ bl[77] br[77] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_80 
+ bl[78] br[78] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_81 
+ bl[79] br[79] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_82 
+ bl[80] br[80] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_83 
+ bl[81] br[81] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_84 
+ bl[82] br[82] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_85 
+ bl[83] br[83] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_86 
+ bl[84] br[84] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_87 
+ bl[85] br[85] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_88 
+ bl[86] br[86] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_89 
+ bl[87] br[87] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_90 
+ bl[88] br[88] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_91 
+ bl[89] br[89] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_92 
+ bl[90] br[90] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_93 
+ bl[91] br[91] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_94 
+ bl[92] br[92] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_95 
+ bl[93] br[93] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_96 
+ bl[94] br[94] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_97 
+ bl[95] br[95] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_98 
+ bl[96] br[96] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_99 
+ bl[97] br[97] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_100 
+ bl[98] br[98] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_101 
+ bl[99] br[99] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_102 
+ bl[100] br[100] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_103 
+ bl[101] br[101] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_104 
+ bl[102] br[102] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_105 
+ bl[103] br[103] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_106 
+ bl[104] br[104] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_107 
+ bl[105] br[105] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_108 
+ bl[106] br[106] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_109 
+ bl[107] br[107] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_110 
+ bl[108] br[108] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_111 
+ bl[109] br[109] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_112 
+ bl[110] br[110] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_113 
+ bl[111] br[111] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_114 
+ bl[112] br[112] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_115 
+ bl[113] br[113] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_116 
+ bl[114] br[114] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_117 
+ bl[115] br[115] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_118 
+ bl[116] br[116] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_119 
+ bl[117] br[117] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_120 
+ bl[118] br[118] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_121 
+ bl[119] br[119] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_122 
+ bl[120] br[120] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_123 
+ bl[121] br[121] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_124 
+ bl[122] br[122] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_125 
+ bl[123] br[123] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_126 
+ bl[124] br[124] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_127 
+ bl[125] br[125] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_128 
+ bl[126] br[126] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_129 
+ bl[127] br[127] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_130 
+ bl[128] br[128] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_131 
+ bl[129] br[129] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_132 
+ bl[130] br[130] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_133 
+ bl[131] br[131] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_134 
+ bl[132] br[132] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_135 
+ bl[133] br[133] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_136 
+ bl[134] br[134] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_137 
+ bl[135] br[135] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_138 
+ bl[136] br[136] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_139 
+ bl[137] br[137] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_140 
+ bl[138] br[138] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_141 
+ bl[139] br[139] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_142 
+ bl[140] br[140] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_143 
+ bl[141] br[141] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_144 
+ bl[142] br[142] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_145 
+ bl[143] br[143] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_146 
+ bl[144] br[144] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_147 
+ bl[145] br[145] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_148 
+ bl[146] br[146] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_149 
+ bl[147] br[147] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_150 
+ bl[148] br[148] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_151 
+ bl[149] br[149] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_152 
+ bl[150] br[150] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_153 
+ bl[151] br[151] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_154 
+ bl[152] br[152] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_155 
+ bl[153] br[153] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_156 
+ bl[154] br[154] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_157 
+ bl[155] br[155] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_158 
+ bl[156] br[156] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_159 
+ bl[157] br[157] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_160 
+ bl[158] br[158] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_161 
+ bl[159] br[159] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_162 
+ bl[160] br[160] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_163 
+ bl[161] br[161] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_164 
+ bl[162] br[162] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_165 
+ bl[163] br[163] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_166 
+ bl[164] br[164] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_167 
+ bl[165] br[165] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_168 
+ bl[166] br[166] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_169 
+ bl[167] br[167] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_170 
+ bl[168] br[168] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_171 
+ bl[169] br[169] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_172 
+ bl[170] br[170] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_173 
+ bl[171] br[171] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_174 
+ bl[172] br[172] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_175 
+ bl[173] br[173] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_176 
+ bl[174] br[174] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_177 
+ bl[175] br[175] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_178 
+ bl[176] br[176] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_179 
+ bl[177] br[177] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_180 
+ bl[178] br[178] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_181 
+ bl[179] br[179] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_182 
+ bl[180] br[180] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_183 
+ bl[181] br[181] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_184 
+ bl[182] br[182] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_185 
+ bl[183] br[183] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_186 
+ bl[184] br[184] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_187 
+ bl[185] br[185] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_188 
+ bl[186] br[186] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_189 
+ bl[187] br[187] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_190 
+ bl[188] br[188] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_191 
+ bl[189] br[189] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_192 
+ bl[190] br[190] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_193 
+ bl[191] br[191] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_194 
+ bl[192] br[192] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_195 
+ bl[193] br[193] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_196 
+ bl[194] br[194] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_197 
+ bl[195] br[195] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_198 
+ bl[196] br[196] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_199 
+ bl[197] br[197] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_200 
+ bl[198] br[198] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_201 
+ bl[199] br[199] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_202 
+ bl[200] br[200] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_203 
+ bl[201] br[201] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_204 
+ bl[202] br[202] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_205 
+ bl[203] br[203] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_206 
+ bl[204] br[204] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_207 
+ bl[205] br[205] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_208 
+ bl[206] br[206] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_209 
+ bl[207] br[207] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_210 
+ bl[208] br[208] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_211 
+ bl[209] br[209] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_212 
+ bl[210] br[210] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_213 
+ bl[211] br[211] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_214 
+ bl[212] br[212] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_215 
+ bl[213] br[213] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_216 
+ bl[214] br[214] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_217 
+ bl[215] br[215] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_218 
+ bl[216] br[216] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_219 
+ bl[217] br[217] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_220 
+ bl[218] br[218] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_221 
+ bl[219] br[219] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_222 
+ bl[220] br[220] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_223 
+ bl[221] br[221] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_224 
+ bl[222] br[222] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_225 
+ bl[223] br[223] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_226 
+ bl[224] br[224] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_227 
+ bl[225] br[225] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_228 
+ bl[226] br[226] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_229 
+ bl[227] br[227] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_230 
+ bl[228] br[228] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_231 
+ bl[229] br[229] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_232 
+ bl[230] br[230] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_233 
+ bl[231] br[231] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_234 
+ bl[232] br[232] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_235 
+ bl[233] br[233] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_236 
+ bl[234] br[234] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_237 
+ bl[235] br[235] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_238 
+ bl[236] br[236] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_239 
+ bl[237] br[237] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_240 
+ bl[238] br[238] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_241 
+ bl[239] br[239] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_242 
+ bl[240] br[240] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_243 
+ bl[241] br[241] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_244 
+ bl[242] br[242] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_245 
+ bl[243] br[243] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_246 
+ bl[244] br[244] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_247 
+ bl[245] br[245] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_248 
+ bl[246] br[246] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_249 
+ bl[247] br[247] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_250 
+ bl[248] br[248] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_251 
+ bl[249] br[249] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_252 
+ bl[250] br[250] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_253 
+ bl[251] br[251] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_254 
+ bl[252] br[252] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_255 
+ bl[253] br[253] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_256 
+ bl[254] br[254] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_257 
+ bl[255] br[255] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_258 
+ vdd vdd vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_259 
+ vdd vdd vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_0 
+ vdd vdd vss vdd vpb vnb wl[52] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_54_1 
+ rbl rbr vss vdd vpb vnb wl[52] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_54_2 
+ bl[0] br[0] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_3 
+ bl[1] br[1] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_4 
+ bl[2] br[2] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_5 
+ bl[3] br[3] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_6 
+ bl[4] br[4] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_7 
+ bl[5] br[5] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_8 
+ bl[6] br[6] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_9 
+ bl[7] br[7] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_10 
+ bl[8] br[8] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_11 
+ bl[9] br[9] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_12 
+ bl[10] br[10] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_13 
+ bl[11] br[11] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_14 
+ bl[12] br[12] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_15 
+ bl[13] br[13] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_16 
+ bl[14] br[14] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_17 
+ bl[15] br[15] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_18 
+ bl[16] br[16] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_19 
+ bl[17] br[17] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_20 
+ bl[18] br[18] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_21 
+ bl[19] br[19] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_22 
+ bl[20] br[20] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_23 
+ bl[21] br[21] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_24 
+ bl[22] br[22] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_25 
+ bl[23] br[23] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_26 
+ bl[24] br[24] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_27 
+ bl[25] br[25] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_28 
+ bl[26] br[26] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_29 
+ bl[27] br[27] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_30 
+ bl[28] br[28] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_31 
+ bl[29] br[29] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_32 
+ bl[30] br[30] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_33 
+ bl[31] br[31] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_34 
+ bl[32] br[32] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_35 
+ bl[33] br[33] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_36 
+ bl[34] br[34] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_37 
+ bl[35] br[35] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_38 
+ bl[36] br[36] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_39 
+ bl[37] br[37] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_40 
+ bl[38] br[38] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_41 
+ bl[39] br[39] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_42 
+ bl[40] br[40] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_43 
+ bl[41] br[41] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_44 
+ bl[42] br[42] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_45 
+ bl[43] br[43] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_46 
+ bl[44] br[44] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_47 
+ bl[45] br[45] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_48 
+ bl[46] br[46] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_49 
+ bl[47] br[47] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_50 
+ bl[48] br[48] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_51 
+ bl[49] br[49] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_52 
+ bl[50] br[50] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_53 
+ bl[51] br[51] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_54 
+ bl[52] br[52] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_55 
+ bl[53] br[53] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_56 
+ bl[54] br[54] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_57 
+ bl[55] br[55] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_58 
+ bl[56] br[56] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_59 
+ bl[57] br[57] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_60 
+ bl[58] br[58] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_61 
+ bl[59] br[59] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_62 
+ bl[60] br[60] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_63 
+ bl[61] br[61] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_64 
+ bl[62] br[62] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_65 
+ bl[63] br[63] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_66 
+ bl[64] br[64] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_67 
+ bl[65] br[65] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_68 
+ bl[66] br[66] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_69 
+ bl[67] br[67] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_70 
+ bl[68] br[68] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_71 
+ bl[69] br[69] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_72 
+ bl[70] br[70] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_73 
+ bl[71] br[71] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_74 
+ bl[72] br[72] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_75 
+ bl[73] br[73] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_76 
+ bl[74] br[74] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_77 
+ bl[75] br[75] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_78 
+ bl[76] br[76] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_79 
+ bl[77] br[77] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_80 
+ bl[78] br[78] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_81 
+ bl[79] br[79] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_82 
+ bl[80] br[80] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_83 
+ bl[81] br[81] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_84 
+ bl[82] br[82] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_85 
+ bl[83] br[83] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_86 
+ bl[84] br[84] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_87 
+ bl[85] br[85] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_88 
+ bl[86] br[86] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_89 
+ bl[87] br[87] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_90 
+ bl[88] br[88] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_91 
+ bl[89] br[89] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_92 
+ bl[90] br[90] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_93 
+ bl[91] br[91] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_94 
+ bl[92] br[92] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_95 
+ bl[93] br[93] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_96 
+ bl[94] br[94] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_97 
+ bl[95] br[95] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_98 
+ bl[96] br[96] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_99 
+ bl[97] br[97] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_100 
+ bl[98] br[98] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_101 
+ bl[99] br[99] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_102 
+ bl[100] br[100] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_103 
+ bl[101] br[101] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_104 
+ bl[102] br[102] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_105 
+ bl[103] br[103] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_106 
+ bl[104] br[104] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_107 
+ bl[105] br[105] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_108 
+ bl[106] br[106] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_109 
+ bl[107] br[107] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_110 
+ bl[108] br[108] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_111 
+ bl[109] br[109] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_112 
+ bl[110] br[110] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_113 
+ bl[111] br[111] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_114 
+ bl[112] br[112] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_115 
+ bl[113] br[113] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_116 
+ bl[114] br[114] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_117 
+ bl[115] br[115] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_118 
+ bl[116] br[116] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_119 
+ bl[117] br[117] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_120 
+ bl[118] br[118] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_121 
+ bl[119] br[119] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_122 
+ bl[120] br[120] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_123 
+ bl[121] br[121] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_124 
+ bl[122] br[122] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_125 
+ bl[123] br[123] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_126 
+ bl[124] br[124] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_127 
+ bl[125] br[125] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_128 
+ bl[126] br[126] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_129 
+ bl[127] br[127] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_130 
+ bl[128] br[128] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_131 
+ bl[129] br[129] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_132 
+ bl[130] br[130] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_133 
+ bl[131] br[131] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_134 
+ bl[132] br[132] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_135 
+ bl[133] br[133] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_136 
+ bl[134] br[134] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_137 
+ bl[135] br[135] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_138 
+ bl[136] br[136] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_139 
+ bl[137] br[137] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_140 
+ bl[138] br[138] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_141 
+ bl[139] br[139] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_142 
+ bl[140] br[140] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_143 
+ bl[141] br[141] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_144 
+ bl[142] br[142] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_145 
+ bl[143] br[143] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_146 
+ bl[144] br[144] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_147 
+ bl[145] br[145] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_148 
+ bl[146] br[146] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_149 
+ bl[147] br[147] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_150 
+ bl[148] br[148] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_151 
+ bl[149] br[149] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_152 
+ bl[150] br[150] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_153 
+ bl[151] br[151] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_154 
+ bl[152] br[152] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_155 
+ bl[153] br[153] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_156 
+ bl[154] br[154] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_157 
+ bl[155] br[155] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_158 
+ bl[156] br[156] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_159 
+ bl[157] br[157] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_160 
+ bl[158] br[158] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_161 
+ bl[159] br[159] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_162 
+ bl[160] br[160] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_163 
+ bl[161] br[161] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_164 
+ bl[162] br[162] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_165 
+ bl[163] br[163] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_166 
+ bl[164] br[164] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_167 
+ bl[165] br[165] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_168 
+ bl[166] br[166] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_169 
+ bl[167] br[167] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_170 
+ bl[168] br[168] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_171 
+ bl[169] br[169] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_172 
+ bl[170] br[170] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_173 
+ bl[171] br[171] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_174 
+ bl[172] br[172] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_175 
+ bl[173] br[173] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_176 
+ bl[174] br[174] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_177 
+ bl[175] br[175] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_178 
+ bl[176] br[176] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_179 
+ bl[177] br[177] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_180 
+ bl[178] br[178] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_181 
+ bl[179] br[179] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_182 
+ bl[180] br[180] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_183 
+ bl[181] br[181] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_184 
+ bl[182] br[182] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_185 
+ bl[183] br[183] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_186 
+ bl[184] br[184] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_187 
+ bl[185] br[185] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_188 
+ bl[186] br[186] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_189 
+ bl[187] br[187] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_190 
+ bl[188] br[188] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_191 
+ bl[189] br[189] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_192 
+ bl[190] br[190] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_193 
+ bl[191] br[191] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_194 
+ bl[192] br[192] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_195 
+ bl[193] br[193] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_196 
+ bl[194] br[194] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_197 
+ bl[195] br[195] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_198 
+ bl[196] br[196] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_199 
+ bl[197] br[197] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_200 
+ bl[198] br[198] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_201 
+ bl[199] br[199] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_202 
+ bl[200] br[200] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_203 
+ bl[201] br[201] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_204 
+ bl[202] br[202] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_205 
+ bl[203] br[203] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_206 
+ bl[204] br[204] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_207 
+ bl[205] br[205] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_208 
+ bl[206] br[206] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_209 
+ bl[207] br[207] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_210 
+ bl[208] br[208] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_211 
+ bl[209] br[209] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_212 
+ bl[210] br[210] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_213 
+ bl[211] br[211] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_214 
+ bl[212] br[212] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_215 
+ bl[213] br[213] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_216 
+ bl[214] br[214] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_217 
+ bl[215] br[215] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_218 
+ bl[216] br[216] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_219 
+ bl[217] br[217] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_220 
+ bl[218] br[218] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_221 
+ bl[219] br[219] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_222 
+ bl[220] br[220] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_223 
+ bl[221] br[221] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_224 
+ bl[222] br[222] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_225 
+ bl[223] br[223] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_226 
+ bl[224] br[224] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_227 
+ bl[225] br[225] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_228 
+ bl[226] br[226] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_229 
+ bl[227] br[227] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_230 
+ bl[228] br[228] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_231 
+ bl[229] br[229] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_232 
+ bl[230] br[230] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_233 
+ bl[231] br[231] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_234 
+ bl[232] br[232] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_235 
+ bl[233] br[233] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_236 
+ bl[234] br[234] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_237 
+ bl[235] br[235] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_238 
+ bl[236] br[236] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_239 
+ bl[237] br[237] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_240 
+ bl[238] br[238] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_241 
+ bl[239] br[239] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_242 
+ bl[240] br[240] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_243 
+ bl[241] br[241] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_244 
+ bl[242] br[242] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_245 
+ bl[243] br[243] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_246 
+ bl[244] br[244] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_247 
+ bl[245] br[245] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_248 
+ bl[246] br[246] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_249 
+ bl[247] br[247] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_250 
+ bl[248] br[248] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_251 
+ bl[249] br[249] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_252 
+ bl[250] br[250] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_253 
+ bl[251] br[251] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_254 
+ bl[252] br[252] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_255 
+ bl[253] br[253] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_256 
+ bl[254] br[254] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_257 
+ bl[255] br[255] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_258 
+ vdd vdd vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_259 
+ vdd vdd vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_0 
+ vdd vdd vss vdd vpb vnb wl[53] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_55_1 
+ rbl rbr vss vdd vpb vnb wl[53] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_55_2 
+ bl[0] br[0] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_3 
+ bl[1] br[1] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_4 
+ bl[2] br[2] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_5 
+ bl[3] br[3] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_6 
+ bl[4] br[4] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_7 
+ bl[5] br[5] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_8 
+ bl[6] br[6] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_9 
+ bl[7] br[7] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_10 
+ bl[8] br[8] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_11 
+ bl[9] br[9] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_12 
+ bl[10] br[10] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_13 
+ bl[11] br[11] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_14 
+ bl[12] br[12] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_15 
+ bl[13] br[13] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_16 
+ bl[14] br[14] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_17 
+ bl[15] br[15] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_18 
+ bl[16] br[16] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_19 
+ bl[17] br[17] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_20 
+ bl[18] br[18] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_21 
+ bl[19] br[19] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_22 
+ bl[20] br[20] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_23 
+ bl[21] br[21] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_24 
+ bl[22] br[22] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_25 
+ bl[23] br[23] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_26 
+ bl[24] br[24] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_27 
+ bl[25] br[25] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_28 
+ bl[26] br[26] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_29 
+ bl[27] br[27] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_30 
+ bl[28] br[28] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_31 
+ bl[29] br[29] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_32 
+ bl[30] br[30] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_33 
+ bl[31] br[31] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_34 
+ bl[32] br[32] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_35 
+ bl[33] br[33] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_36 
+ bl[34] br[34] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_37 
+ bl[35] br[35] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_38 
+ bl[36] br[36] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_39 
+ bl[37] br[37] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_40 
+ bl[38] br[38] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_41 
+ bl[39] br[39] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_42 
+ bl[40] br[40] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_43 
+ bl[41] br[41] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_44 
+ bl[42] br[42] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_45 
+ bl[43] br[43] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_46 
+ bl[44] br[44] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_47 
+ bl[45] br[45] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_48 
+ bl[46] br[46] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_49 
+ bl[47] br[47] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_50 
+ bl[48] br[48] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_51 
+ bl[49] br[49] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_52 
+ bl[50] br[50] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_53 
+ bl[51] br[51] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_54 
+ bl[52] br[52] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_55 
+ bl[53] br[53] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_56 
+ bl[54] br[54] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_57 
+ bl[55] br[55] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_58 
+ bl[56] br[56] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_59 
+ bl[57] br[57] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_60 
+ bl[58] br[58] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_61 
+ bl[59] br[59] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_62 
+ bl[60] br[60] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_63 
+ bl[61] br[61] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_64 
+ bl[62] br[62] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_65 
+ bl[63] br[63] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_66 
+ bl[64] br[64] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_67 
+ bl[65] br[65] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_68 
+ bl[66] br[66] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_69 
+ bl[67] br[67] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_70 
+ bl[68] br[68] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_71 
+ bl[69] br[69] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_72 
+ bl[70] br[70] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_73 
+ bl[71] br[71] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_74 
+ bl[72] br[72] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_75 
+ bl[73] br[73] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_76 
+ bl[74] br[74] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_77 
+ bl[75] br[75] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_78 
+ bl[76] br[76] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_79 
+ bl[77] br[77] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_80 
+ bl[78] br[78] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_81 
+ bl[79] br[79] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_82 
+ bl[80] br[80] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_83 
+ bl[81] br[81] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_84 
+ bl[82] br[82] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_85 
+ bl[83] br[83] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_86 
+ bl[84] br[84] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_87 
+ bl[85] br[85] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_88 
+ bl[86] br[86] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_89 
+ bl[87] br[87] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_90 
+ bl[88] br[88] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_91 
+ bl[89] br[89] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_92 
+ bl[90] br[90] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_93 
+ bl[91] br[91] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_94 
+ bl[92] br[92] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_95 
+ bl[93] br[93] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_96 
+ bl[94] br[94] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_97 
+ bl[95] br[95] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_98 
+ bl[96] br[96] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_99 
+ bl[97] br[97] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_100 
+ bl[98] br[98] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_101 
+ bl[99] br[99] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_102 
+ bl[100] br[100] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_103 
+ bl[101] br[101] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_104 
+ bl[102] br[102] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_105 
+ bl[103] br[103] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_106 
+ bl[104] br[104] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_107 
+ bl[105] br[105] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_108 
+ bl[106] br[106] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_109 
+ bl[107] br[107] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_110 
+ bl[108] br[108] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_111 
+ bl[109] br[109] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_112 
+ bl[110] br[110] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_113 
+ bl[111] br[111] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_114 
+ bl[112] br[112] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_115 
+ bl[113] br[113] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_116 
+ bl[114] br[114] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_117 
+ bl[115] br[115] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_118 
+ bl[116] br[116] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_119 
+ bl[117] br[117] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_120 
+ bl[118] br[118] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_121 
+ bl[119] br[119] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_122 
+ bl[120] br[120] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_123 
+ bl[121] br[121] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_124 
+ bl[122] br[122] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_125 
+ bl[123] br[123] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_126 
+ bl[124] br[124] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_127 
+ bl[125] br[125] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_128 
+ bl[126] br[126] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_129 
+ bl[127] br[127] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_130 
+ bl[128] br[128] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_131 
+ bl[129] br[129] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_132 
+ bl[130] br[130] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_133 
+ bl[131] br[131] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_134 
+ bl[132] br[132] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_135 
+ bl[133] br[133] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_136 
+ bl[134] br[134] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_137 
+ bl[135] br[135] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_138 
+ bl[136] br[136] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_139 
+ bl[137] br[137] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_140 
+ bl[138] br[138] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_141 
+ bl[139] br[139] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_142 
+ bl[140] br[140] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_143 
+ bl[141] br[141] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_144 
+ bl[142] br[142] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_145 
+ bl[143] br[143] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_146 
+ bl[144] br[144] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_147 
+ bl[145] br[145] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_148 
+ bl[146] br[146] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_149 
+ bl[147] br[147] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_150 
+ bl[148] br[148] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_151 
+ bl[149] br[149] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_152 
+ bl[150] br[150] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_153 
+ bl[151] br[151] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_154 
+ bl[152] br[152] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_155 
+ bl[153] br[153] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_156 
+ bl[154] br[154] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_157 
+ bl[155] br[155] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_158 
+ bl[156] br[156] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_159 
+ bl[157] br[157] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_160 
+ bl[158] br[158] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_161 
+ bl[159] br[159] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_162 
+ bl[160] br[160] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_163 
+ bl[161] br[161] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_164 
+ bl[162] br[162] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_165 
+ bl[163] br[163] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_166 
+ bl[164] br[164] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_167 
+ bl[165] br[165] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_168 
+ bl[166] br[166] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_169 
+ bl[167] br[167] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_170 
+ bl[168] br[168] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_171 
+ bl[169] br[169] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_172 
+ bl[170] br[170] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_173 
+ bl[171] br[171] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_174 
+ bl[172] br[172] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_175 
+ bl[173] br[173] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_176 
+ bl[174] br[174] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_177 
+ bl[175] br[175] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_178 
+ bl[176] br[176] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_179 
+ bl[177] br[177] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_180 
+ bl[178] br[178] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_181 
+ bl[179] br[179] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_182 
+ bl[180] br[180] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_183 
+ bl[181] br[181] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_184 
+ bl[182] br[182] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_185 
+ bl[183] br[183] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_186 
+ bl[184] br[184] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_187 
+ bl[185] br[185] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_188 
+ bl[186] br[186] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_189 
+ bl[187] br[187] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_190 
+ bl[188] br[188] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_191 
+ bl[189] br[189] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_192 
+ bl[190] br[190] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_193 
+ bl[191] br[191] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_194 
+ bl[192] br[192] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_195 
+ bl[193] br[193] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_196 
+ bl[194] br[194] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_197 
+ bl[195] br[195] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_198 
+ bl[196] br[196] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_199 
+ bl[197] br[197] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_200 
+ bl[198] br[198] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_201 
+ bl[199] br[199] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_202 
+ bl[200] br[200] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_203 
+ bl[201] br[201] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_204 
+ bl[202] br[202] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_205 
+ bl[203] br[203] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_206 
+ bl[204] br[204] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_207 
+ bl[205] br[205] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_208 
+ bl[206] br[206] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_209 
+ bl[207] br[207] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_210 
+ bl[208] br[208] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_211 
+ bl[209] br[209] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_212 
+ bl[210] br[210] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_213 
+ bl[211] br[211] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_214 
+ bl[212] br[212] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_215 
+ bl[213] br[213] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_216 
+ bl[214] br[214] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_217 
+ bl[215] br[215] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_218 
+ bl[216] br[216] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_219 
+ bl[217] br[217] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_220 
+ bl[218] br[218] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_221 
+ bl[219] br[219] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_222 
+ bl[220] br[220] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_223 
+ bl[221] br[221] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_224 
+ bl[222] br[222] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_225 
+ bl[223] br[223] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_226 
+ bl[224] br[224] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_227 
+ bl[225] br[225] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_228 
+ bl[226] br[226] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_229 
+ bl[227] br[227] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_230 
+ bl[228] br[228] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_231 
+ bl[229] br[229] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_232 
+ bl[230] br[230] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_233 
+ bl[231] br[231] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_234 
+ bl[232] br[232] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_235 
+ bl[233] br[233] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_236 
+ bl[234] br[234] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_237 
+ bl[235] br[235] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_238 
+ bl[236] br[236] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_239 
+ bl[237] br[237] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_240 
+ bl[238] br[238] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_241 
+ bl[239] br[239] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_242 
+ bl[240] br[240] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_243 
+ bl[241] br[241] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_244 
+ bl[242] br[242] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_245 
+ bl[243] br[243] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_246 
+ bl[244] br[244] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_247 
+ bl[245] br[245] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_248 
+ bl[246] br[246] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_249 
+ bl[247] br[247] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_250 
+ bl[248] br[248] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_251 
+ bl[249] br[249] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_252 
+ bl[250] br[250] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_253 
+ bl[251] br[251] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_254 
+ bl[252] br[252] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_255 
+ bl[253] br[253] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_256 
+ bl[254] br[254] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_257 
+ bl[255] br[255] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_258 
+ vdd vdd vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_259 
+ vdd vdd vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_0 
+ vdd vdd vss vdd vpb vnb wl[54] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_56_1 
+ rbl rbr vss vdd vpb vnb wl[54] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_56_2 
+ bl[0] br[0] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_3 
+ bl[1] br[1] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_4 
+ bl[2] br[2] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_5 
+ bl[3] br[3] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_6 
+ bl[4] br[4] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_7 
+ bl[5] br[5] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_8 
+ bl[6] br[6] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_9 
+ bl[7] br[7] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_10 
+ bl[8] br[8] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_11 
+ bl[9] br[9] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_12 
+ bl[10] br[10] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_13 
+ bl[11] br[11] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_14 
+ bl[12] br[12] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_15 
+ bl[13] br[13] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_16 
+ bl[14] br[14] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_17 
+ bl[15] br[15] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_18 
+ bl[16] br[16] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_19 
+ bl[17] br[17] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_20 
+ bl[18] br[18] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_21 
+ bl[19] br[19] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_22 
+ bl[20] br[20] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_23 
+ bl[21] br[21] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_24 
+ bl[22] br[22] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_25 
+ bl[23] br[23] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_26 
+ bl[24] br[24] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_27 
+ bl[25] br[25] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_28 
+ bl[26] br[26] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_29 
+ bl[27] br[27] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_30 
+ bl[28] br[28] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_31 
+ bl[29] br[29] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_32 
+ bl[30] br[30] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_33 
+ bl[31] br[31] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_34 
+ bl[32] br[32] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_35 
+ bl[33] br[33] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_36 
+ bl[34] br[34] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_37 
+ bl[35] br[35] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_38 
+ bl[36] br[36] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_39 
+ bl[37] br[37] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_40 
+ bl[38] br[38] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_41 
+ bl[39] br[39] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_42 
+ bl[40] br[40] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_43 
+ bl[41] br[41] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_44 
+ bl[42] br[42] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_45 
+ bl[43] br[43] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_46 
+ bl[44] br[44] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_47 
+ bl[45] br[45] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_48 
+ bl[46] br[46] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_49 
+ bl[47] br[47] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_50 
+ bl[48] br[48] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_51 
+ bl[49] br[49] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_52 
+ bl[50] br[50] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_53 
+ bl[51] br[51] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_54 
+ bl[52] br[52] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_55 
+ bl[53] br[53] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_56 
+ bl[54] br[54] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_57 
+ bl[55] br[55] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_58 
+ bl[56] br[56] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_59 
+ bl[57] br[57] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_60 
+ bl[58] br[58] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_61 
+ bl[59] br[59] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_62 
+ bl[60] br[60] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_63 
+ bl[61] br[61] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_64 
+ bl[62] br[62] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_65 
+ bl[63] br[63] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_66 
+ bl[64] br[64] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_67 
+ bl[65] br[65] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_68 
+ bl[66] br[66] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_69 
+ bl[67] br[67] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_70 
+ bl[68] br[68] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_71 
+ bl[69] br[69] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_72 
+ bl[70] br[70] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_73 
+ bl[71] br[71] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_74 
+ bl[72] br[72] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_75 
+ bl[73] br[73] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_76 
+ bl[74] br[74] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_77 
+ bl[75] br[75] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_78 
+ bl[76] br[76] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_79 
+ bl[77] br[77] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_80 
+ bl[78] br[78] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_81 
+ bl[79] br[79] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_82 
+ bl[80] br[80] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_83 
+ bl[81] br[81] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_84 
+ bl[82] br[82] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_85 
+ bl[83] br[83] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_86 
+ bl[84] br[84] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_87 
+ bl[85] br[85] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_88 
+ bl[86] br[86] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_89 
+ bl[87] br[87] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_90 
+ bl[88] br[88] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_91 
+ bl[89] br[89] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_92 
+ bl[90] br[90] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_93 
+ bl[91] br[91] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_94 
+ bl[92] br[92] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_95 
+ bl[93] br[93] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_96 
+ bl[94] br[94] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_97 
+ bl[95] br[95] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_98 
+ bl[96] br[96] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_99 
+ bl[97] br[97] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_100 
+ bl[98] br[98] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_101 
+ bl[99] br[99] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_102 
+ bl[100] br[100] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_103 
+ bl[101] br[101] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_104 
+ bl[102] br[102] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_105 
+ bl[103] br[103] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_106 
+ bl[104] br[104] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_107 
+ bl[105] br[105] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_108 
+ bl[106] br[106] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_109 
+ bl[107] br[107] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_110 
+ bl[108] br[108] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_111 
+ bl[109] br[109] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_112 
+ bl[110] br[110] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_113 
+ bl[111] br[111] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_114 
+ bl[112] br[112] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_115 
+ bl[113] br[113] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_116 
+ bl[114] br[114] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_117 
+ bl[115] br[115] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_118 
+ bl[116] br[116] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_119 
+ bl[117] br[117] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_120 
+ bl[118] br[118] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_121 
+ bl[119] br[119] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_122 
+ bl[120] br[120] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_123 
+ bl[121] br[121] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_124 
+ bl[122] br[122] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_125 
+ bl[123] br[123] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_126 
+ bl[124] br[124] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_127 
+ bl[125] br[125] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_128 
+ bl[126] br[126] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_129 
+ bl[127] br[127] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_130 
+ bl[128] br[128] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_131 
+ bl[129] br[129] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_132 
+ bl[130] br[130] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_133 
+ bl[131] br[131] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_134 
+ bl[132] br[132] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_135 
+ bl[133] br[133] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_136 
+ bl[134] br[134] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_137 
+ bl[135] br[135] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_138 
+ bl[136] br[136] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_139 
+ bl[137] br[137] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_140 
+ bl[138] br[138] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_141 
+ bl[139] br[139] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_142 
+ bl[140] br[140] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_143 
+ bl[141] br[141] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_144 
+ bl[142] br[142] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_145 
+ bl[143] br[143] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_146 
+ bl[144] br[144] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_147 
+ bl[145] br[145] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_148 
+ bl[146] br[146] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_149 
+ bl[147] br[147] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_150 
+ bl[148] br[148] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_151 
+ bl[149] br[149] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_152 
+ bl[150] br[150] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_153 
+ bl[151] br[151] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_154 
+ bl[152] br[152] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_155 
+ bl[153] br[153] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_156 
+ bl[154] br[154] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_157 
+ bl[155] br[155] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_158 
+ bl[156] br[156] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_159 
+ bl[157] br[157] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_160 
+ bl[158] br[158] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_161 
+ bl[159] br[159] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_162 
+ bl[160] br[160] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_163 
+ bl[161] br[161] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_164 
+ bl[162] br[162] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_165 
+ bl[163] br[163] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_166 
+ bl[164] br[164] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_167 
+ bl[165] br[165] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_168 
+ bl[166] br[166] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_169 
+ bl[167] br[167] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_170 
+ bl[168] br[168] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_171 
+ bl[169] br[169] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_172 
+ bl[170] br[170] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_173 
+ bl[171] br[171] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_174 
+ bl[172] br[172] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_175 
+ bl[173] br[173] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_176 
+ bl[174] br[174] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_177 
+ bl[175] br[175] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_178 
+ bl[176] br[176] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_179 
+ bl[177] br[177] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_180 
+ bl[178] br[178] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_181 
+ bl[179] br[179] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_182 
+ bl[180] br[180] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_183 
+ bl[181] br[181] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_184 
+ bl[182] br[182] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_185 
+ bl[183] br[183] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_186 
+ bl[184] br[184] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_187 
+ bl[185] br[185] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_188 
+ bl[186] br[186] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_189 
+ bl[187] br[187] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_190 
+ bl[188] br[188] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_191 
+ bl[189] br[189] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_192 
+ bl[190] br[190] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_193 
+ bl[191] br[191] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_194 
+ bl[192] br[192] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_195 
+ bl[193] br[193] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_196 
+ bl[194] br[194] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_197 
+ bl[195] br[195] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_198 
+ bl[196] br[196] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_199 
+ bl[197] br[197] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_200 
+ bl[198] br[198] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_201 
+ bl[199] br[199] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_202 
+ bl[200] br[200] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_203 
+ bl[201] br[201] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_204 
+ bl[202] br[202] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_205 
+ bl[203] br[203] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_206 
+ bl[204] br[204] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_207 
+ bl[205] br[205] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_208 
+ bl[206] br[206] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_209 
+ bl[207] br[207] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_210 
+ bl[208] br[208] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_211 
+ bl[209] br[209] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_212 
+ bl[210] br[210] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_213 
+ bl[211] br[211] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_214 
+ bl[212] br[212] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_215 
+ bl[213] br[213] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_216 
+ bl[214] br[214] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_217 
+ bl[215] br[215] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_218 
+ bl[216] br[216] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_219 
+ bl[217] br[217] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_220 
+ bl[218] br[218] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_221 
+ bl[219] br[219] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_222 
+ bl[220] br[220] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_223 
+ bl[221] br[221] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_224 
+ bl[222] br[222] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_225 
+ bl[223] br[223] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_226 
+ bl[224] br[224] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_227 
+ bl[225] br[225] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_228 
+ bl[226] br[226] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_229 
+ bl[227] br[227] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_230 
+ bl[228] br[228] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_231 
+ bl[229] br[229] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_232 
+ bl[230] br[230] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_233 
+ bl[231] br[231] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_234 
+ bl[232] br[232] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_235 
+ bl[233] br[233] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_236 
+ bl[234] br[234] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_237 
+ bl[235] br[235] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_238 
+ bl[236] br[236] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_239 
+ bl[237] br[237] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_240 
+ bl[238] br[238] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_241 
+ bl[239] br[239] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_242 
+ bl[240] br[240] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_243 
+ bl[241] br[241] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_244 
+ bl[242] br[242] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_245 
+ bl[243] br[243] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_246 
+ bl[244] br[244] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_247 
+ bl[245] br[245] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_248 
+ bl[246] br[246] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_249 
+ bl[247] br[247] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_250 
+ bl[248] br[248] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_251 
+ bl[249] br[249] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_252 
+ bl[250] br[250] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_253 
+ bl[251] br[251] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_254 
+ bl[252] br[252] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_255 
+ bl[253] br[253] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_256 
+ bl[254] br[254] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_257 
+ bl[255] br[255] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_258 
+ vdd vdd vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_259 
+ vdd vdd vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_0 
+ vdd vdd vss vdd vpb vnb wl[55] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_57_1 
+ rbl rbr vss vdd vpb vnb wl[55] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_57_2 
+ bl[0] br[0] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_3 
+ bl[1] br[1] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_4 
+ bl[2] br[2] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_5 
+ bl[3] br[3] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_6 
+ bl[4] br[4] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_7 
+ bl[5] br[5] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_8 
+ bl[6] br[6] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_9 
+ bl[7] br[7] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_10 
+ bl[8] br[8] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_11 
+ bl[9] br[9] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_12 
+ bl[10] br[10] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_13 
+ bl[11] br[11] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_14 
+ bl[12] br[12] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_15 
+ bl[13] br[13] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_16 
+ bl[14] br[14] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_17 
+ bl[15] br[15] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_18 
+ bl[16] br[16] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_19 
+ bl[17] br[17] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_20 
+ bl[18] br[18] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_21 
+ bl[19] br[19] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_22 
+ bl[20] br[20] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_23 
+ bl[21] br[21] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_24 
+ bl[22] br[22] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_25 
+ bl[23] br[23] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_26 
+ bl[24] br[24] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_27 
+ bl[25] br[25] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_28 
+ bl[26] br[26] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_29 
+ bl[27] br[27] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_30 
+ bl[28] br[28] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_31 
+ bl[29] br[29] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_32 
+ bl[30] br[30] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_33 
+ bl[31] br[31] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_34 
+ bl[32] br[32] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_35 
+ bl[33] br[33] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_36 
+ bl[34] br[34] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_37 
+ bl[35] br[35] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_38 
+ bl[36] br[36] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_39 
+ bl[37] br[37] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_40 
+ bl[38] br[38] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_41 
+ bl[39] br[39] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_42 
+ bl[40] br[40] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_43 
+ bl[41] br[41] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_44 
+ bl[42] br[42] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_45 
+ bl[43] br[43] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_46 
+ bl[44] br[44] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_47 
+ bl[45] br[45] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_48 
+ bl[46] br[46] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_49 
+ bl[47] br[47] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_50 
+ bl[48] br[48] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_51 
+ bl[49] br[49] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_52 
+ bl[50] br[50] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_53 
+ bl[51] br[51] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_54 
+ bl[52] br[52] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_55 
+ bl[53] br[53] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_56 
+ bl[54] br[54] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_57 
+ bl[55] br[55] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_58 
+ bl[56] br[56] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_59 
+ bl[57] br[57] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_60 
+ bl[58] br[58] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_61 
+ bl[59] br[59] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_62 
+ bl[60] br[60] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_63 
+ bl[61] br[61] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_64 
+ bl[62] br[62] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_65 
+ bl[63] br[63] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_66 
+ bl[64] br[64] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_67 
+ bl[65] br[65] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_68 
+ bl[66] br[66] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_69 
+ bl[67] br[67] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_70 
+ bl[68] br[68] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_71 
+ bl[69] br[69] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_72 
+ bl[70] br[70] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_73 
+ bl[71] br[71] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_74 
+ bl[72] br[72] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_75 
+ bl[73] br[73] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_76 
+ bl[74] br[74] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_77 
+ bl[75] br[75] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_78 
+ bl[76] br[76] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_79 
+ bl[77] br[77] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_80 
+ bl[78] br[78] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_81 
+ bl[79] br[79] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_82 
+ bl[80] br[80] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_83 
+ bl[81] br[81] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_84 
+ bl[82] br[82] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_85 
+ bl[83] br[83] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_86 
+ bl[84] br[84] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_87 
+ bl[85] br[85] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_88 
+ bl[86] br[86] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_89 
+ bl[87] br[87] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_90 
+ bl[88] br[88] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_91 
+ bl[89] br[89] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_92 
+ bl[90] br[90] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_93 
+ bl[91] br[91] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_94 
+ bl[92] br[92] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_95 
+ bl[93] br[93] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_96 
+ bl[94] br[94] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_97 
+ bl[95] br[95] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_98 
+ bl[96] br[96] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_99 
+ bl[97] br[97] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_100 
+ bl[98] br[98] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_101 
+ bl[99] br[99] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_102 
+ bl[100] br[100] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_103 
+ bl[101] br[101] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_104 
+ bl[102] br[102] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_105 
+ bl[103] br[103] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_106 
+ bl[104] br[104] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_107 
+ bl[105] br[105] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_108 
+ bl[106] br[106] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_109 
+ bl[107] br[107] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_110 
+ bl[108] br[108] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_111 
+ bl[109] br[109] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_112 
+ bl[110] br[110] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_113 
+ bl[111] br[111] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_114 
+ bl[112] br[112] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_115 
+ bl[113] br[113] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_116 
+ bl[114] br[114] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_117 
+ bl[115] br[115] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_118 
+ bl[116] br[116] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_119 
+ bl[117] br[117] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_120 
+ bl[118] br[118] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_121 
+ bl[119] br[119] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_122 
+ bl[120] br[120] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_123 
+ bl[121] br[121] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_124 
+ bl[122] br[122] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_125 
+ bl[123] br[123] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_126 
+ bl[124] br[124] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_127 
+ bl[125] br[125] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_128 
+ bl[126] br[126] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_129 
+ bl[127] br[127] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_130 
+ bl[128] br[128] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_131 
+ bl[129] br[129] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_132 
+ bl[130] br[130] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_133 
+ bl[131] br[131] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_134 
+ bl[132] br[132] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_135 
+ bl[133] br[133] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_136 
+ bl[134] br[134] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_137 
+ bl[135] br[135] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_138 
+ bl[136] br[136] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_139 
+ bl[137] br[137] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_140 
+ bl[138] br[138] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_141 
+ bl[139] br[139] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_142 
+ bl[140] br[140] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_143 
+ bl[141] br[141] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_144 
+ bl[142] br[142] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_145 
+ bl[143] br[143] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_146 
+ bl[144] br[144] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_147 
+ bl[145] br[145] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_148 
+ bl[146] br[146] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_149 
+ bl[147] br[147] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_150 
+ bl[148] br[148] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_151 
+ bl[149] br[149] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_152 
+ bl[150] br[150] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_153 
+ bl[151] br[151] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_154 
+ bl[152] br[152] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_155 
+ bl[153] br[153] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_156 
+ bl[154] br[154] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_157 
+ bl[155] br[155] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_158 
+ bl[156] br[156] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_159 
+ bl[157] br[157] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_160 
+ bl[158] br[158] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_161 
+ bl[159] br[159] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_162 
+ bl[160] br[160] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_163 
+ bl[161] br[161] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_164 
+ bl[162] br[162] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_165 
+ bl[163] br[163] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_166 
+ bl[164] br[164] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_167 
+ bl[165] br[165] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_168 
+ bl[166] br[166] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_169 
+ bl[167] br[167] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_170 
+ bl[168] br[168] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_171 
+ bl[169] br[169] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_172 
+ bl[170] br[170] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_173 
+ bl[171] br[171] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_174 
+ bl[172] br[172] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_175 
+ bl[173] br[173] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_176 
+ bl[174] br[174] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_177 
+ bl[175] br[175] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_178 
+ bl[176] br[176] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_179 
+ bl[177] br[177] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_180 
+ bl[178] br[178] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_181 
+ bl[179] br[179] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_182 
+ bl[180] br[180] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_183 
+ bl[181] br[181] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_184 
+ bl[182] br[182] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_185 
+ bl[183] br[183] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_186 
+ bl[184] br[184] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_187 
+ bl[185] br[185] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_188 
+ bl[186] br[186] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_189 
+ bl[187] br[187] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_190 
+ bl[188] br[188] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_191 
+ bl[189] br[189] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_192 
+ bl[190] br[190] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_193 
+ bl[191] br[191] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_194 
+ bl[192] br[192] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_195 
+ bl[193] br[193] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_196 
+ bl[194] br[194] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_197 
+ bl[195] br[195] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_198 
+ bl[196] br[196] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_199 
+ bl[197] br[197] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_200 
+ bl[198] br[198] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_201 
+ bl[199] br[199] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_202 
+ bl[200] br[200] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_203 
+ bl[201] br[201] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_204 
+ bl[202] br[202] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_205 
+ bl[203] br[203] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_206 
+ bl[204] br[204] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_207 
+ bl[205] br[205] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_208 
+ bl[206] br[206] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_209 
+ bl[207] br[207] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_210 
+ bl[208] br[208] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_211 
+ bl[209] br[209] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_212 
+ bl[210] br[210] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_213 
+ bl[211] br[211] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_214 
+ bl[212] br[212] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_215 
+ bl[213] br[213] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_216 
+ bl[214] br[214] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_217 
+ bl[215] br[215] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_218 
+ bl[216] br[216] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_219 
+ bl[217] br[217] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_220 
+ bl[218] br[218] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_221 
+ bl[219] br[219] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_222 
+ bl[220] br[220] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_223 
+ bl[221] br[221] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_224 
+ bl[222] br[222] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_225 
+ bl[223] br[223] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_226 
+ bl[224] br[224] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_227 
+ bl[225] br[225] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_228 
+ bl[226] br[226] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_229 
+ bl[227] br[227] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_230 
+ bl[228] br[228] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_231 
+ bl[229] br[229] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_232 
+ bl[230] br[230] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_233 
+ bl[231] br[231] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_234 
+ bl[232] br[232] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_235 
+ bl[233] br[233] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_236 
+ bl[234] br[234] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_237 
+ bl[235] br[235] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_238 
+ bl[236] br[236] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_239 
+ bl[237] br[237] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_240 
+ bl[238] br[238] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_241 
+ bl[239] br[239] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_242 
+ bl[240] br[240] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_243 
+ bl[241] br[241] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_244 
+ bl[242] br[242] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_245 
+ bl[243] br[243] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_246 
+ bl[244] br[244] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_247 
+ bl[245] br[245] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_248 
+ bl[246] br[246] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_249 
+ bl[247] br[247] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_250 
+ bl[248] br[248] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_251 
+ bl[249] br[249] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_252 
+ bl[250] br[250] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_253 
+ bl[251] br[251] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_254 
+ bl[252] br[252] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_255 
+ bl[253] br[253] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_256 
+ bl[254] br[254] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_257 
+ bl[255] br[255] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_258 
+ vdd vdd vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_259 
+ vdd vdd vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_0 
+ vdd vdd vss vdd vpb vnb wl[56] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_58_1 
+ rbl rbr vss vdd vpb vnb wl[56] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_58_2 
+ bl[0] br[0] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_3 
+ bl[1] br[1] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_4 
+ bl[2] br[2] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_5 
+ bl[3] br[3] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_6 
+ bl[4] br[4] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_7 
+ bl[5] br[5] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_8 
+ bl[6] br[6] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_9 
+ bl[7] br[7] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_10 
+ bl[8] br[8] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_11 
+ bl[9] br[9] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_12 
+ bl[10] br[10] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_13 
+ bl[11] br[11] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_14 
+ bl[12] br[12] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_15 
+ bl[13] br[13] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_16 
+ bl[14] br[14] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_17 
+ bl[15] br[15] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_18 
+ bl[16] br[16] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_19 
+ bl[17] br[17] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_20 
+ bl[18] br[18] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_21 
+ bl[19] br[19] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_22 
+ bl[20] br[20] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_23 
+ bl[21] br[21] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_24 
+ bl[22] br[22] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_25 
+ bl[23] br[23] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_26 
+ bl[24] br[24] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_27 
+ bl[25] br[25] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_28 
+ bl[26] br[26] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_29 
+ bl[27] br[27] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_30 
+ bl[28] br[28] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_31 
+ bl[29] br[29] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_32 
+ bl[30] br[30] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_33 
+ bl[31] br[31] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_34 
+ bl[32] br[32] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_35 
+ bl[33] br[33] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_36 
+ bl[34] br[34] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_37 
+ bl[35] br[35] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_38 
+ bl[36] br[36] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_39 
+ bl[37] br[37] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_40 
+ bl[38] br[38] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_41 
+ bl[39] br[39] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_42 
+ bl[40] br[40] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_43 
+ bl[41] br[41] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_44 
+ bl[42] br[42] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_45 
+ bl[43] br[43] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_46 
+ bl[44] br[44] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_47 
+ bl[45] br[45] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_48 
+ bl[46] br[46] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_49 
+ bl[47] br[47] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_50 
+ bl[48] br[48] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_51 
+ bl[49] br[49] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_52 
+ bl[50] br[50] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_53 
+ bl[51] br[51] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_54 
+ bl[52] br[52] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_55 
+ bl[53] br[53] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_56 
+ bl[54] br[54] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_57 
+ bl[55] br[55] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_58 
+ bl[56] br[56] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_59 
+ bl[57] br[57] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_60 
+ bl[58] br[58] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_61 
+ bl[59] br[59] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_62 
+ bl[60] br[60] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_63 
+ bl[61] br[61] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_64 
+ bl[62] br[62] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_65 
+ bl[63] br[63] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_66 
+ bl[64] br[64] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_67 
+ bl[65] br[65] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_68 
+ bl[66] br[66] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_69 
+ bl[67] br[67] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_70 
+ bl[68] br[68] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_71 
+ bl[69] br[69] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_72 
+ bl[70] br[70] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_73 
+ bl[71] br[71] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_74 
+ bl[72] br[72] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_75 
+ bl[73] br[73] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_76 
+ bl[74] br[74] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_77 
+ bl[75] br[75] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_78 
+ bl[76] br[76] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_79 
+ bl[77] br[77] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_80 
+ bl[78] br[78] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_81 
+ bl[79] br[79] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_82 
+ bl[80] br[80] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_83 
+ bl[81] br[81] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_84 
+ bl[82] br[82] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_85 
+ bl[83] br[83] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_86 
+ bl[84] br[84] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_87 
+ bl[85] br[85] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_88 
+ bl[86] br[86] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_89 
+ bl[87] br[87] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_90 
+ bl[88] br[88] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_91 
+ bl[89] br[89] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_92 
+ bl[90] br[90] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_93 
+ bl[91] br[91] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_94 
+ bl[92] br[92] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_95 
+ bl[93] br[93] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_96 
+ bl[94] br[94] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_97 
+ bl[95] br[95] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_98 
+ bl[96] br[96] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_99 
+ bl[97] br[97] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_100 
+ bl[98] br[98] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_101 
+ bl[99] br[99] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_102 
+ bl[100] br[100] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_103 
+ bl[101] br[101] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_104 
+ bl[102] br[102] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_105 
+ bl[103] br[103] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_106 
+ bl[104] br[104] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_107 
+ bl[105] br[105] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_108 
+ bl[106] br[106] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_109 
+ bl[107] br[107] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_110 
+ bl[108] br[108] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_111 
+ bl[109] br[109] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_112 
+ bl[110] br[110] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_113 
+ bl[111] br[111] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_114 
+ bl[112] br[112] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_115 
+ bl[113] br[113] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_116 
+ bl[114] br[114] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_117 
+ bl[115] br[115] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_118 
+ bl[116] br[116] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_119 
+ bl[117] br[117] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_120 
+ bl[118] br[118] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_121 
+ bl[119] br[119] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_122 
+ bl[120] br[120] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_123 
+ bl[121] br[121] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_124 
+ bl[122] br[122] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_125 
+ bl[123] br[123] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_126 
+ bl[124] br[124] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_127 
+ bl[125] br[125] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_128 
+ bl[126] br[126] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_129 
+ bl[127] br[127] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_130 
+ bl[128] br[128] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_131 
+ bl[129] br[129] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_132 
+ bl[130] br[130] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_133 
+ bl[131] br[131] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_134 
+ bl[132] br[132] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_135 
+ bl[133] br[133] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_136 
+ bl[134] br[134] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_137 
+ bl[135] br[135] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_138 
+ bl[136] br[136] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_139 
+ bl[137] br[137] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_140 
+ bl[138] br[138] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_141 
+ bl[139] br[139] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_142 
+ bl[140] br[140] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_143 
+ bl[141] br[141] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_144 
+ bl[142] br[142] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_145 
+ bl[143] br[143] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_146 
+ bl[144] br[144] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_147 
+ bl[145] br[145] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_148 
+ bl[146] br[146] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_149 
+ bl[147] br[147] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_150 
+ bl[148] br[148] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_151 
+ bl[149] br[149] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_152 
+ bl[150] br[150] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_153 
+ bl[151] br[151] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_154 
+ bl[152] br[152] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_155 
+ bl[153] br[153] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_156 
+ bl[154] br[154] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_157 
+ bl[155] br[155] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_158 
+ bl[156] br[156] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_159 
+ bl[157] br[157] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_160 
+ bl[158] br[158] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_161 
+ bl[159] br[159] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_162 
+ bl[160] br[160] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_163 
+ bl[161] br[161] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_164 
+ bl[162] br[162] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_165 
+ bl[163] br[163] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_166 
+ bl[164] br[164] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_167 
+ bl[165] br[165] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_168 
+ bl[166] br[166] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_169 
+ bl[167] br[167] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_170 
+ bl[168] br[168] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_171 
+ bl[169] br[169] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_172 
+ bl[170] br[170] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_173 
+ bl[171] br[171] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_174 
+ bl[172] br[172] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_175 
+ bl[173] br[173] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_176 
+ bl[174] br[174] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_177 
+ bl[175] br[175] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_178 
+ bl[176] br[176] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_179 
+ bl[177] br[177] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_180 
+ bl[178] br[178] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_181 
+ bl[179] br[179] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_182 
+ bl[180] br[180] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_183 
+ bl[181] br[181] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_184 
+ bl[182] br[182] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_185 
+ bl[183] br[183] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_186 
+ bl[184] br[184] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_187 
+ bl[185] br[185] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_188 
+ bl[186] br[186] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_189 
+ bl[187] br[187] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_190 
+ bl[188] br[188] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_191 
+ bl[189] br[189] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_192 
+ bl[190] br[190] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_193 
+ bl[191] br[191] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_194 
+ bl[192] br[192] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_195 
+ bl[193] br[193] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_196 
+ bl[194] br[194] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_197 
+ bl[195] br[195] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_198 
+ bl[196] br[196] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_199 
+ bl[197] br[197] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_200 
+ bl[198] br[198] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_201 
+ bl[199] br[199] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_202 
+ bl[200] br[200] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_203 
+ bl[201] br[201] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_204 
+ bl[202] br[202] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_205 
+ bl[203] br[203] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_206 
+ bl[204] br[204] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_207 
+ bl[205] br[205] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_208 
+ bl[206] br[206] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_209 
+ bl[207] br[207] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_210 
+ bl[208] br[208] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_211 
+ bl[209] br[209] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_212 
+ bl[210] br[210] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_213 
+ bl[211] br[211] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_214 
+ bl[212] br[212] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_215 
+ bl[213] br[213] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_216 
+ bl[214] br[214] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_217 
+ bl[215] br[215] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_218 
+ bl[216] br[216] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_219 
+ bl[217] br[217] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_220 
+ bl[218] br[218] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_221 
+ bl[219] br[219] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_222 
+ bl[220] br[220] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_223 
+ bl[221] br[221] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_224 
+ bl[222] br[222] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_225 
+ bl[223] br[223] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_226 
+ bl[224] br[224] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_227 
+ bl[225] br[225] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_228 
+ bl[226] br[226] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_229 
+ bl[227] br[227] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_230 
+ bl[228] br[228] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_231 
+ bl[229] br[229] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_232 
+ bl[230] br[230] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_233 
+ bl[231] br[231] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_234 
+ bl[232] br[232] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_235 
+ bl[233] br[233] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_236 
+ bl[234] br[234] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_237 
+ bl[235] br[235] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_238 
+ bl[236] br[236] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_239 
+ bl[237] br[237] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_240 
+ bl[238] br[238] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_241 
+ bl[239] br[239] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_242 
+ bl[240] br[240] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_243 
+ bl[241] br[241] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_244 
+ bl[242] br[242] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_245 
+ bl[243] br[243] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_246 
+ bl[244] br[244] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_247 
+ bl[245] br[245] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_248 
+ bl[246] br[246] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_249 
+ bl[247] br[247] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_250 
+ bl[248] br[248] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_251 
+ bl[249] br[249] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_252 
+ bl[250] br[250] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_253 
+ bl[251] br[251] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_254 
+ bl[252] br[252] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_255 
+ bl[253] br[253] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_256 
+ bl[254] br[254] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_257 
+ bl[255] br[255] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_258 
+ vdd vdd vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_259 
+ vdd vdd vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_0 
+ vdd vdd vss vdd vpb vnb wl[57] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_59_1 
+ rbl rbr vss vdd vpb vnb wl[57] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_59_2 
+ bl[0] br[0] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_3 
+ bl[1] br[1] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_4 
+ bl[2] br[2] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_5 
+ bl[3] br[3] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_6 
+ bl[4] br[4] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_7 
+ bl[5] br[5] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_8 
+ bl[6] br[6] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_9 
+ bl[7] br[7] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_10 
+ bl[8] br[8] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_11 
+ bl[9] br[9] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_12 
+ bl[10] br[10] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_13 
+ bl[11] br[11] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_14 
+ bl[12] br[12] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_15 
+ bl[13] br[13] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_16 
+ bl[14] br[14] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_17 
+ bl[15] br[15] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_18 
+ bl[16] br[16] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_19 
+ bl[17] br[17] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_20 
+ bl[18] br[18] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_21 
+ bl[19] br[19] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_22 
+ bl[20] br[20] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_23 
+ bl[21] br[21] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_24 
+ bl[22] br[22] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_25 
+ bl[23] br[23] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_26 
+ bl[24] br[24] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_27 
+ bl[25] br[25] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_28 
+ bl[26] br[26] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_29 
+ bl[27] br[27] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_30 
+ bl[28] br[28] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_31 
+ bl[29] br[29] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_32 
+ bl[30] br[30] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_33 
+ bl[31] br[31] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_34 
+ bl[32] br[32] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_35 
+ bl[33] br[33] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_36 
+ bl[34] br[34] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_37 
+ bl[35] br[35] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_38 
+ bl[36] br[36] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_39 
+ bl[37] br[37] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_40 
+ bl[38] br[38] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_41 
+ bl[39] br[39] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_42 
+ bl[40] br[40] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_43 
+ bl[41] br[41] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_44 
+ bl[42] br[42] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_45 
+ bl[43] br[43] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_46 
+ bl[44] br[44] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_47 
+ bl[45] br[45] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_48 
+ bl[46] br[46] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_49 
+ bl[47] br[47] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_50 
+ bl[48] br[48] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_51 
+ bl[49] br[49] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_52 
+ bl[50] br[50] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_53 
+ bl[51] br[51] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_54 
+ bl[52] br[52] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_55 
+ bl[53] br[53] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_56 
+ bl[54] br[54] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_57 
+ bl[55] br[55] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_58 
+ bl[56] br[56] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_59 
+ bl[57] br[57] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_60 
+ bl[58] br[58] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_61 
+ bl[59] br[59] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_62 
+ bl[60] br[60] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_63 
+ bl[61] br[61] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_64 
+ bl[62] br[62] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_65 
+ bl[63] br[63] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_66 
+ bl[64] br[64] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_67 
+ bl[65] br[65] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_68 
+ bl[66] br[66] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_69 
+ bl[67] br[67] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_70 
+ bl[68] br[68] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_71 
+ bl[69] br[69] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_72 
+ bl[70] br[70] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_73 
+ bl[71] br[71] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_74 
+ bl[72] br[72] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_75 
+ bl[73] br[73] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_76 
+ bl[74] br[74] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_77 
+ bl[75] br[75] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_78 
+ bl[76] br[76] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_79 
+ bl[77] br[77] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_80 
+ bl[78] br[78] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_81 
+ bl[79] br[79] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_82 
+ bl[80] br[80] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_83 
+ bl[81] br[81] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_84 
+ bl[82] br[82] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_85 
+ bl[83] br[83] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_86 
+ bl[84] br[84] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_87 
+ bl[85] br[85] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_88 
+ bl[86] br[86] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_89 
+ bl[87] br[87] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_90 
+ bl[88] br[88] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_91 
+ bl[89] br[89] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_92 
+ bl[90] br[90] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_93 
+ bl[91] br[91] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_94 
+ bl[92] br[92] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_95 
+ bl[93] br[93] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_96 
+ bl[94] br[94] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_97 
+ bl[95] br[95] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_98 
+ bl[96] br[96] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_99 
+ bl[97] br[97] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_100 
+ bl[98] br[98] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_101 
+ bl[99] br[99] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_102 
+ bl[100] br[100] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_103 
+ bl[101] br[101] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_104 
+ bl[102] br[102] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_105 
+ bl[103] br[103] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_106 
+ bl[104] br[104] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_107 
+ bl[105] br[105] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_108 
+ bl[106] br[106] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_109 
+ bl[107] br[107] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_110 
+ bl[108] br[108] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_111 
+ bl[109] br[109] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_112 
+ bl[110] br[110] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_113 
+ bl[111] br[111] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_114 
+ bl[112] br[112] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_115 
+ bl[113] br[113] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_116 
+ bl[114] br[114] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_117 
+ bl[115] br[115] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_118 
+ bl[116] br[116] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_119 
+ bl[117] br[117] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_120 
+ bl[118] br[118] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_121 
+ bl[119] br[119] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_122 
+ bl[120] br[120] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_123 
+ bl[121] br[121] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_124 
+ bl[122] br[122] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_125 
+ bl[123] br[123] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_126 
+ bl[124] br[124] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_127 
+ bl[125] br[125] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_128 
+ bl[126] br[126] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_129 
+ bl[127] br[127] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_130 
+ bl[128] br[128] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_131 
+ bl[129] br[129] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_132 
+ bl[130] br[130] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_133 
+ bl[131] br[131] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_134 
+ bl[132] br[132] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_135 
+ bl[133] br[133] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_136 
+ bl[134] br[134] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_137 
+ bl[135] br[135] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_138 
+ bl[136] br[136] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_139 
+ bl[137] br[137] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_140 
+ bl[138] br[138] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_141 
+ bl[139] br[139] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_142 
+ bl[140] br[140] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_143 
+ bl[141] br[141] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_144 
+ bl[142] br[142] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_145 
+ bl[143] br[143] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_146 
+ bl[144] br[144] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_147 
+ bl[145] br[145] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_148 
+ bl[146] br[146] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_149 
+ bl[147] br[147] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_150 
+ bl[148] br[148] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_151 
+ bl[149] br[149] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_152 
+ bl[150] br[150] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_153 
+ bl[151] br[151] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_154 
+ bl[152] br[152] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_155 
+ bl[153] br[153] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_156 
+ bl[154] br[154] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_157 
+ bl[155] br[155] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_158 
+ bl[156] br[156] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_159 
+ bl[157] br[157] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_160 
+ bl[158] br[158] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_161 
+ bl[159] br[159] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_162 
+ bl[160] br[160] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_163 
+ bl[161] br[161] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_164 
+ bl[162] br[162] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_165 
+ bl[163] br[163] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_166 
+ bl[164] br[164] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_167 
+ bl[165] br[165] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_168 
+ bl[166] br[166] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_169 
+ bl[167] br[167] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_170 
+ bl[168] br[168] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_171 
+ bl[169] br[169] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_172 
+ bl[170] br[170] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_173 
+ bl[171] br[171] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_174 
+ bl[172] br[172] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_175 
+ bl[173] br[173] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_176 
+ bl[174] br[174] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_177 
+ bl[175] br[175] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_178 
+ bl[176] br[176] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_179 
+ bl[177] br[177] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_180 
+ bl[178] br[178] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_181 
+ bl[179] br[179] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_182 
+ bl[180] br[180] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_183 
+ bl[181] br[181] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_184 
+ bl[182] br[182] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_185 
+ bl[183] br[183] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_186 
+ bl[184] br[184] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_187 
+ bl[185] br[185] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_188 
+ bl[186] br[186] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_189 
+ bl[187] br[187] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_190 
+ bl[188] br[188] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_191 
+ bl[189] br[189] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_192 
+ bl[190] br[190] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_193 
+ bl[191] br[191] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_194 
+ bl[192] br[192] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_195 
+ bl[193] br[193] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_196 
+ bl[194] br[194] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_197 
+ bl[195] br[195] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_198 
+ bl[196] br[196] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_199 
+ bl[197] br[197] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_200 
+ bl[198] br[198] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_201 
+ bl[199] br[199] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_202 
+ bl[200] br[200] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_203 
+ bl[201] br[201] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_204 
+ bl[202] br[202] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_205 
+ bl[203] br[203] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_206 
+ bl[204] br[204] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_207 
+ bl[205] br[205] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_208 
+ bl[206] br[206] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_209 
+ bl[207] br[207] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_210 
+ bl[208] br[208] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_211 
+ bl[209] br[209] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_212 
+ bl[210] br[210] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_213 
+ bl[211] br[211] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_214 
+ bl[212] br[212] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_215 
+ bl[213] br[213] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_216 
+ bl[214] br[214] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_217 
+ bl[215] br[215] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_218 
+ bl[216] br[216] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_219 
+ bl[217] br[217] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_220 
+ bl[218] br[218] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_221 
+ bl[219] br[219] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_222 
+ bl[220] br[220] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_223 
+ bl[221] br[221] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_224 
+ bl[222] br[222] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_225 
+ bl[223] br[223] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_226 
+ bl[224] br[224] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_227 
+ bl[225] br[225] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_228 
+ bl[226] br[226] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_229 
+ bl[227] br[227] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_230 
+ bl[228] br[228] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_231 
+ bl[229] br[229] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_232 
+ bl[230] br[230] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_233 
+ bl[231] br[231] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_234 
+ bl[232] br[232] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_235 
+ bl[233] br[233] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_236 
+ bl[234] br[234] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_237 
+ bl[235] br[235] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_238 
+ bl[236] br[236] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_239 
+ bl[237] br[237] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_240 
+ bl[238] br[238] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_241 
+ bl[239] br[239] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_242 
+ bl[240] br[240] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_243 
+ bl[241] br[241] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_244 
+ bl[242] br[242] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_245 
+ bl[243] br[243] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_246 
+ bl[244] br[244] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_247 
+ bl[245] br[245] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_248 
+ bl[246] br[246] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_249 
+ bl[247] br[247] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_250 
+ bl[248] br[248] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_251 
+ bl[249] br[249] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_252 
+ bl[250] br[250] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_253 
+ bl[251] br[251] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_254 
+ bl[252] br[252] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_255 
+ bl[253] br[253] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_256 
+ bl[254] br[254] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_257 
+ bl[255] br[255] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_258 
+ vdd vdd vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_259 
+ vdd vdd vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_0 
+ vdd vdd vss vdd vpb vnb wl[58] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_60_1 
+ rbl rbr vss vdd vpb vnb wl[58] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_60_2 
+ bl[0] br[0] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_3 
+ bl[1] br[1] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_4 
+ bl[2] br[2] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_5 
+ bl[3] br[3] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_6 
+ bl[4] br[4] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_7 
+ bl[5] br[5] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_8 
+ bl[6] br[6] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_9 
+ bl[7] br[7] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_10 
+ bl[8] br[8] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_11 
+ bl[9] br[9] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_12 
+ bl[10] br[10] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_13 
+ bl[11] br[11] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_14 
+ bl[12] br[12] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_15 
+ bl[13] br[13] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_16 
+ bl[14] br[14] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_17 
+ bl[15] br[15] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_18 
+ bl[16] br[16] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_19 
+ bl[17] br[17] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_20 
+ bl[18] br[18] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_21 
+ bl[19] br[19] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_22 
+ bl[20] br[20] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_23 
+ bl[21] br[21] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_24 
+ bl[22] br[22] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_25 
+ bl[23] br[23] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_26 
+ bl[24] br[24] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_27 
+ bl[25] br[25] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_28 
+ bl[26] br[26] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_29 
+ bl[27] br[27] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_30 
+ bl[28] br[28] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_31 
+ bl[29] br[29] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_32 
+ bl[30] br[30] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_33 
+ bl[31] br[31] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_34 
+ bl[32] br[32] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_35 
+ bl[33] br[33] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_36 
+ bl[34] br[34] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_37 
+ bl[35] br[35] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_38 
+ bl[36] br[36] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_39 
+ bl[37] br[37] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_40 
+ bl[38] br[38] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_41 
+ bl[39] br[39] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_42 
+ bl[40] br[40] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_43 
+ bl[41] br[41] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_44 
+ bl[42] br[42] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_45 
+ bl[43] br[43] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_46 
+ bl[44] br[44] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_47 
+ bl[45] br[45] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_48 
+ bl[46] br[46] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_49 
+ bl[47] br[47] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_50 
+ bl[48] br[48] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_51 
+ bl[49] br[49] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_52 
+ bl[50] br[50] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_53 
+ bl[51] br[51] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_54 
+ bl[52] br[52] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_55 
+ bl[53] br[53] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_56 
+ bl[54] br[54] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_57 
+ bl[55] br[55] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_58 
+ bl[56] br[56] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_59 
+ bl[57] br[57] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_60 
+ bl[58] br[58] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_61 
+ bl[59] br[59] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_62 
+ bl[60] br[60] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_63 
+ bl[61] br[61] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_64 
+ bl[62] br[62] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_65 
+ bl[63] br[63] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_66 
+ bl[64] br[64] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_67 
+ bl[65] br[65] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_68 
+ bl[66] br[66] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_69 
+ bl[67] br[67] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_70 
+ bl[68] br[68] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_71 
+ bl[69] br[69] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_72 
+ bl[70] br[70] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_73 
+ bl[71] br[71] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_74 
+ bl[72] br[72] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_75 
+ bl[73] br[73] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_76 
+ bl[74] br[74] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_77 
+ bl[75] br[75] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_78 
+ bl[76] br[76] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_79 
+ bl[77] br[77] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_80 
+ bl[78] br[78] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_81 
+ bl[79] br[79] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_82 
+ bl[80] br[80] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_83 
+ bl[81] br[81] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_84 
+ bl[82] br[82] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_85 
+ bl[83] br[83] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_86 
+ bl[84] br[84] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_87 
+ bl[85] br[85] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_88 
+ bl[86] br[86] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_89 
+ bl[87] br[87] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_90 
+ bl[88] br[88] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_91 
+ bl[89] br[89] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_92 
+ bl[90] br[90] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_93 
+ bl[91] br[91] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_94 
+ bl[92] br[92] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_95 
+ bl[93] br[93] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_96 
+ bl[94] br[94] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_97 
+ bl[95] br[95] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_98 
+ bl[96] br[96] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_99 
+ bl[97] br[97] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_100 
+ bl[98] br[98] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_101 
+ bl[99] br[99] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_102 
+ bl[100] br[100] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_103 
+ bl[101] br[101] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_104 
+ bl[102] br[102] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_105 
+ bl[103] br[103] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_106 
+ bl[104] br[104] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_107 
+ bl[105] br[105] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_108 
+ bl[106] br[106] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_109 
+ bl[107] br[107] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_110 
+ bl[108] br[108] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_111 
+ bl[109] br[109] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_112 
+ bl[110] br[110] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_113 
+ bl[111] br[111] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_114 
+ bl[112] br[112] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_115 
+ bl[113] br[113] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_116 
+ bl[114] br[114] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_117 
+ bl[115] br[115] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_118 
+ bl[116] br[116] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_119 
+ bl[117] br[117] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_120 
+ bl[118] br[118] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_121 
+ bl[119] br[119] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_122 
+ bl[120] br[120] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_123 
+ bl[121] br[121] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_124 
+ bl[122] br[122] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_125 
+ bl[123] br[123] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_126 
+ bl[124] br[124] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_127 
+ bl[125] br[125] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_128 
+ bl[126] br[126] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_129 
+ bl[127] br[127] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_130 
+ bl[128] br[128] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_131 
+ bl[129] br[129] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_132 
+ bl[130] br[130] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_133 
+ bl[131] br[131] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_134 
+ bl[132] br[132] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_135 
+ bl[133] br[133] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_136 
+ bl[134] br[134] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_137 
+ bl[135] br[135] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_138 
+ bl[136] br[136] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_139 
+ bl[137] br[137] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_140 
+ bl[138] br[138] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_141 
+ bl[139] br[139] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_142 
+ bl[140] br[140] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_143 
+ bl[141] br[141] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_144 
+ bl[142] br[142] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_145 
+ bl[143] br[143] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_146 
+ bl[144] br[144] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_147 
+ bl[145] br[145] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_148 
+ bl[146] br[146] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_149 
+ bl[147] br[147] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_150 
+ bl[148] br[148] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_151 
+ bl[149] br[149] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_152 
+ bl[150] br[150] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_153 
+ bl[151] br[151] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_154 
+ bl[152] br[152] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_155 
+ bl[153] br[153] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_156 
+ bl[154] br[154] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_157 
+ bl[155] br[155] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_158 
+ bl[156] br[156] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_159 
+ bl[157] br[157] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_160 
+ bl[158] br[158] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_161 
+ bl[159] br[159] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_162 
+ bl[160] br[160] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_163 
+ bl[161] br[161] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_164 
+ bl[162] br[162] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_165 
+ bl[163] br[163] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_166 
+ bl[164] br[164] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_167 
+ bl[165] br[165] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_168 
+ bl[166] br[166] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_169 
+ bl[167] br[167] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_170 
+ bl[168] br[168] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_171 
+ bl[169] br[169] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_172 
+ bl[170] br[170] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_173 
+ bl[171] br[171] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_174 
+ bl[172] br[172] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_175 
+ bl[173] br[173] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_176 
+ bl[174] br[174] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_177 
+ bl[175] br[175] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_178 
+ bl[176] br[176] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_179 
+ bl[177] br[177] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_180 
+ bl[178] br[178] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_181 
+ bl[179] br[179] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_182 
+ bl[180] br[180] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_183 
+ bl[181] br[181] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_184 
+ bl[182] br[182] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_185 
+ bl[183] br[183] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_186 
+ bl[184] br[184] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_187 
+ bl[185] br[185] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_188 
+ bl[186] br[186] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_189 
+ bl[187] br[187] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_190 
+ bl[188] br[188] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_191 
+ bl[189] br[189] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_192 
+ bl[190] br[190] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_193 
+ bl[191] br[191] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_194 
+ bl[192] br[192] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_195 
+ bl[193] br[193] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_196 
+ bl[194] br[194] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_197 
+ bl[195] br[195] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_198 
+ bl[196] br[196] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_199 
+ bl[197] br[197] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_200 
+ bl[198] br[198] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_201 
+ bl[199] br[199] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_202 
+ bl[200] br[200] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_203 
+ bl[201] br[201] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_204 
+ bl[202] br[202] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_205 
+ bl[203] br[203] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_206 
+ bl[204] br[204] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_207 
+ bl[205] br[205] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_208 
+ bl[206] br[206] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_209 
+ bl[207] br[207] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_210 
+ bl[208] br[208] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_211 
+ bl[209] br[209] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_212 
+ bl[210] br[210] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_213 
+ bl[211] br[211] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_214 
+ bl[212] br[212] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_215 
+ bl[213] br[213] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_216 
+ bl[214] br[214] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_217 
+ bl[215] br[215] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_218 
+ bl[216] br[216] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_219 
+ bl[217] br[217] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_220 
+ bl[218] br[218] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_221 
+ bl[219] br[219] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_222 
+ bl[220] br[220] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_223 
+ bl[221] br[221] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_224 
+ bl[222] br[222] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_225 
+ bl[223] br[223] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_226 
+ bl[224] br[224] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_227 
+ bl[225] br[225] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_228 
+ bl[226] br[226] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_229 
+ bl[227] br[227] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_230 
+ bl[228] br[228] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_231 
+ bl[229] br[229] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_232 
+ bl[230] br[230] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_233 
+ bl[231] br[231] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_234 
+ bl[232] br[232] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_235 
+ bl[233] br[233] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_236 
+ bl[234] br[234] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_237 
+ bl[235] br[235] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_238 
+ bl[236] br[236] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_239 
+ bl[237] br[237] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_240 
+ bl[238] br[238] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_241 
+ bl[239] br[239] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_242 
+ bl[240] br[240] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_243 
+ bl[241] br[241] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_244 
+ bl[242] br[242] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_245 
+ bl[243] br[243] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_246 
+ bl[244] br[244] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_247 
+ bl[245] br[245] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_248 
+ bl[246] br[246] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_249 
+ bl[247] br[247] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_250 
+ bl[248] br[248] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_251 
+ bl[249] br[249] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_252 
+ bl[250] br[250] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_253 
+ bl[251] br[251] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_254 
+ bl[252] br[252] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_255 
+ bl[253] br[253] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_256 
+ bl[254] br[254] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_257 
+ bl[255] br[255] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_258 
+ vdd vdd vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_259 
+ vdd vdd vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_0 
+ vdd vdd vss vdd vpb vnb wl[59] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_61_1 
+ rbl rbr vss vdd vpb vnb wl[59] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_61_2 
+ bl[0] br[0] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_3 
+ bl[1] br[1] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_4 
+ bl[2] br[2] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_5 
+ bl[3] br[3] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_6 
+ bl[4] br[4] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_7 
+ bl[5] br[5] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_8 
+ bl[6] br[6] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_9 
+ bl[7] br[7] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_10 
+ bl[8] br[8] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_11 
+ bl[9] br[9] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_12 
+ bl[10] br[10] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_13 
+ bl[11] br[11] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_14 
+ bl[12] br[12] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_15 
+ bl[13] br[13] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_16 
+ bl[14] br[14] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_17 
+ bl[15] br[15] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_18 
+ bl[16] br[16] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_19 
+ bl[17] br[17] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_20 
+ bl[18] br[18] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_21 
+ bl[19] br[19] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_22 
+ bl[20] br[20] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_23 
+ bl[21] br[21] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_24 
+ bl[22] br[22] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_25 
+ bl[23] br[23] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_26 
+ bl[24] br[24] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_27 
+ bl[25] br[25] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_28 
+ bl[26] br[26] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_29 
+ bl[27] br[27] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_30 
+ bl[28] br[28] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_31 
+ bl[29] br[29] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_32 
+ bl[30] br[30] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_33 
+ bl[31] br[31] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_34 
+ bl[32] br[32] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_35 
+ bl[33] br[33] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_36 
+ bl[34] br[34] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_37 
+ bl[35] br[35] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_38 
+ bl[36] br[36] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_39 
+ bl[37] br[37] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_40 
+ bl[38] br[38] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_41 
+ bl[39] br[39] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_42 
+ bl[40] br[40] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_43 
+ bl[41] br[41] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_44 
+ bl[42] br[42] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_45 
+ bl[43] br[43] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_46 
+ bl[44] br[44] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_47 
+ bl[45] br[45] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_48 
+ bl[46] br[46] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_49 
+ bl[47] br[47] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_50 
+ bl[48] br[48] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_51 
+ bl[49] br[49] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_52 
+ bl[50] br[50] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_53 
+ bl[51] br[51] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_54 
+ bl[52] br[52] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_55 
+ bl[53] br[53] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_56 
+ bl[54] br[54] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_57 
+ bl[55] br[55] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_58 
+ bl[56] br[56] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_59 
+ bl[57] br[57] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_60 
+ bl[58] br[58] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_61 
+ bl[59] br[59] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_62 
+ bl[60] br[60] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_63 
+ bl[61] br[61] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_64 
+ bl[62] br[62] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_65 
+ bl[63] br[63] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_66 
+ bl[64] br[64] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_67 
+ bl[65] br[65] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_68 
+ bl[66] br[66] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_69 
+ bl[67] br[67] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_70 
+ bl[68] br[68] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_71 
+ bl[69] br[69] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_72 
+ bl[70] br[70] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_73 
+ bl[71] br[71] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_74 
+ bl[72] br[72] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_75 
+ bl[73] br[73] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_76 
+ bl[74] br[74] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_77 
+ bl[75] br[75] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_78 
+ bl[76] br[76] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_79 
+ bl[77] br[77] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_80 
+ bl[78] br[78] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_81 
+ bl[79] br[79] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_82 
+ bl[80] br[80] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_83 
+ bl[81] br[81] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_84 
+ bl[82] br[82] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_85 
+ bl[83] br[83] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_86 
+ bl[84] br[84] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_87 
+ bl[85] br[85] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_88 
+ bl[86] br[86] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_89 
+ bl[87] br[87] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_90 
+ bl[88] br[88] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_91 
+ bl[89] br[89] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_92 
+ bl[90] br[90] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_93 
+ bl[91] br[91] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_94 
+ bl[92] br[92] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_95 
+ bl[93] br[93] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_96 
+ bl[94] br[94] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_97 
+ bl[95] br[95] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_98 
+ bl[96] br[96] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_99 
+ bl[97] br[97] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_100 
+ bl[98] br[98] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_101 
+ bl[99] br[99] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_102 
+ bl[100] br[100] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_103 
+ bl[101] br[101] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_104 
+ bl[102] br[102] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_105 
+ bl[103] br[103] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_106 
+ bl[104] br[104] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_107 
+ bl[105] br[105] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_108 
+ bl[106] br[106] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_109 
+ bl[107] br[107] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_110 
+ bl[108] br[108] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_111 
+ bl[109] br[109] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_112 
+ bl[110] br[110] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_113 
+ bl[111] br[111] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_114 
+ bl[112] br[112] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_115 
+ bl[113] br[113] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_116 
+ bl[114] br[114] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_117 
+ bl[115] br[115] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_118 
+ bl[116] br[116] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_119 
+ bl[117] br[117] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_120 
+ bl[118] br[118] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_121 
+ bl[119] br[119] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_122 
+ bl[120] br[120] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_123 
+ bl[121] br[121] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_124 
+ bl[122] br[122] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_125 
+ bl[123] br[123] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_126 
+ bl[124] br[124] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_127 
+ bl[125] br[125] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_128 
+ bl[126] br[126] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_129 
+ bl[127] br[127] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_130 
+ bl[128] br[128] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_131 
+ bl[129] br[129] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_132 
+ bl[130] br[130] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_133 
+ bl[131] br[131] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_134 
+ bl[132] br[132] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_135 
+ bl[133] br[133] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_136 
+ bl[134] br[134] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_137 
+ bl[135] br[135] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_138 
+ bl[136] br[136] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_139 
+ bl[137] br[137] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_140 
+ bl[138] br[138] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_141 
+ bl[139] br[139] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_142 
+ bl[140] br[140] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_143 
+ bl[141] br[141] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_144 
+ bl[142] br[142] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_145 
+ bl[143] br[143] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_146 
+ bl[144] br[144] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_147 
+ bl[145] br[145] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_148 
+ bl[146] br[146] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_149 
+ bl[147] br[147] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_150 
+ bl[148] br[148] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_151 
+ bl[149] br[149] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_152 
+ bl[150] br[150] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_153 
+ bl[151] br[151] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_154 
+ bl[152] br[152] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_155 
+ bl[153] br[153] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_156 
+ bl[154] br[154] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_157 
+ bl[155] br[155] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_158 
+ bl[156] br[156] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_159 
+ bl[157] br[157] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_160 
+ bl[158] br[158] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_161 
+ bl[159] br[159] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_162 
+ bl[160] br[160] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_163 
+ bl[161] br[161] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_164 
+ bl[162] br[162] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_165 
+ bl[163] br[163] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_166 
+ bl[164] br[164] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_167 
+ bl[165] br[165] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_168 
+ bl[166] br[166] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_169 
+ bl[167] br[167] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_170 
+ bl[168] br[168] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_171 
+ bl[169] br[169] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_172 
+ bl[170] br[170] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_173 
+ bl[171] br[171] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_174 
+ bl[172] br[172] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_175 
+ bl[173] br[173] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_176 
+ bl[174] br[174] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_177 
+ bl[175] br[175] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_178 
+ bl[176] br[176] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_179 
+ bl[177] br[177] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_180 
+ bl[178] br[178] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_181 
+ bl[179] br[179] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_182 
+ bl[180] br[180] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_183 
+ bl[181] br[181] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_184 
+ bl[182] br[182] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_185 
+ bl[183] br[183] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_186 
+ bl[184] br[184] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_187 
+ bl[185] br[185] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_188 
+ bl[186] br[186] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_189 
+ bl[187] br[187] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_190 
+ bl[188] br[188] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_191 
+ bl[189] br[189] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_192 
+ bl[190] br[190] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_193 
+ bl[191] br[191] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_194 
+ bl[192] br[192] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_195 
+ bl[193] br[193] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_196 
+ bl[194] br[194] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_197 
+ bl[195] br[195] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_198 
+ bl[196] br[196] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_199 
+ bl[197] br[197] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_200 
+ bl[198] br[198] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_201 
+ bl[199] br[199] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_202 
+ bl[200] br[200] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_203 
+ bl[201] br[201] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_204 
+ bl[202] br[202] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_205 
+ bl[203] br[203] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_206 
+ bl[204] br[204] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_207 
+ bl[205] br[205] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_208 
+ bl[206] br[206] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_209 
+ bl[207] br[207] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_210 
+ bl[208] br[208] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_211 
+ bl[209] br[209] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_212 
+ bl[210] br[210] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_213 
+ bl[211] br[211] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_214 
+ bl[212] br[212] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_215 
+ bl[213] br[213] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_216 
+ bl[214] br[214] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_217 
+ bl[215] br[215] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_218 
+ bl[216] br[216] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_219 
+ bl[217] br[217] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_220 
+ bl[218] br[218] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_221 
+ bl[219] br[219] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_222 
+ bl[220] br[220] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_223 
+ bl[221] br[221] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_224 
+ bl[222] br[222] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_225 
+ bl[223] br[223] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_226 
+ bl[224] br[224] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_227 
+ bl[225] br[225] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_228 
+ bl[226] br[226] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_229 
+ bl[227] br[227] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_230 
+ bl[228] br[228] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_231 
+ bl[229] br[229] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_232 
+ bl[230] br[230] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_233 
+ bl[231] br[231] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_234 
+ bl[232] br[232] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_235 
+ bl[233] br[233] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_236 
+ bl[234] br[234] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_237 
+ bl[235] br[235] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_238 
+ bl[236] br[236] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_239 
+ bl[237] br[237] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_240 
+ bl[238] br[238] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_241 
+ bl[239] br[239] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_242 
+ bl[240] br[240] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_243 
+ bl[241] br[241] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_244 
+ bl[242] br[242] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_245 
+ bl[243] br[243] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_246 
+ bl[244] br[244] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_247 
+ bl[245] br[245] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_248 
+ bl[246] br[246] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_249 
+ bl[247] br[247] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_250 
+ bl[248] br[248] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_251 
+ bl[249] br[249] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_252 
+ bl[250] br[250] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_253 
+ bl[251] br[251] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_254 
+ bl[252] br[252] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_255 
+ bl[253] br[253] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_256 
+ bl[254] br[254] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_257 
+ bl[255] br[255] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_258 
+ vdd vdd vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_259 
+ vdd vdd vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_0 
+ vdd vdd vss vdd vpb vnb wl[60] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_62_1 
+ rbl rbr vss vdd vpb vnb wl[60] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_62_2 
+ bl[0] br[0] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_3 
+ bl[1] br[1] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_4 
+ bl[2] br[2] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_5 
+ bl[3] br[3] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_6 
+ bl[4] br[4] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_7 
+ bl[5] br[5] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_8 
+ bl[6] br[6] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_9 
+ bl[7] br[7] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_10 
+ bl[8] br[8] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_11 
+ bl[9] br[9] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_12 
+ bl[10] br[10] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_13 
+ bl[11] br[11] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_14 
+ bl[12] br[12] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_15 
+ bl[13] br[13] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_16 
+ bl[14] br[14] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_17 
+ bl[15] br[15] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_18 
+ bl[16] br[16] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_19 
+ bl[17] br[17] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_20 
+ bl[18] br[18] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_21 
+ bl[19] br[19] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_22 
+ bl[20] br[20] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_23 
+ bl[21] br[21] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_24 
+ bl[22] br[22] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_25 
+ bl[23] br[23] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_26 
+ bl[24] br[24] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_27 
+ bl[25] br[25] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_28 
+ bl[26] br[26] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_29 
+ bl[27] br[27] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_30 
+ bl[28] br[28] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_31 
+ bl[29] br[29] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_32 
+ bl[30] br[30] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_33 
+ bl[31] br[31] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_34 
+ bl[32] br[32] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_35 
+ bl[33] br[33] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_36 
+ bl[34] br[34] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_37 
+ bl[35] br[35] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_38 
+ bl[36] br[36] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_39 
+ bl[37] br[37] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_40 
+ bl[38] br[38] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_41 
+ bl[39] br[39] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_42 
+ bl[40] br[40] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_43 
+ bl[41] br[41] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_44 
+ bl[42] br[42] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_45 
+ bl[43] br[43] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_46 
+ bl[44] br[44] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_47 
+ bl[45] br[45] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_48 
+ bl[46] br[46] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_49 
+ bl[47] br[47] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_50 
+ bl[48] br[48] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_51 
+ bl[49] br[49] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_52 
+ bl[50] br[50] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_53 
+ bl[51] br[51] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_54 
+ bl[52] br[52] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_55 
+ bl[53] br[53] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_56 
+ bl[54] br[54] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_57 
+ bl[55] br[55] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_58 
+ bl[56] br[56] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_59 
+ bl[57] br[57] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_60 
+ bl[58] br[58] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_61 
+ bl[59] br[59] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_62 
+ bl[60] br[60] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_63 
+ bl[61] br[61] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_64 
+ bl[62] br[62] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_65 
+ bl[63] br[63] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_66 
+ bl[64] br[64] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_67 
+ bl[65] br[65] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_68 
+ bl[66] br[66] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_69 
+ bl[67] br[67] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_70 
+ bl[68] br[68] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_71 
+ bl[69] br[69] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_72 
+ bl[70] br[70] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_73 
+ bl[71] br[71] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_74 
+ bl[72] br[72] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_75 
+ bl[73] br[73] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_76 
+ bl[74] br[74] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_77 
+ bl[75] br[75] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_78 
+ bl[76] br[76] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_79 
+ bl[77] br[77] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_80 
+ bl[78] br[78] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_81 
+ bl[79] br[79] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_82 
+ bl[80] br[80] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_83 
+ bl[81] br[81] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_84 
+ bl[82] br[82] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_85 
+ bl[83] br[83] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_86 
+ bl[84] br[84] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_87 
+ bl[85] br[85] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_88 
+ bl[86] br[86] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_89 
+ bl[87] br[87] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_90 
+ bl[88] br[88] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_91 
+ bl[89] br[89] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_92 
+ bl[90] br[90] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_93 
+ bl[91] br[91] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_94 
+ bl[92] br[92] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_95 
+ bl[93] br[93] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_96 
+ bl[94] br[94] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_97 
+ bl[95] br[95] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_98 
+ bl[96] br[96] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_99 
+ bl[97] br[97] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_100 
+ bl[98] br[98] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_101 
+ bl[99] br[99] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_102 
+ bl[100] br[100] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_103 
+ bl[101] br[101] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_104 
+ bl[102] br[102] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_105 
+ bl[103] br[103] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_106 
+ bl[104] br[104] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_107 
+ bl[105] br[105] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_108 
+ bl[106] br[106] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_109 
+ bl[107] br[107] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_110 
+ bl[108] br[108] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_111 
+ bl[109] br[109] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_112 
+ bl[110] br[110] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_113 
+ bl[111] br[111] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_114 
+ bl[112] br[112] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_115 
+ bl[113] br[113] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_116 
+ bl[114] br[114] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_117 
+ bl[115] br[115] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_118 
+ bl[116] br[116] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_119 
+ bl[117] br[117] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_120 
+ bl[118] br[118] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_121 
+ bl[119] br[119] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_122 
+ bl[120] br[120] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_123 
+ bl[121] br[121] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_124 
+ bl[122] br[122] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_125 
+ bl[123] br[123] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_126 
+ bl[124] br[124] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_127 
+ bl[125] br[125] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_128 
+ bl[126] br[126] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_129 
+ bl[127] br[127] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_130 
+ bl[128] br[128] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_131 
+ bl[129] br[129] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_132 
+ bl[130] br[130] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_133 
+ bl[131] br[131] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_134 
+ bl[132] br[132] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_135 
+ bl[133] br[133] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_136 
+ bl[134] br[134] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_137 
+ bl[135] br[135] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_138 
+ bl[136] br[136] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_139 
+ bl[137] br[137] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_140 
+ bl[138] br[138] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_141 
+ bl[139] br[139] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_142 
+ bl[140] br[140] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_143 
+ bl[141] br[141] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_144 
+ bl[142] br[142] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_145 
+ bl[143] br[143] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_146 
+ bl[144] br[144] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_147 
+ bl[145] br[145] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_148 
+ bl[146] br[146] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_149 
+ bl[147] br[147] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_150 
+ bl[148] br[148] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_151 
+ bl[149] br[149] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_152 
+ bl[150] br[150] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_153 
+ bl[151] br[151] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_154 
+ bl[152] br[152] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_155 
+ bl[153] br[153] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_156 
+ bl[154] br[154] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_157 
+ bl[155] br[155] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_158 
+ bl[156] br[156] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_159 
+ bl[157] br[157] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_160 
+ bl[158] br[158] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_161 
+ bl[159] br[159] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_162 
+ bl[160] br[160] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_163 
+ bl[161] br[161] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_164 
+ bl[162] br[162] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_165 
+ bl[163] br[163] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_166 
+ bl[164] br[164] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_167 
+ bl[165] br[165] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_168 
+ bl[166] br[166] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_169 
+ bl[167] br[167] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_170 
+ bl[168] br[168] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_171 
+ bl[169] br[169] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_172 
+ bl[170] br[170] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_173 
+ bl[171] br[171] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_174 
+ bl[172] br[172] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_175 
+ bl[173] br[173] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_176 
+ bl[174] br[174] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_177 
+ bl[175] br[175] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_178 
+ bl[176] br[176] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_179 
+ bl[177] br[177] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_180 
+ bl[178] br[178] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_181 
+ bl[179] br[179] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_182 
+ bl[180] br[180] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_183 
+ bl[181] br[181] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_184 
+ bl[182] br[182] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_185 
+ bl[183] br[183] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_186 
+ bl[184] br[184] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_187 
+ bl[185] br[185] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_188 
+ bl[186] br[186] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_189 
+ bl[187] br[187] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_190 
+ bl[188] br[188] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_191 
+ bl[189] br[189] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_192 
+ bl[190] br[190] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_193 
+ bl[191] br[191] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_194 
+ bl[192] br[192] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_195 
+ bl[193] br[193] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_196 
+ bl[194] br[194] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_197 
+ bl[195] br[195] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_198 
+ bl[196] br[196] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_199 
+ bl[197] br[197] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_200 
+ bl[198] br[198] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_201 
+ bl[199] br[199] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_202 
+ bl[200] br[200] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_203 
+ bl[201] br[201] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_204 
+ bl[202] br[202] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_205 
+ bl[203] br[203] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_206 
+ bl[204] br[204] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_207 
+ bl[205] br[205] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_208 
+ bl[206] br[206] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_209 
+ bl[207] br[207] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_210 
+ bl[208] br[208] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_211 
+ bl[209] br[209] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_212 
+ bl[210] br[210] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_213 
+ bl[211] br[211] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_214 
+ bl[212] br[212] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_215 
+ bl[213] br[213] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_216 
+ bl[214] br[214] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_217 
+ bl[215] br[215] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_218 
+ bl[216] br[216] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_219 
+ bl[217] br[217] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_220 
+ bl[218] br[218] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_221 
+ bl[219] br[219] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_222 
+ bl[220] br[220] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_223 
+ bl[221] br[221] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_224 
+ bl[222] br[222] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_225 
+ bl[223] br[223] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_226 
+ bl[224] br[224] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_227 
+ bl[225] br[225] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_228 
+ bl[226] br[226] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_229 
+ bl[227] br[227] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_230 
+ bl[228] br[228] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_231 
+ bl[229] br[229] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_232 
+ bl[230] br[230] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_233 
+ bl[231] br[231] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_234 
+ bl[232] br[232] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_235 
+ bl[233] br[233] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_236 
+ bl[234] br[234] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_237 
+ bl[235] br[235] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_238 
+ bl[236] br[236] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_239 
+ bl[237] br[237] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_240 
+ bl[238] br[238] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_241 
+ bl[239] br[239] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_242 
+ bl[240] br[240] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_243 
+ bl[241] br[241] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_244 
+ bl[242] br[242] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_245 
+ bl[243] br[243] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_246 
+ bl[244] br[244] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_247 
+ bl[245] br[245] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_248 
+ bl[246] br[246] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_249 
+ bl[247] br[247] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_250 
+ bl[248] br[248] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_251 
+ bl[249] br[249] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_252 
+ bl[250] br[250] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_253 
+ bl[251] br[251] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_254 
+ bl[252] br[252] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_255 
+ bl[253] br[253] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_256 
+ bl[254] br[254] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_257 
+ bl[255] br[255] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_258 
+ vdd vdd vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_259 
+ vdd vdd vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_0 
+ vdd vdd vss vdd vpb vnb wl[61] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_63_1 
+ rbl rbr vss vdd vpb vnb wl[61] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_63_2 
+ bl[0] br[0] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_3 
+ bl[1] br[1] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_4 
+ bl[2] br[2] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_5 
+ bl[3] br[3] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_6 
+ bl[4] br[4] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_7 
+ bl[5] br[5] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_8 
+ bl[6] br[6] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_9 
+ bl[7] br[7] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_10 
+ bl[8] br[8] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_11 
+ bl[9] br[9] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_12 
+ bl[10] br[10] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_13 
+ bl[11] br[11] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_14 
+ bl[12] br[12] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_15 
+ bl[13] br[13] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_16 
+ bl[14] br[14] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_17 
+ bl[15] br[15] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_18 
+ bl[16] br[16] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_19 
+ bl[17] br[17] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_20 
+ bl[18] br[18] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_21 
+ bl[19] br[19] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_22 
+ bl[20] br[20] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_23 
+ bl[21] br[21] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_24 
+ bl[22] br[22] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_25 
+ bl[23] br[23] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_26 
+ bl[24] br[24] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_27 
+ bl[25] br[25] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_28 
+ bl[26] br[26] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_29 
+ bl[27] br[27] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_30 
+ bl[28] br[28] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_31 
+ bl[29] br[29] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_32 
+ bl[30] br[30] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_33 
+ bl[31] br[31] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_34 
+ bl[32] br[32] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_35 
+ bl[33] br[33] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_36 
+ bl[34] br[34] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_37 
+ bl[35] br[35] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_38 
+ bl[36] br[36] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_39 
+ bl[37] br[37] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_40 
+ bl[38] br[38] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_41 
+ bl[39] br[39] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_42 
+ bl[40] br[40] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_43 
+ bl[41] br[41] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_44 
+ bl[42] br[42] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_45 
+ bl[43] br[43] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_46 
+ bl[44] br[44] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_47 
+ bl[45] br[45] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_48 
+ bl[46] br[46] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_49 
+ bl[47] br[47] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_50 
+ bl[48] br[48] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_51 
+ bl[49] br[49] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_52 
+ bl[50] br[50] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_53 
+ bl[51] br[51] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_54 
+ bl[52] br[52] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_55 
+ bl[53] br[53] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_56 
+ bl[54] br[54] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_57 
+ bl[55] br[55] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_58 
+ bl[56] br[56] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_59 
+ bl[57] br[57] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_60 
+ bl[58] br[58] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_61 
+ bl[59] br[59] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_62 
+ bl[60] br[60] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_63 
+ bl[61] br[61] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_64 
+ bl[62] br[62] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_65 
+ bl[63] br[63] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_66 
+ bl[64] br[64] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_67 
+ bl[65] br[65] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_68 
+ bl[66] br[66] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_69 
+ bl[67] br[67] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_70 
+ bl[68] br[68] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_71 
+ bl[69] br[69] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_72 
+ bl[70] br[70] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_73 
+ bl[71] br[71] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_74 
+ bl[72] br[72] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_75 
+ bl[73] br[73] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_76 
+ bl[74] br[74] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_77 
+ bl[75] br[75] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_78 
+ bl[76] br[76] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_79 
+ bl[77] br[77] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_80 
+ bl[78] br[78] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_81 
+ bl[79] br[79] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_82 
+ bl[80] br[80] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_83 
+ bl[81] br[81] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_84 
+ bl[82] br[82] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_85 
+ bl[83] br[83] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_86 
+ bl[84] br[84] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_87 
+ bl[85] br[85] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_88 
+ bl[86] br[86] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_89 
+ bl[87] br[87] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_90 
+ bl[88] br[88] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_91 
+ bl[89] br[89] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_92 
+ bl[90] br[90] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_93 
+ bl[91] br[91] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_94 
+ bl[92] br[92] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_95 
+ bl[93] br[93] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_96 
+ bl[94] br[94] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_97 
+ bl[95] br[95] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_98 
+ bl[96] br[96] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_99 
+ bl[97] br[97] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_100 
+ bl[98] br[98] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_101 
+ bl[99] br[99] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_102 
+ bl[100] br[100] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_103 
+ bl[101] br[101] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_104 
+ bl[102] br[102] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_105 
+ bl[103] br[103] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_106 
+ bl[104] br[104] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_107 
+ bl[105] br[105] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_108 
+ bl[106] br[106] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_109 
+ bl[107] br[107] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_110 
+ bl[108] br[108] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_111 
+ bl[109] br[109] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_112 
+ bl[110] br[110] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_113 
+ bl[111] br[111] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_114 
+ bl[112] br[112] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_115 
+ bl[113] br[113] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_116 
+ bl[114] br[114] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_117 
+ bl[115] br[115] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_118 
+ bl[116] br[116] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_119 
+ bl[117] br[117] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_120 
+ bl[118] br[118] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_121 
+ bl[119] br[119] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_122 
+ bl[120] br[120] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_123 
+ bl[121] br[121] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_124 
+ bl[122] br[122] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_125 
+ bl[123] br[123] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_126 
+ bl[124] br[124] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_127 
+ bl[125] br[125] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_128 
+ bl[126] br[126] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_129 
+ bl[127] br[127] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_130 
+ bl[128] br[128] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_131 
+ bl[129] br[129] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_132 
+ bl[130] br[130] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_133 
+ bl[131] br[131] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_134 
+ bl[132] br[132] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_135 
+ bl[133] br[133] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_136 
+ bl[134] br[134] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_137 
+ bl[135] br[135] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_138 
+ bl[136] br[136] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_139 
+ bl[137] br[137] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_140 
+ bl[138] br[138] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_141 
+ bl[139] br[139] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_142 
+ bl[140] br[140] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_143 
+ bl[141] br[141] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_144 
+ bl[142] br[142] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_145 
+ bl[143] br[143] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_146 
+ bl[144] br[144] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_147 
+ bl[145] br[145] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_148 
+ bl[146] br[146] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_149 
+ bl[147] br[147] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_150 
+ bl[148] br[148] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_151 
+ bl[149] br[149] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_152 
+ bl[150] br[150] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_153 
+ bl[151] br[151] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_154 
+ bl[152] br[152] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_155 
+ bl[153] br[153] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_156 
+ bl[154] br[154] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_157 
+ bl[155] br[155] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_158 
+ bl[156] br[156] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_159 
+ bl[157] br[157] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_160 
+ bl[158] br[158] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_161 
+ bl[159] br[159] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_162 
+ bl[160] br[160] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_163 
+ bl[161] br[161] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_164 
+ bl[162] br[162] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_165 
+ bl[163] br[163] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_166 
+ bl[164] br[164] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_167 
+ bl[165] br[165] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_168 
+ bl[166] br[166] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_169 
+ bl[167] br[167] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_170 
+ bl[168] br[168] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_171 
+ bl[169] br[169] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_172 
+ bl[170] br[170] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_173 
+ bl[171] br[171] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_174 
+ bl[172] br[172] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_175 
+ bl[173] br[173] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_176 
+ bl[174] br[174] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_177 
+ bl[175] br[175] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_178 
+ bl[176] br[176] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_179 
+ bl[177] br[177] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_180 
+ bl[178] br[178] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_181 
+ bl[179] br[179] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_182 
+ bl[180] br[180] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_183 
+ bl[181] br[181] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_184 
+ bl[182] br[182] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_185 
+ bl[183] br[183] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_186 
+ bl[184] br[184] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_187 
+ bl[185] br[185] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_188 
+ bl[186] br[186] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_189 
+ bl[187] br[187] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_190 
+ bl[188] br[188] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_191 
+ bl[189] br[189] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_192 
+ bl[190] br[190] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_193 
+ bl[191] br[191] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_194 
+ bl[192] br[192] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_195 
+ bl[193] br[193] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_196 
+ bl[194] br[194] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_197 
+ bl[195] br[195] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_198 
+ bl[196] br[196] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_199 
+ bl[197] br[197] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_200 
+ bl[198] br[198] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_201 
+ bl[199] br[199] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_202 
+ bl[200] br[200] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_203 
+ bl[201] br[201] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_204 
+ bl[202] br[202] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_205 
+ bl[203] br[203] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_206 
+ bl[204] br[204] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_207 
+ bl[205] br[205] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_208 
+ bl[206] br[206] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_209 
+ bl[207] br[207] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_210 
+ bl[208] br[208] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_211 
+ bl[209] br[209] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_212 
+ bl[210] br[210] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_213 
+ bl[211] br[211] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_214 
+ bl[212] br[212] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_215 
+ bl[213] br[213] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_216 
+ bl[214] br[214] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_217 
+ bl[215] br[215] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_218 
+ bl[216] br[216] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_219 
+ bl[217] br[217] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_220 
+ bl[218] br[218] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_221 
+ bl[219] br[219] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_222 
+ bl[220] br[220] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_223 
+ bl[221] br[221] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_224 
+ bl[222] br[222] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_225 
+ bl[223] br[223] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_226 
+ bl[224] br[224] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_227 
+ bl[225] br[225] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_228 
+ bl[226] br[226] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_229 
+ bl[227] br[227] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_230 
+ bl[228] br[228] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_231 
+ bl[229] br[229] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_232 
+ bl[230] br[230] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_233 
+ bl[231] br[231] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_234 
+ bl[232] br[232] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_235 
+ bl[233] br[233] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_236 
+ bl[234] br[234] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_237 
+ bl[235] br[235] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_238 
+ bl[236] br[236] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_239 
+ bl[237] br[237] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_240 
+ bl[238] br[238] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_241 
+ bl[239] br[239] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_242 
+ bl[240] br[240] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_243 
+ bl[241] br[241] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_244 
+ bl[242] br[242] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_245 
+ bl[243] br[243] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_246 
+ bl[244] br[244] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_247 
+ bl[245] br[245] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_248 
+ bl[246] br[246] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_249 
+ bl[247] br[247] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_250 
+ bl[248] br[248] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_251 
+ bl[249] br[249] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_252 
+ bl[250] br[250] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_253 
+ bl[251] br[251] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_254 
+ bl[252] br[252] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_255 
+ bl[253] br[253] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_256 
+ bl[254] br[254] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_257 
+ bl[255] br[255] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_258 
+ vdd vdd vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_259 
+ vdd vdd vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_0 
+ vdd vdd vss vdd vpb vnb wl[62] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_64_1 
+ rbl rbr vss vdd vpb vnb wl[62] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_64_2 
+ bl[0] br[0] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_3 
+ bl[1] br[1] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_4 
+ bl[2] br[2] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_5 
+ bl[3] br[3] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_6 
+ bl[4] br[4] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_7 
+ bl[5] br[5] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_8 
+ bl[6] br[6] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_9 
+ bl[7] br[7] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_10 
+ bl[8] br[8] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_11 
+ bl[9] br[9] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_12 
+ bl[10] br[10] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_13 
+ bl[11] br[11] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_14 
+ bl[12] br[12] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_15 
+ bl[13] br[13] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_16 
+ bl[14] br[14] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_17 
+ bl[15] br[15] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_18 
+ bl[16] br[16] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_19 
+ bl[17] br[17] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_20 
+ bl[18] br[18] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_21 
+ bl[19] br[19] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_22 
+ bl[20] br[20] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_23 
+ bl[21] br[21] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_24 
+ bl[22] br[22] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_25 
+ bl[23] br[23] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_26 
+ bl[24] br[24] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_27 
+ bl[25] br[25] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_28 
+ bl[26] br[26] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_29 
+ bl[27] br[27] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_30 
+ bl[28] br[28] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_31 
+ bl[29] br[29] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_32 
+ bl[30] br[30] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_33 
+ bl[31] br[31] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_34 
+ bl[32] br[32] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_35 
+ bl[33] br[33] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_36 
+ bl[34] br[34] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_37 
+ bl[35] br[35] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_38 
+ bl[36] br[36] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_39 
+ bl[37] br[37] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_40 
+ bl[38] br[38] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_41 
+ bl[39] br[39] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_42 
+ bl[40] br[40] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_43 
+ bl[41] br[41] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_44 
+ bl[42] br[42] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_45 
+ bl[43] br[43] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_46 
+ bl[44] br[44] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_47 
+ bl[45] br[45] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_48 
+ bl[46] br[46] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_49 
+ bl[47] br[47] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_50 
+ bl[48] br[48] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_51 
+ bl[49] br[49] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_52 
+ bl[50] br[50] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_53 
+ bl[51] br[51] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_54 
+ bl[52] br[52] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_55 
+ bl[53] br[53] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_56 
+ bl[54] br[54] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_57 
+ bl[55] br[55] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_58 
+ bl[56] br[56] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_59 
+ bl[57] br[57] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_60 
+ bl[58] br[58] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_61 
+ bl[59] br[59] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_62 
+ bl[60] br[60] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_63 
+ bl[61] br[61] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_64 
+ bl[62] br[62] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_65 
+ bl[63] br[63] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_66 
+ bl[64] br[64] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_67 
+ bl[65] br[65] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_68 
+ bl[66] br[66] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_69 
+ bl[67] br[67] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_70 
+ bl[68] br[68] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_71 
+ bl[69] br[69] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_72 
+ bl[70] br[70] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_73 
+ bl[71] br[71] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_74 
+ bl[72] br[72] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_75 
+ bl[73] br[73] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_76 
+ bl[74] br[74] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_77 
+ bl[75] br[75] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_78 
+ bl[76] br[76] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_79 
+ bl[77] br[77] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_80 
+ bl[78] br[78] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_81 
+ bl[79] br[79] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_82 
+ bl[80] br[80] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_83 
+ bl[81] br[81] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_84 
+ bl[82] br[82] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_85 
+ bl[83] br[83] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_86 
+ bl[84] br[84] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_87 
+ bl[85] br[85] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_88 
+ bl[86] br[86] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_89 
+ bl[87] br[87] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_90 
+ bl[88] br[88] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_91 
+ bl[89] br[89] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_92 
+ bl[90] br[90] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_93 
+ bl[91] br[91] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_94 
+ bl[92] br[92] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_95 
+ bl[93] br[93] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_96 
+ bl[94] br[94] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_97 
+ bl[95] br[95] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_98 
+ bl[96] br[96] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_99 
+ bl[97] br[97] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_100 
+ bl[98] br[98] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_101 
+ bl[99] br[99] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_102 
+ bl[100] br[100] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_103 
+ bl[101] br[101] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_104 
+ bl[102] br[102] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_105 
+ bl[103] br[103] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_106 
+ bl[104] br[104] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_107 
+ bl[105] br[105] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_108 
+ bl[106] br[106] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_109 
+ bl[107] br[107] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_110 
+ bl[108] br[108] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_111 
+ bl[109] br[109] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_112 
+ bl[110] br[110] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_113 
+ bl[111] br[111] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_114 
+ bl[112] br[112] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_115 
+ bl[113] br[113] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_116 
+ bl[114] br[114] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_117 
+ bl[115] br[115] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_118 
+ bl[116] br[116] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_119 
+ bl[117] br[117] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_120 
+ bl[118] br[118] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_121 
+ bl[119] br[119] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_122 
+ bl[120] br[120] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_123 
+ bl[121] br[121] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_124 
+ bl[122] br[122] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_125 
+ bl[123] br[123] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_126 
+ bl[124] br[124] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_127 
+ bl[125] br[125] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_128 
+ bl[126] br[126] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_129 
+ bl[127] br[127] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_130 
+ bl[128] br[128] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_131 
+ bl[129] br[129] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_132 
+ bl[130] br[130] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_133 
+ bl[131] br[131] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_134 
+ bl[132] br[132] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_135 
+ bl[133] br[133] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_136 
+ bl[134] br[134] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_137 
+ bl[135] br[135] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_138 
+ bl[136] br[136] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_139 
+ bl[137] br[137] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_140 
+ bl[138] br[138] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_141 
+ bl[139] br[139] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_142 
+ bl[140] br[140] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_143 
+ bl[141] br[141] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_144 
+ bl[142] br[142] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_145 
+ bl[143] br[143] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_146 
+ bl[144] br[144] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_147 
+ bl[145] br[145] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_148 
+ bl[146] br[146] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_149 
+ bl[147] br[147] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_150 
+ bl[148] br[148] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_151 
+ bl[149] br[149] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_152 
+ bl[150] br[150] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_153 
+ bl[151] br[151] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_154 
+ bl[152] br[152] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_155 
+ bl[153] br[153] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_156 
+ bl[154] br[154] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_157 
+ bl[155] br[155] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_158 
+ bl[156] br[156] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_159 
+ bl[157] br[157] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_160 
+ bl[158] br[158] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_161 
+ bl[159] br[159] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_162 
+ bl[160] br[160] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_163 
+ bl[161] br[161] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_164 
+ bl[162] br[162] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_165 
+ bl[163] br[163] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_166 
+ bl[164] br[164] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_167 
+ bl[165] br[165] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_168 
+ bl[166] br[166] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_169 
+ bl[167] br[167] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_170 
+ bl[168] br[168] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_171 
+ bl[169] br[169] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_172 
+ bl[170] br[170] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_173 
+ bl[171] br[171] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_174 
+ bl[172] br[172] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_175 
+ bl[173] br[173] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_176 
+ bl[174] br[174] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_177 
+ bl[175] br[175] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_178 
+ bl[176] br[176] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_179 
+ bl[177] br[177] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_180 
+ bl[178] br[178] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_181 
+ bl[179] br[179] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_182 
+ bl[180] br[180] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_183 
+ bl[181] br[181] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_184 
+ bl[182] br[182] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_185 
+ bl[183] br[183] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_186 
+ bl[184] br[184] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_187 
+ bl[185] br[185] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_188 
+ bl[186] br[186] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_189 
+ bl[187] br[187] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_190 
+ bl[188] br[188] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_191 
+ bl[189] br[189] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_192 
+ bl[190] br[190] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_193 
+ bl[191] br[191] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_194 
+ bl[192] br[192] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_195 
+ bl[193] br[193] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_196 
+ bl[194] br[194] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_197 
+ bl[195] br[195] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_198 
+ bl[196] br[196] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_199 
+ bl[197] br[197] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_200 
+ bl[198] br[198] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_201 
+ bl[199] br[199] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_202 
+ bl[200] br[200] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_203 
+ bl[201] br[201] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_204 
+ bl[202] br[202] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_205 
+ bl[203] br[203] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_206 
+ bl[204] br[204] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_207 
+ bl[205] br[205] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_208 
+ bl[206] br[206] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_209 
+ bl[207] br[207] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_210 
+ bl[208] br[208] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_211 
+ bl[209] br[209] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_212 
+ bl[210] br[210] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_213 
+ bl[211] br[211] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_214 
+ bl[212] br[212] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_215 
+ bl[213] br[213] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_216 
+ bl[214] br[214] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_217 
+ bl[215] br[215] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_218 
+ bl[216] br[216] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_219 
+ bl[217] br[217] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_220 
+ bl[218] br[218] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_221 
+ bl[219] br[219] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_222 
+ bl[220] br[220] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_223 
+ bl[221] br[221] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_224 
+ bl[222] br[222] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_225 
+ bl[223] br[223] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_226 
+ bl[224] br[224] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_227 
+ bl[225] br[225] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_228 
+ bl[226] br[226] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_229 
+ bl[227] br[227] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_230 
+ bl[228] br[228] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_231 
+ bl[229] br[229] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_232 
+ bl[230] br[230] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_233 
+ bl[231] br[231] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_234 
+ bl[232] br[232] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_235 
+ bl[233] br[233] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_236 
+ bl[234] br[234] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_237 
+ bl[235] br[235] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_238 
+ bl[236] br[236] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_239 
+ bl[237] br[237] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_240 
+ bl[238] br[238] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_241 
+ bl[239] br[239] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_242 
+ bl[240] br[240] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_243 
+ bl[241] br[241] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_244 
+ bl[242] br[242] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_245 
+ bl[243] br[243] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_246 
+ bl[244] br[244] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_247 
+ bl[245] br[245] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_248 
+ bl[246] br[246] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_249 
+ bl[247] br[247] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_250 
+ bl[248] br[248] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_251 
+ bl[249] br[249] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_252 
+ bl[250] br[250] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_253 
+ bl[251] br[251] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_254 
+ bl[252] br[252] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_255 
+ bl[253] br[253] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_256 
+ bl[254] br[254] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_257 
+ bl[255] br[255] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_258 
+ vdd vdd vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_259 
+ vdd vdd vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_0 
+ vdd vdd vss vdd vpb vnb wl[63] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_65_1 
+ rbl rbr vss vdd vpb vnb wl[63] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_65_2 
+ bl[0] br[0] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_3 
+ bl[1] br[1] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_4 
+ bl[2] br[2] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_5 
+ bl[3] br[3] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_6 
+ bl[4] br[4] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_7 
+ bl[5] br[5] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_8 
+ bl[6] br[6] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_9 
+ bl[7] br[7] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_10 
+ bl[8] br[8] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_11 
+ bl[9] br[9] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_12 
+ bl[10] br[10] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_13 
+ bl[11] br[11] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_14 
+ bl[12] br[12] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_15 
+ bl[13] br[13] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_16 
+ bl[14] br[14] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_17 
+ bl[15] br[15] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_18 
+ bl[16] br[16] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_19 
+ bl[17] br[17] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_20 
+ bl[18] br[18] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_21 
+ bl[19] br[19] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_22 
+ bl[20] br[20] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_23 
+ bl[21] br[21] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_24 
+ bl[22] br[22] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_25 
+ bl[23] br[23] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_26 
+ bl[24] br[24] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_27 
+ bl[25] br[25] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_28 
+ bl[26] br[26] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_29 
+ bl[27] br[27] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_30 
+ bl[28] br[28] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_31 
+ bl[29] br[29] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_32 
+ bl[30] br[30] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_33 
+ bl[31] br[31] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_34 
+ bl[32] br[32] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_35 
+ bl[33] br[33] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_36 
+ bl[34] br[34] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_37 
+ bl[35] br[35] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_38 
+ bl[36] br[36] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_39 
+ bl[37] br[37] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_40 
+ bl[38] br[38] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_41 
+ bl[39] br[39] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_42 
+ bl[40] br[40] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_43 
+ bl[41] br[41] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_44 
+ bl[42] br[42] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_45 
+ bl[43] br[43] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_46 
+ bl[44] br[44] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_47 
+ bl[45] br[45] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_48 
+ bl[46] br[46] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_49 
+ bl[47] br[47] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_50 
+ bl[48] br[48] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_51 
+ bl[49] br[49] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_52 
+ bl[50] br[50] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_53 
+ bl[51] br[51] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_54 
+ bl[52] br[52] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_55 
+ bl[53] br[53] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_56 
+ bl[54] br[54] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_57 
+ bl[55] br[55] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_58 
+ bl[56] br[56] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_59 
+ bl[57] br[57] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_60 
+ bl[58] br[58] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_61 
+ bl[59] br[59] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_62 
+ bl[60] br[60] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_63 
+ bl[61] br[61] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_64 
+ bl[62] br[62] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_65 
+ bl[63] br[63] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_66 
+ bl[64] br[64] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_67 
+ bl[65] br[65] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_68 
+ bl[66] br[66] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_69 
+ bl[67] br[67] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_70 
+ bl[68] br[68] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_71 
+ bl[69] br[69] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_72 
+ bl[70] br[70] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_73 
+ bl[71] br[71] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_74 
+ bl[72] br[72] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_75 
+ bl[73] br[73] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_76 
+ bl[74] br[74] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_77 
+ bl[75] br[75] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_78 
+ bl[76] br[76] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_79 
+ bl[77] br[77] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_80 
+ bl[78] br[78] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_81 
+ bl[79] br[79] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_82 
+ bl[80] br[80] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_83 
+ bl[81] br[81] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_84 
+ bl[82] br[82] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_85 
+ bl[83] br[83] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_86 
+ bl[84] br[84] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_87 
+ bl[85] br[85] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_88 
+ bl[86] br[86] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_89 
+ bl[87] br[87] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_90 
+ bl[88] br[88] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_91 
+ bl[89] br[89] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_92 
+ bl[90] br[90] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_93 
+ bl[91] br[91] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_94 
+ bl[92] br[92] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_95 
+ bl[93] br[93] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_96 
+ bl[94] br[94] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_97 
+ bl[95] br[95] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_98 
+ bl[96] br[96] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_99 
+ bl[97] br[97] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_100 
+ bl[98] br[98] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_101 
+ bl[99] br[99] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_102 
+ bl[100] br[100] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_103 
+ bl[101] br[101] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_104 
+ bl[102] br[102] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_105 
+ bl[103] br[103] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_106 
+ bl[104] br[104] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_107 
+ bl[105] br[105] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_108 
+ bl[106] br[106] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_109 
+ bl[107] br[107] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_110 
+ bl[108] br[108] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_111 
+ bl[109] br[109] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_112 
+ bl[110] br[110] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_113 
+ bl[111] br[111] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_114 
+ bl[112] br[112] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_115 
+ bl[113] br[113] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_116 
+ bl[114] br[114] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_117 
+ bl[115] br[115] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_118 
+ bl[116] br[116] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_119 
+ bl[117] br[117] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_120 
+ bl[118] br[118] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_121 
+ bl[119] br[119] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_122 
+ bl[120] br[120] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_123 
+ bl[121] br[121] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_124 
+ bl[122] br[122] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_125 
+ bl[123] br[123] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_126 
+ bl[124] br[124] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_127 
+ bl[125] br[125] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_128 
+ bl[126] br[126] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_129 
+ bl[127] br[127] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_130 
+ bl[128] br[128] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_131 
+ bl[129] br[129] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_132 
+ bl[130] br[130] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_133 
+ bl[131] br[131] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_134 
+ bl[132] br[132] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_135 
+ bl[133] br[133] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_136 
+ bl[134] br[134] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_137 
+ bl[135] br[135] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_138 
+ bl[136] br[136] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_139 
+ bl[137] br[137] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_140 
+ bl[138] br[138] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_141 
+ bl[139] br[139] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_142 
+ bl[140] br[140] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_143 
+ bl[141] br[141] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_144 
+ bl[142] br[142] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_145 
+ bl[143] br[143] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_146 
+ bl[144] br[144] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_147 
+ bl[145] br[145] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_148 
+ bl[146] br[146] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_149 
+ bl[147] br[147] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_150 
+ bl[148] br[148] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_151 
+ bl[149] br[149] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_152 
+ bl[150] br[150] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_153 
+ bl[151] br[151] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_154 
+ bl[152] br[152] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_155 
+ bl[153] br[153] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_156 
+ bl[154] br[154] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_157 
+ bl[155] br[155] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_158 
+ bl[156] br[156] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_159 
+ bl[157] br[157] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_160 
+ bl[158] br[158] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_161 
+ bl[159] br[159] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_162 
+ bl[160] br[160] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_163 
+ bl[161] br[161] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_164 
+ bl[162] br[162] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_165 
+ bl[163] br[163] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_166 
+ bl[164] br[164] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_167 
+ bl[165] br[165] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_168 
+ bl[166] br[166] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_169 
+ bl[167] br[167] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_170 
+ bl[168] br[168] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_171 
+ bl[169] br[169] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_172 
+ bl[170] br[170] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_173 
+ bl[171] br[171] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_174 
+ bl[172] br[172] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_175 
+ bl[173] br[173] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_176 
+ bl[174] br[174] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_177 
+ bl[175] br[175] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_178 
+ bl[176] br[176] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_179 
+ bl[177] br[177] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_180 
+ bl[178] br[178] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_181 
+ bl[179] br[179] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_182 
+ bl[180] br[180] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_183 
+ bl[181] br[181] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_184 
+ bl[182] br[182] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_185 
+ bl[183] br[183] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_186 
+ bl[184] br[184] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_187 
+ bl[185] br[185] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_188 
+ bl[186] br[186] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_189 
+ bl[187] br[187] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_190 
+ bl[188] br[188] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_191 
+ bl[189] br[189] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_192 
+ bl[190] br[190] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_193 
+ bl[191] br[191] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_194 
+ bl[192] br[192] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_195 
+ bl[193] br[193] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_196 
+ bl[194] br[194] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_197 
+ bl[195] br[195] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_198 
+ bl[196] br[196] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_199 
+ bl[197] br[197] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_200 
+ bl[198] br[198] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_201 
+ bl[199] br[199] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_202 
+ bl[200] br[200] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_203 
+ bl[201] br[201] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_204 
+ bl[202] br[202] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_205 
+ bl[203] br[203] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_206 
+ bl[204] br[204] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_207 
+ bl[205] br[205] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_208 
+ bl[206] br[206] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_209 
+ bl[207] br[207] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_210 
+ bl[208] br[208] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_211 
+ bl[209] br[209] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_212 
+ bl[210] br[210] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_213 
+ bl[211] br[211] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_214 
+ bl[212] br[212] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_215 
+ bl[213] br[213] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_216 
+ bl[214] br[214] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_217 
+ bl[215] br[215] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_218 
+ bl[216] br[216] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_219 
+ bl[217] br[217] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_220 
+ bl[218] br[218] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_221 
+ bl[219] br[219] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_222 
+ bl[220] br[220] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_223 
+ bl[221] br[221] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_224 
+ bl[222] br[222] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_225 
+ bl[223] br[223] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_226 
+ bl[224] br[224] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_227 
+ bl[225] br[225] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_228 
+ bl[226] br[226] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_229 
+ bl[227] br[227] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_230 
+ bl[228] br[228] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_231 
+ bl[229] br[229] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_232 
+ bl[230] br[230] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_233 
+ bl[231] br[231] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_234 
+ bl[232] br[232] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_235 
+ bl[233] br[233] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_236 
+ bl[234] br[234] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_237 
+ bl[235] br[235] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_238 
+ bl[236] br[236] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_239 
+ bl[237] br[237] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_240 
+ bl[238] br[238] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_241 
+ bl[239] br[239] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_242 
+ bl[240] br[240] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_243 
+ bl[241] br[241] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_244 
+ bl[242] br[242] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_245 
+ bl[243] br[243] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_246 
+ bl[244] br[244] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_247 
+ bl[245] br[245] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_248 
+ bl[246] br[246] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_249 
+ bl[247] br[247] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_250 
+ bl[248] br[248] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_251 
+ bl[249] br[249] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_252 
+ bl[250] br[250] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_253 
+ bl[251] br[251] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_254 
+ bl[252] br[252] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_255 
+ bl[253] br[253] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_256 
+ bl[254] br[254] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_257 
+ bl[255] br[255] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_258 
+ vdd vdd vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_259 
+ vdd vdd vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_0 
+ vdd vdd vss vdd vpb vnb wl[64] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_66_1 
+ rbl rbr vss vdd vpb vnb wl[64] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_66_2 
+ bl[0] br[0] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_3 
+ bl[1] br[1] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_4 
+ bl[2] br[2] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_5 
+ bl[3] br[3] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_6 
+ bl[4] br[4] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_7 
+ bl[5] br[5] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_8 
+ bl[6] br[6] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_9 
+ bl[7] br[7] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_10 
+ bl[8] br[8] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_11 
+ bl[9] br[9] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_12 
+ bl[10] br[10] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_13 
+ bl[11] br[11] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_14 
+ bl[12] br[12] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_15 
+ bl[13] br[13] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_16 
+ bl[14] br[14] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_17 
+ bl[15] br[15] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_18 
+ bl[16] br[16] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_19 
+ bl[17] br[17] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_20 
+ bl[18] br[18] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_21 
+ bl[19] br[19] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_22 
+ bl[20] br[20] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_23 
+ bl[21] br[21] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_24 
+ bl[22] br[22] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_25 
+ bl[23] br[23] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_26 
+ bl[24] br[24] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_27 
+ bl[25] br[25] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_28 
+ bl[26] br[26] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_29 
+ bl[27] br[27] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_30 
+ bl[28] br[28] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_31 
+ bl[29] br[29] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_32 
+ bl[30] br[30] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_33 
+ bl[31] br[31] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_34 
+ bl[32] br[32] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_35 
+ bl[33] br[33] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_36 
+ bl[34] br[34] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_37 
+ bl[35] br[35] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_38 
+ bl[36] br[36] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_39 
+ bl[37] br[37] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_40 
+ bl[38] br[38] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_41 
+ bl[39] br[39] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_42 
+ bl[40] br[40] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_43 
+ bl[41] br[41] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_44 
+ bl[42] br[42] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_45 
+ bl[43] br[43] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_46 
+ bl[44] br[44] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_47 
+ bl[45] br[45] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_48 
+ bl[46] br[46] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_49 
+ bl[47] br[47] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_50 
+ bl[48] br[48] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_51 
+ bl[49] br[49] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_52 
+ bl[50] br[50] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_53 
+ bl[51] br[51] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_54 
+ bl[52] br[52] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_55 
+ bl[53] br[53] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_56 
+ bl[54] br[54] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_57 
+ bl[55] br[55] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_58 
+ bl[56] br[56] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_59 
+ bl[57] br[57] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_60 
+ bl[58] br[58] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_61 
+ bl[59] br[59] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_62 
+ bl[60] br[60] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_63 
+ bl[61] br[61] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_64 
+ bl[62] br[62] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_65 
+ bl[63] br[63] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_66 
+ bl[64] br[64] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_67 
+ bl[65] br[65] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_68 
+ bl[66] br[66] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_69 
+ bl[67] br[67] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_70 
+ bl[68] br[68] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_71 
+ bl[69] br[69] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_72 
+ bl[70] br[70] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_73 
+ bl[71] br[71] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_74 
+ bl[72] br[72] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_75 
+ bl[73] br[73] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_76 
+ bl[74] br[74] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_77 
+ bl[75] br[75] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_78 
+ bl[76] br[76] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_79 
+ bl[77] br[77] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_80 
+ bl[78] br[78] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_81 
+ bl[79] br[79] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_82 
+ bl[80] br[80] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_83 
+ bl[81] br[81] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_84 
+ bl[82] br[82] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_85 
+ bl[83] br[83] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_86 
+ bl[84] br[84] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_87 
+ bl[85] br[85] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_88 
+ bl[86] br[86] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_89 
+ bl[87] br[87] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_90 
+ bl[88] br[88] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_91 
+ bl[89] br[89] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_92 
+ bl[90] br[90] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_93 
+ bl[91] br[91] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_94 
+ bl[92] br[92] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_95 
+ bl[93] br[93] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_96 
+ bl[94] br[94] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_97 
+ bl[95] br[95] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_98 
+ bl[96] br[96] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_99 
+ bl[97] br[97] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_100 
+ bl[98] br[98] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_101 
+ bl[99] br[99] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_102 
+ bl[100] br[100] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_103 
+ bl[101] br[101] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_104 
+ bl[102] br[102] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_105 
+ bl[103] br[103] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_106 
+ bl[104] br[104] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_107 
+ bl[105] br[105] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_108 
+ bl[106] br[106] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_109 
+ bl[107] br[107] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_110 
+ bl[108] br[108] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_111 
+ bl[109] br[109] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_112 
+ bl[110] br[110] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_113 
+ bl[111] br[111] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_114 
+ bl[112] br[112] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_115 
+ bl[113] br[113] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_116 
+ bl[114] br[114] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_117 
+ bl[115] br[115] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_118 
+ bl[116] br[116] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_119 
+ bl[117] br[117] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_120 
+ bl[118] br[118] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_121 
+ bl[119] br[119] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_122 
+ bl[120] br[120] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_123 
+ bl[121] br[121] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_124 
+ bl[122] br[122] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_125 
+ bl[123] br[123] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_126 
+ bl[124] br[124] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_127 
+ bl[125] br[125] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_128 
+ bl[126] br[126] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_129 
+ bl[127] br[127] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_130 
+ bl[128] br[128] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_131 
+ bl[129] br[129] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_132 
+ bl[130] br[130] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_133 
+ bl[131] br[131] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_134 
+ bl[132] br[132] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_135 
+ bl[133] br[133] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_136 
+ bl[134] br[134] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_137 
+ bl[135] br[135] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_138 
+ bl[136] br[136] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_139 
+ bl[137] br[137] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_140 
+ bl[138] br[138] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_141 
+ bl[139] br[139] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_142 
+ bl[140] br[140] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_143 
+ bl[141] br[141] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_144 
+ bl[142] br[142] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_145 
+ bl[143] br[143] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_146 
+ bl[144] br[144] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_147 
+ bl[145] br[145] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_148 
+ bl[146] br[146] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_149 
+ bl[147] br[147] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_150 
+ bl[148] br[148] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_151 
+ bl[149] br[149] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_152 
+ bl[150] br[150] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_153 
+ bl[151] br[151] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_154 
+ bl[152] br[152] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_155 
+ bl[153] br[153] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_156 
+ bl[154] br[154] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_157 
+ bl[155] br[155] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_158 
+ bl[156] br[156] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_159 
+ bl[157] br[157] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_160 
+ bl[158] br[158] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_161 
+ bl[159] br[159] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_162 
+ bl[160] br[160] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_163 
+ bl[161] br[161] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_164 
+ bl[162] br[162] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_165 
+ bl[163] br[163] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_166 
+ bl[164] br[164] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_167 
+ bl[165] br[165] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_168 
+ bl[166] br[166] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_169 
+ bl[167] br[167] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_170 
+ bl[168] br[168] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_171 
+ bl[169] br[169] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_172 
+ bl[170] br[170] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_173 
+ bl[171] br[171] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_174 
+ bl[172] br[172] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_175 
+ bl[173] br[173] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_176 
+ bl[174] br[174] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_177 
+ bl[175] br[175] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_178 
+ bl[176] br[176] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_179 
+ bl[177] br[177] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_180 
+ bl[178] br[178] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_181 
+ bl[179] br[179] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_182 
+ bl[180] br[180] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_183 
+ bl[181] br[181] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_184 
+ bl[182] br[182] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_185 
+ bl[183] br[183] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_186 
+ bl[184] br[184] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_187 
+ bl[185] br[185] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_188 
+ bl[186] br[186] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_189 
+ bl[187] br[187] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_190 
+ bl[188] br[188] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_191 
+ bl[189] br[189] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_192 
+ bl[190] br[190] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_193 
+ bl[191] br[191] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_194 
+ bl[192] br[192] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_195 
+ bl[193] br[193] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_196 
+ bl[194] br[194] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_197 
+ bl[195] br[195] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_198 
+ bl[196] br[196] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_199 
+ bl[197] br[197] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_200 
+ bl[198] br[198] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_201 
+ bl[199] br[199] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_202 
+ bl[200] br[200] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_203 
+ bl[201] br[201] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_204 
+ bl[202] br[202] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_205 
+ bl[203] br[203] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_206 
+ bl[204] br[204] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_207 
+ bl[205] br[205] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_208 
+ bl[206] br[206] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_209 
+ bl[207] br[207] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_210 
+ bl[208] br[208] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_211 
+ bl[209] br[209] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_212 
+ bl[210] br[210] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_213 
+ bl[211] br[211] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_214 
+ bl[212] br[212] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_215 
+ bl[213] br[213] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_216 
+ bl[214] br[214] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_217 
+ bl[215] br[215] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_218 
+ bl[216] br[216] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_219 
+ bl[217] br[217] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_220 
+ bl[218] br[218] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_221 
+ bl[219] br[219] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_222 
+ bl[220] br[220] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_223 
+ bl[221] br[221] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_224 
+ bl[222] br[222] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_225 
+ bl[223] br[223] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_226 
+ bl[224] br[224] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_227 
+ bl[225] br[225] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_228 
+ bl[226] br[226] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_229 
+ bl[227] br[227] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_230 
+ bl[228] br[228] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_231 
+ bl[229] br[229] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_232 
+ bl[230] br[230] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_233 
+ bl[231] br[231] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_234 
+ bl[232] br[232] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_235 
+ bl[233] br[233] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_236 
+ bl[234] br[234] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_237 
+ bl[235] br[235] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_238 
+ bl[236] br[236] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_239 
+ bl[237] br[237] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_240 
+ bl[238] br[238] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_241 
+ bl[239] br[239] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_242 
+ bl[240] br[240] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_243 
+ bl[241] br[241] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_244 
+ bl[242] br[242] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_245 
+ bl[243] br[243] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_246 
+ bl[244] br[244] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_247 
+ bl[245] br[245] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_248 
+ bl[246] br[246] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_249 
+ bl[247] br[247] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_250 
+ bl[248] br[248] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_251 
+ bl[249] br[249] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_252 
+ bl[250] br[250] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_253 
+ bl[251] br[251] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_254 
+ bl[252] br[252] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_255 
+ bl[253] br[253] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_256 
+ bl[254] br[254] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_257 
+ bl[255] br[255] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_258 
+ vdd vdd vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_259 
+ vdd vdd vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_0 
+ vdd vdd vss vdd vpb vnb wl[65] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_67_1 
+ rbl rbr vss vdd vpb vnb wl[65] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_67_2 
+ bl[0] br[0] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_3 
+ bl[1] br[1] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_4 
+ bl[2] br[2] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_5 
+ bl[3] br[3] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_6 
+ bl[4] br[4] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_7 
+ bl[5] br[5] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_8 
+ bl[6] br[6] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_9 
+ bl[7] br[7] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_10 
+ bl[8] br[8] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_11 
+ bl[9] br[9] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_12 
+ bl[10] br[10] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_13 
+ bl[11] br[11] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_14 
+ bl[12] br[12] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_15 
+ bl[13] br[13] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_16 
+ bl[14] br[14] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_17 
+ bl[15] br[15] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_18 
+ bl[16] br[16] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_19 
+ bl[17] br[17] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_20 
+ bl[18] br[18] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_21 
+ bl[19] br[19] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_22 
+ bl[20] br[20] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_23 
+ bl[21] br[21] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_24 
+ bl[22] br[22] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_25 
+ bl[23] br[23] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_26 
+ bl[24] br[24] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_27 
+ bl[25] br[25] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_28 
+ bl[26] br[26] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_29 
+ bl[27] br[27] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_30 
+ bl[28] br[28] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_31 
+ bl[29] br[29] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_32 
+ bl[30] br[30] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_33 
+ bl[31] br[31] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_34 
+ bl[32] br[32] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_35 
+ bl[33] br[33] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_36 
+ bl[34] br[34] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_37 
+ bl[35] br[35] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_38 
+ bl[36] br[36] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_39 
+ bl[37] br[37] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_40 
+ bl[38] br[38] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_41 
+ bl[39] br[39] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_42 
+ bl[40] br[40] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_43 
+ bl[41] br[41] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_44 
+ bl[42] br[42] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_45 
+ bl[43] br[43] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_46 
+ bl[44] br[44] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_47 
+ bl[45] br[45] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_48 
+ bl[46] br[46] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_49 
+ bl[47] br[47] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_50 
+ bl[48] br[48] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_51 
+ bl[49] br[49] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_52 
+ bl[50] br[50] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_53 
+ bl[51] br[51] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_54 
+ bl[52] br[52] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_55 
+ bl[53] br[53] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_56 
+ bl[54] br[54] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_57 
+ bl[55] br[55] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_58 
+ bl[56] br[56] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_59 
+ bl[57] br[57] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_60 
+ bl[58] br[58] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_61 
+ bl[59] br[59] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_62 
+ bl[60] br[60] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_63 
+ bl[61] br[61] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_64 
+ bl[62] br[62] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_65 
+ bl[63] br[63] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_66 
+ bl[64] br[64] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_67 
+ bl[65] br[65] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_68 
+ bl[66] br[66] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_69 
+ bl[67] br[67] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_70 
+ bl[68] br[68] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_71 
+ bl[69] br[69] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_72 
+ bl[70] br[70] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_73 
+ bl[71] br[71] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_74 
+ bl[72] br[72] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_75 
+ bl[73] br[73] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_76 
+ bl[74] br[74] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_77 
+ bl[75] br[75] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_78 
+ bl[76] br[76] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_79 
+ bl[77] br[77] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_80 
+ bl[78] br[78] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_81 
+ bl[79] br[79] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_82 
+ bl[80] br[80] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_83 
+ bl[81] br[81] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_84 
+ bl[82] br[82] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_85 
+ bl[83] br[83] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_86 
+ bl[84] br[84] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_87 
+ bl[85] br[85] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_88 
+ bl[86] br[86] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_89 
+ bl[87] br[87] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_90 
+ bl[88] br[88] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_91 
+ bl[89] br[89] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_92 
+ bl[90] br[90] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_93 
+ bl[91] br[91] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_94 
+ bl[92] br[92] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_95 
+ bl[93] br[93] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_96 
+ bl[94] br[94] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_97 
+ bl[95] br[95] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_98 
+ bl[96] br[96] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_99 
+ bl[97] br[97] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_100 
+ bl[98] br[98] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_101 
+ bl[99] br[99] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_102 
+ bl[100] br[100] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_103 
+ bl[101] br[101] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_104 
+ bl[102] br[102] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_105 
+ bl[103] br[103] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_106 
+ bl[104] br[104] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_107 
+ bl[105] br[105] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_108 
+ bl[106] br[106] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_109 
+ bl[107] br[107] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_110 
+ bl[108] br[108] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_111 
+ bl[109] br[109] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_112 
+ bl[110] br[110] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_113 
+ bl[111] br[111] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_114 
+ bl[112] br[112] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_115 
+ bl[113] br[113] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_116 
+ bl[114] br[114] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_117 
+ bl[115] br[115] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_118 
+ bl[116] br[116] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_119 
+ bl[117] br[117] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_120 
+ bl[118] br[118] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_121 
+ bl[119] br[119] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_122 
+ bl[120] br[120] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_123 
+ bl[121] br[121] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_124 
+ bl[122] br[122] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_125 
+ bl[123] br[123] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_126 
+ bl[124] br[124] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_127 
+ bl[125] br[125] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_128 
+ bl[126] br[126] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_129 
+ bl[127] br[127] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_130 
+ bl[128] br[128] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_131 
+ bl[129] br[129] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_132 
+ bl[130] br[130] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_133 
+ bl[131] br[131] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_134 
+ bl[132] br[132] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_135 
+ bl[133] br[133] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_136 
+ bl[134] br[134] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_137 
+ bl[135] br[135] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_138 
+ bl[136] br[136] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_139 
+ bl[137] br[137] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_140 
+ bl[138] br[138] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_141 
+ bl[139] br[139] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_142 
+ bl[140] br[140] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_143 
+ bl[141] br[141] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_144 
+ bl[142] br[142] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_145 
+ bl[143] br[143] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_146 
+ bl[144] br[144] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_147 
+ bl[145] br[145] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_148 
+ bl[146] br[146] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_149 
+ bl[147] br[147] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_150 
+ bl[148] br[148] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_151 
+ bl[149] br[149] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_152 
+ bl[150] br[150] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_153 
+ bl[151] br[151] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_154 
+ bl[152] br[152] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_155 
+ bl[153] br[153] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_156 
+ bl[154] br[154] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_157 
+ bl[155] br[155] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_158 
+ bl[156] br[156] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_159 
+ bl[157] br[157] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_160 
+ bl[158] br[158] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_161 
+ bl[159] br[159] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_162 
+ bl[160] br[160] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_163 
+ bl[161] br[161] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_164 
+ bl[162] br[162] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_165 
+ bl[163] br[163] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_166 
+ bl[164] br[164] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_167 
+ bl[165] br[165] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_168 
+ bl[166] br[166] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_169 
+ bl[167] br[167] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_170 
+ bl[168] br[168] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_171 
+ bl[169] br[169] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_172 
+ bl[170] br[170] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_173 
+ bl[171] br[171] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_174 
+ bl[172] br[172] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_175 
+ bl[173] br[173] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_176 
+ bl[174] br[174] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_177 
+ bl[175] br[175] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_178 
+ bl[176] br[176] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_179 
+ bl[177] br[177] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_180 
+ bl[178] br[178] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_181 
+ bl[179] br[179] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_182 
+ bl[180] br[180] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_183 
+ bl[181] br[181] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_184 
+ bl[182] br[182] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_185 
+ bl[183] br[183] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_186 
+ bl[184] br[184] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_187 
+ bl[185] br[185] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_188 
+ bl[186] br[186] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_189 
+ bl[187] br[187] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_190 
+ bl[188] br[188] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_191 
+ bl[189] br[189] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_192 
+ bl[190] br[190] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_193 
+ bl[191] br[191] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_194 
+ bl[192] br[192] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_195 
+ bl[193] br[193] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_196 
+ bl[194] br[194] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_197 
+ bl[195] br[195] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_198 
+ bl[196] br[196] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_199 
+ bl[197] br[197] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_200 
+ bl[198] br[198] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_201 
+ bl[199] br[199] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_202 
+ bl[200] br[200] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_203 
+ bl[201] br[201] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_204 
+ bl[202] br[202] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_205 
+ bl[203] br[203] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_206 
+ bl[204] br[204] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_207 
+ bl[205] br[205] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_208 
+ bl[206] br[206] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_209 
+ bl[207] br[207] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_210 
+ bl[208] br[208] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_211 
+ bl[209] br[209] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_212 
+ bl[210] br[210] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_213 
+ bl[211] br[211] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_214 
+ bl[212] br[212] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_215 
+ bl[213] br[213] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_216 
+ bl[214] br[214] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_217 
+ bl[215] br[215] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_218 
+ bl[216] br[216] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_219 
+ bl[217] br[217] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_220 
+ bl[218] br[218] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_221 
+ bl[219] br[219] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_222 
+ bl[220] br[220] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_223 
+ bl[221] br[221] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_224 
+ bl[222] br[222] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_225 
+ bl[223] br[223] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_226 
+ bl[224] br[224] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_227 
+ bl[225] br[225] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_228 
+ bl[226] br[226] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_229 
+ bl[227] br[227] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_230 
+ bl[228] br[228] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_231 
+ bl[229] br[229] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_232 
+ bl[230] br[230] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_233 
+ bl[231] br[231] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_234 
+ bl[232] br[232] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_235 
+ bl[233] br[233] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_236 
+ bl[234] br[234] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_237 
+ bl[235] br[235] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_238 
+ bl[236] br[236] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_239 
+ bl[237] br[237] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_240 
+ bl[238] br[238] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_241 
+ bl[239] br[239] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_242 
+ bl[240] br[240] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_243 
+ bl[241] br[241] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_244 
+ bl[242] br[242] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_245 
+ bl[243] br[243] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_246 
+ bl[244] br[244] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_247 
+ bl[245] br[245] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_248 
+ bl[246] br[246] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_249 
+ bl[247] br[247] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_250 
+ bl[248] br[248] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_251 
+ bl[249] br[249] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_252 
+ bl[250] br[250] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_253 
+ bl[251] br[251] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_254 
+ bl[252] br[252] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_255 
+ bl[253] br[253] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_256 
+ bl[254] br[254] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_257 
+ bl[255] br[255] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_258 
+ vdd vdd vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_259 
+ vdd vdd vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_0 
+ vdd vdd vss vdd vpb vnb wl[66] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_68_1 
+ rbl rbr vss vdd vpb vnb wl[66] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_68_2 
+ bl[0] br[0] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_3 
+ bl[1] br[1] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_4 
+ bl[2] br[2] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_5 
+ bl[3] br[3] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_6 
+ bl[4] br[4] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_7 
+ bl[5] br[5] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_8 
+ bl[6] br[6] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_9 
+ bl[7] br[7] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_10 
+ bl[8] br[8] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_11 
+ bl[9] br[9] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_12 
+ bl[10] br[10] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_13 
+ bl[11] br[11] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_14 
+ bl[12] br[12] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_15 
+ bl[13] br[13] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_16 
+ bl[14] br[14] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_17 
+ bl[15] br[15] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_18 
+ bl[16] br[16] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_19 
+ bl[17] br[17] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_20 
+ bl[18] br[18] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_21 
+ bl[19] br[19] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_22 
+ bl[20] br[20] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_23 
+ bl[21] br[21] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_24 
+ bl[22] br[22] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_25 
+ bl[23] br[23] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_26 
+ bl[24] br[24] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_27 
+ bl[25] br[25] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_28 
+ bl[26] br[26] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_29 
+ bl[27] br[27] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_30 
+ bl[28] br[28] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_31 
+ bl[29] br[29] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_32 
+ bl[30] br[30] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_33 
+ bl[31] br[31] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_34 
+ bl[32] br[32] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_35 
+ bl[33] br[33] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_36 
+ bl[34] br[34] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_37 
+ bl[35] br[35] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_38 
+ bl[36] br[36] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_39 
+ bl[37] br[37] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_40 
+ bl[38] br[38] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_41 
+ bl[39] br[39] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_42 
+ bl[40] br[40] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_43 
+ bl[41] br[41] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_44 
+ bl[42] br[42] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_45 
+ bl[43] br[43] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_46 
+ bl[44] br[44] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_47 
+ bl[45] br[45] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_48 
+ bl[46] br[46] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_49 
+ bl[47] br[47] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_50 
+ bl[48] br[48] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_51 
+ bl[49] br[49] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_52 
+ bl[50] br[50] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_53 
+ bl[51] br[51] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_54 
+ bl[52] br[52] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_55 
+ bl[53] br[53] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_56 
+ bl[54] br[54] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_57 
+ bl[55] br[55] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_58 
+ bl[56] br[56] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_59 
+ bl[57] br[57] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_60 
+ bl[58] br[58] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_61 
+ bl[59] br[59] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_62 
+ bl[60] br[60] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_63 
+ bl[61] br[61] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_64 
+ bl[62] br[62] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_65 
+ bl[63] br[63] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_66 
+ bl[64] br[64] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_67 
+ bl[65] br[65] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_68 
+ bl[66] br[66] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_69 
+ bl[67] br[67] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_70 
+ bl[68] br[68] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_71 
+ bl[69] br[69] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_72 
+ bl[70] br[70] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_73 
+ bl[71] br[71] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_74 
+ bl[72] br[72] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_75 
+ bl[73] br[73] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_76 
+ bl[74] br[74] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_77 
+ bl[75] br[75] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_78 
+ bl[76] br[76] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_79 
+ bl[77] br[77] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_80 
+ bl[78] br[78] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_81 
+ bl[79] br[79] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_82 
+ bl[80] br[80] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_83 
+ bl[81] br[81] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_84 
+ bl[82] br[82] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_85 
+ bl[83] br[83] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_86 
+ bl[84] br[84] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_87 
+ bl[85] br[85] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_88 
+ bl[86] br[86] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_89 
+ bl[87] br[87] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_90 
+ bl[88] br[88] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_91 
+ bl[89] br[89] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_92 
+ bl[90] br[90] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_93 
+ bl[91] br[91] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_94 
+ bl[92] br[92] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_95 
+ bl[93] br[93] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_96 
+ bl[94] br[94] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_97 
+ bl[95] br[95] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_98 
+ bl[96] br[96] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_99 
+ bl[97] br[97] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_100 
+ bl[98] br[98] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_101 
+ bl[99] br[99] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_102 
+ bl[100] br[100] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_103 
+ bl[101] br[101] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_104 
+ bl[102] br[102] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_105 
+ bl[103] br[103] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_106 
+ bl[104] br[104] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_107 
+ bl[105] br[105] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_108 
+ bl[106] br[106] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_109 
+ bl[107] br[107] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_110 
+ bl[108] br[108] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_111 
+ bl[109] br[109] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_112 
+ bl[110] br[110] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_113 
+ bl[111] br[111] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_114 
+ bl[112] br[112] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_115 
+ bl[113] br[113] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_116 
+ bl[114] br[114] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_117 
+ bl[115] br[115] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_118 
+ bl[116] br[116] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_119 
+ bl[117] br[117] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_120 
+ bl[118] br[118] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_121 
+ bl[119] br[119] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_122 
+ bl[120] br[120] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_123 
+ bl[121] br[121] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_124 
+ bl[122] br[122] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_125 
+ bl[123] br[123] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_126 
+ bl[124] br[124] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_127 
+ bl[125] br[125] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_128 
+ bl[126] br[126] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_129 
+ bl[127] br[127] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_130 
+ bl[128] br[128] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_131 
+ bl[129] br[129] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_132 
+ bl[130] br[130] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_133 
+ bl[131] br[131] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_134 
+ bl[132] br[132] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_135 
+ bl[133] br[133] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_136 
+ bl[134] br[134] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_137 
+ bl[135] br[135] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_138 
+ bl[136] br[136] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_139 
+ bl[137] br[137] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_140 
+ bl[138] br[138] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_141 
+ bl[139] br[139] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_142 
+ bl[140] br[140] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_143 
+ bl[141] br[141] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_144 
+ bl[142] br[142] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_145 
+ bl[143] br[143] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_146 
+ bl[144] br[144] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_147 
+ bl[145] br[145] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_148 
+ bl[146] br[146] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_149 
+ bl[147] br[147] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_150 
+ bl[148] br[148] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_151 
+ bl[149] br[149] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_152 
+ bl[150] br[150] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_153 
+ bl[151] br[151] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_154 
+ bl[152] br[152] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_155 
+ bl[153] br[153] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_156 
+ bl[154] br[154] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_157 
+ bl[155] br[155] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_158 
+ bl[156] br[156] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_159 
+ bl[157] br[157] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_160 
+ bl[158] br[158] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_161 
+ bl[159] br[159] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_162 
+ bl[160] br[160] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_163 
+ bl[161] br[161] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_164 
+ bl[162] br[162] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_165 
+ bl[163] br[163] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_166 
+ bl[164] br[164] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_167 
+ bl[165] br[165] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_168 
+ bl[166] br[166] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_169 
+ bl[167] br[167] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_170 
+ bl[168] br[168] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_171 
+ bl[169] br[169] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_172 
+ bl[170] br[170] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_173 
+ bl[171] br[171] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_174 
+ bl[172] br[172] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_175 
+ bl[173] br[173] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_176 
+ bl[174] br[174] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_177 
+ bl[175] br[175] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_178 
+ bl[176] br[176] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_179 
+ bl[177] br[177] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_180 
+ bl[178] br[178] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_181 
+ bl[179] br[179] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_182 
+ bl[180] br[180] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_183 
+ bl[181] br[181] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_184 
+ bl[182] br[182] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_185 
+ bl[183] br[183] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_186 
+ bl[184] br[184] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_187 
+ bl[185] br[185] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_188 
+ bl[186] br[186] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_189 
+ bl[187] br[187] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_190 
+ bl[188] br[188] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_191 
+ bl[189] br[189] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_192 
+ bl[190] br[190] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_193 
+ bl[191] br[191] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_194 
+ bl[192] br[192] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_195 
+ bl[193] br[193] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_196 
+ bl[194] br[194] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_197 
+ bl[195] br[195] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_198 
+ bl[196] br[196] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_199 
+ bl[197] br[197] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_200 
+ bl[198] br[198] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_201 
+ bl[199] br[199] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_202 
+ bl[200] br[200] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_203 
+ bl[201] br[201] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_204 
+ bl[202] br[202] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_205 
+ bl[203] br[203] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_206 
+ bl[204] br[204] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_207 
+ bl[205] br[205] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_208 
+ bl[206] br[206] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_209 
+ bl[207] br[207] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_210 
+ bl[208] br[208] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_211 
+ bl[209] br[209] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_212 
+ bl[210] br[210] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_213 
+ bl[211] br[211] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_214 
+ bl[212] br[212] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_215 
+ bl[213] br[213] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_216 
+ bl[214] br[214] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_217 
+ bl[215] br[215] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_218 
+ bl[216] br[216] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_219 
+ bl[217] br[217] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_220 
+ bl[218] br[218] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_221 
+ bl[219] br[219] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_222 
+ bl[220] br[220] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_223 
+ bl[221] br[221] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_224 
+ bl[222] br[222] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_225 
+ bl[223] br[223] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_226 
+ bl[224] br[224] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_227 
+ bl[225] br[225] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_228 
+ bl[226] br[226] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_229 
+ bl[227] br[227] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_230 
+ bl[228] br[228] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_231 
+ bl[229] br[229] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_232 
+ bl[230] br[230] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_233 
+ bl[231] br[231] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_234 
+ bl[232] br[232] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_235 
+ bl[233] br[233] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_236 
+ bl[234] br[234] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_237 
+ bl[235] br[235] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_238 
+ bl[236] br[236] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_239 
+ bl[237] br[237] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_240 
+ bl[238] br[238] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_241 
+ bl[239] br[239] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_242 
+ bl[240] br[240] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_243 
+ bl[241] br[241] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_244 
+ bl[242] br[242] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_245 
+ bl[243] br[243] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_246 
+ bl[244] br[244] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_247 
+ bl[245] br[245] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_248 
+ bl[246] br[246] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_249 
+ bl[247] br[247] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_250 
+ bl[248] br[248] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_251 
+ bl[249] br[249] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_252 
+ bl[250] br[250] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_253 
+ bl[251] br[251] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_254 
+ bl[252] br[252] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_255 
+ bl[253] br[253] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_256 
+ bl[254] br[254] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_257 
+ bl[255] br[255] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_258 
+ vdd vdd vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_259 
+ vdd vdd vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_0 
+ vdd vdd vss vdd vpb vnb wl[67] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_69_1 
+ rbl rbr vss vdd vpb vnb wl[67] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_69_2 
+ bl[0] br[0] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_3 
+ bl[1] br[1] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_4 
+ bl[2] br[2] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_5 
+ bl[3] br[3] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_6 
+ bl[4] br[4] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_7 
+ bl[5] br[5] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_8 
+ bl[6] br[6] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_9 
+ bl[7] br[7] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_10 
+ bl[8] br[8] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_11 
+ bl[9] br[9] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_12 
+ bl[10] br[10] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_13 
+ bl[11] br[11] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_14 
+ bl[12] br[12] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_15 
+ bl[13] br[13] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_16 
+ bl[14] br[14] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_17 
+ bl[15] br[15] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_18 
+ bl[16] br[16] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_19 
+ bl[17] br[17] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_20 
+ bl[18] br[18] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_21 
+ bl[19] br[19] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_22 
+ bl[20] br[20] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_23 
+ bl[21] br[21] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_24 
+ bl[22] br[22] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_25 
+ bl[23] br[23] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_26 
+ bl[24] br[24] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_27 
+ bl[25] br[25] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_28 
+ bl[26] br[26] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_29 
+ bl[27] br[27] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_30 
+ bl[28] br[28] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_31 
+ bl[29] br[29] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_32 
+ bl[30] br[30] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_33 
+ bl[31] br[31] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_34 
+ bl[32] br[32] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_35 
+ bl[33] br[33] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_36 
+ bl[34] br[34] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_37 
+ bl[35] br[35] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_38 
+ bl[36] br[36] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_39 
+ bl[37] br[37] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_40 
+ bl[38] br[38] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_41 
+ bl[39] br[39] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_42 
+ bl[40] br[40] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_43 
+ bl[41] br[41] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_44 
+ bl[42] br[42] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_45 
+ bl[43] br[43] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_46 
+ bl[44] br[44] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_47 
+ bl[45] br[45] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_48 
+ bl[46] br[46] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_49 
+ bl[47] br[47] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_50 
+ bl[48] br[48] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_51 
+ bl[49] br[49] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_52 
+ bl[50] br[50] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_53 
+ bl[51] br[51] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_54 
+ bl[52] br[52] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_55 
+ bl[53] br[53] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_56 
+ bl[54] br[54] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_57 
+ bl[55] br[55] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_58 
+ bl[56] br[56] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_59 
+ bl[57] br[57] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_60 
+ bl[58] br[58] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_61 
+ bl[59] br[59] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_62 
+ bl[60] br[60] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_63 
+ bl[61] br[61] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_64 
+ bl[62] br[62] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_65 
+ bl[63] br[63] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_66 
+ bl[64] br[64] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_67 
+ bl[65] br[65] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_68 
+ bl[66] br[66] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_69 
+ bl[67] br[67] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_70 
+ bl[68] br[68] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_71 
+ bl[69] br[69] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_72 
+ bl[70] br[70] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_73 
+ bl[71] br[71] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_74 
+ bl[72] br[72] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_75 
+ bl[73] br[73] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_76 
+ bl[74] br[74] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_77 
+ bl[75] br[75] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_78 
+ bl[76] br[76] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_79 
+ bl[77] br[77] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_80 
+ bl[78] br[78] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_81 
+ bl[79] br[79] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_82 
+ bl[80] br[80] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_83 
+ bl[81] br[81] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_84 
+ bl[82] br[82] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_85 
+ bl[83] br[83] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_86 
+ bl[84] br[84] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_87 
+ bl[85] br[85] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_88 
+ bl[86] br[86] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_89 
+ bl[87] br[87] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_90 
+ bl[88] br[88] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_91 
+ bl[89] br[89] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_92 
+ bl[90] br[90] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_93 
+ bl[91] br[91] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_94 
+ bl[92] br[92] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_95 
+ bl[93] br[93] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_96 
+ bl[94] br[94] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_97 
+ bl[95] br[95] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_98 
+ bl[96] br[96] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_99 
+ bl[97] br[97] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_100 
+ bl[98] br[98] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_101 
+ bl[99] br[99] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_102 
+ bl[100] br[100] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_103 
+ bl[101] br[101] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_104 
+ bl[102] br[102] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_105 
+ bl[103] br[103] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_106 
+ bl[104] br[104] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_107 
+ bl[105] br[105] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_108 
+ bl[106] br[106] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_109 
+ bl[107] br[107] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_110 
+ bl[108] br[108] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_111 
+ bl[109] br[109] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_112 
+ bl[110] br[110] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_113 
+ bl[111] br[111] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_114 
+ bl[112] br[112] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_115 
+ bl[113] br[113] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_116 
+ bl[114] br[114] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_117 
+ bl[115] br[115] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_118 
+ bl[116] br[116] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_119 
+ bl[117] br[117] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_120 
+ bl[118] br[118] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_121 
+ bl[119] br[119] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_122 
+ bl[120] br[120] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_123 
+ bl[121] br[121] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_124 
+ bl[122] br[122] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_125 
+ bl[123] br[123] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_126 
+ bl[124] br[124] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_127 
+ bl[125] br[125] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_128 
+ bl[126] br[126] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_129 
+ bl[127] br[127] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_130 
+ bl[128] br[128] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_131 
+ bl[129] br[129] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_132 
+ bl[130] br[130] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_133 
+ bl[131] br[131] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_134 
+ bl[132] br[132] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_135 
+ bl[133] br[133] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_136 
+ bl[134] br[134] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_137 
+ bl[135] br[135] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_138 
+ bl[136] br[136] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_139 
+ bl[137] br[137] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_140 
+ bl[138] br[138] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_141 
+ bl[139] br[139] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_142 
+ bl[140] br[140] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_143 
+ bl[141] br[141] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_144 
+ bl[142] br[142] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_145 
+ bl[143] br[143] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_146 
+ bl[144] br[144] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_147 
+ bl[145] br[145] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_148 
+ bl[146] br[146] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_149 
+ bl[147] br[147] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_150 
+ bl[148] br[148] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_151 
+ bl[149] br[149] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_152 
+ bl[150] br[150] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_153 
+ bl[151] br[151] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_154 
+ bl[152] br[152] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_155 
+ bl[153] br[153] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_156 
+ bl[154] br[154] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_157 
+ bl[155] br[155] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_158 
+ bl[156] br[156] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_159 
+ bl[157] br[157] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_160 
+ bl[158] br[158] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_161 
+ bl[159] br[159] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_162 
+ bl[160] br[160] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_163 
+ bl[161] br[161] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_164 
+ bl[162] br[162] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_165 
+ bl[163] br[163] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_166 
+ bl[164] br[164] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_167 
+ bl[165] br[165] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_168 
+ bl[166] br[166] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_169 
+ bl[167] br[167] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_170 
+ bl[168] br[168] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_171 
+ bl[169] br[169] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_172 
+ bl[170] br[170] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_173 
+ bl[171] br[171] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_174 
+ bl[172] br[172] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_175 
+ bl[173] br[173] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_176 
+ bl[174] br[174] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_177 
+ bl[175] br[175] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_178 
+ bl[176] br[176] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_179 
+ bl[177] br[177] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_180 
+ bl[178] br[178] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_181 
+ bl[179] br[179] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_182 
+ bl[180] br[180] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_183 
+ bl[181] br[181] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_184 
+ bl[182] br[182] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_185 
+ bl[183] br[183] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_186 
+ bl[184] br[184] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_187 
+ bl[185] br[185] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_188 
+ bl[186] br[186] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_189 
+ bl[187] br[187] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_190 
+ bl[188] br[188] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_191 
+ bl[189] br[189] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_192 
+ bl[190] br[190] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_193 
+ bl[191] br[191] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_194 
+ bl[192] br[192] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_195 
+ bl[193] br[193] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_196 
+ bl[194] br[194] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_197 
+ bl[195] br[195] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_198 
+ bl[196] br[196] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_199 
+ bl[197] br[197] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_200 
+ bl[198] br[198] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_201 
+ bl[199] br[199] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_202 
+ bl[200] br[200] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_203 
+ bl[201] br[201] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_204 
+ bl[202] br[202] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_205 
+ bl[203] br[203] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_206 
+ bl[204] br[204] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_207 
+ bl[205] br[205] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_208 
+ bl[206] br[206] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_209 
+ bl[207] br[207] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_210 
+ bl[208] br[208] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_211 
+ bl[209] br[209] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_212 
+ bl[210] br[210] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_213 
+ bl[211] br[211] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_214 
+ bl[212] br[212] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_215 
+ bl[213] br[213] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_216 
+ bl[214] br[214] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_217 
+ bl[215] br[215] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_218 
+ bl[216] br[216] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_219 
+ bl[217] br[217] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_220 
+ bl[218] br[218] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_221 
+ bl[219] br[219] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_222 
+ bl[220] br[220] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_223 
+ bl[221] br[221] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_224 
+ bl[222] br[222] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_225 
+ bl[223] br[223] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_226 
+ bl[224] br[224] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_227 
+ bl[225] br[225] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_228 
+ bl[226] br[226] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_229 
+ bl[227] br[227] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_230 
+ bl[228] br[228] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_231 
+ bl[229] br[229] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_232 
+ bl[230] br[230] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_233 
+ bl[231] br[231] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_234 
+ bl[232] br[232] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_235 
+ bl[233] br[233] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_236 
+ bl[234] br[234] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_237 
+ bl[235] br[235] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_238 
+ bl[236] br[236] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_239 
+ bl[237] br[237] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_240 
+ bl[238] br[238] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_241 
+ bl[239] br[239] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_242 
+ bl[240] br[240] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_243 
+ bl[241] br[241] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_244 
+ bl[242] br[242] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_245 
+ bl[243] br[243] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_246 
+ bl[244] br[244] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_247 
+ bl[245] br[245] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_248 
+ bl[246] br[246] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_249 
+ bl[247] br[247] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_250 
+ bl[248] br[248] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_251 
+ bl[249] br[249] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_252 
+ bl[250] br[250] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_253 
+ bl[251] br[251] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_254 
+ bl[252] br[252] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_255 
+ bl[253] br[253] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_256 
+ bl[254] br[254] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_257 
+ bl[255] br[255] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_258 
+ vdd vdd vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_259 
+ vdd vdd vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_0 
+ vdd vdd vss vdd vpb vnb wl[68] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_70_1 
+ rbl rbr vss vdd vpb vnb wl[68] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_70_2 
+ bl[0] br[0] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_3 
+ bl[1] br[1] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_4 
+ bl[2] br[2] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_5 
+ bl[3] br[3] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_6 
+ bl[4] br[4] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_7 
+ bl[5] br[5] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_8 
+ bl[6] br[6] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_9 
+ bl[7] br[7] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_10 
+ bl[8] br[8] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_11 
+ bl[9] br[9] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_12 
+ bl[10] br[10] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_13 
+ bl[11] br[11] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_14 
+ bl[12] br[12] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_15 
+ bl[13] br[13] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_16 
+ bl[14] br[14] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_17 
+ bl[15] br[15] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_18 
+ bl[16] br[16] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_19 
+ bl[17] br[17] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_20 
+ bl[18] br[18] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_21 
+ bl[19] br[19] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_22 
+ bl[20] br[20] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_23 
+ bl[21] br[21] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_24 
+ bl[22] br[22] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_25 
+ bl[23] br[23] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_26 
+ bl[24] br[24] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_27 
+ bl[25] br[25] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_28 
+ bl[26] br[26] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_29 
+ bl[27] br[27] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_30 
+ bl[28] br[28] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_31 
+ bl[29] br[29] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_32 
+ bl[30] br[30] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_33 
+ bl[31] br[31] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_34 
+ bl[32] br[32] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_35 
+ bl[33] br[33] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_36 
+ bl[34] br[34] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_37 
+ bl[35] br[35] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_38 
+ bl[36] br[36] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_39 
+ bl[37] br[37] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_40 
+ bl[38] br[38] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_41 
+ bl[39] br[39] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_42 
+ bl[40] br[40] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_43 
+ bl[41] br[41] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_44 
+ bl[42] br[42] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_45 
+ bl[43] br[43] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_46 
+ bl[44] br[44] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_47 
+ bl[45] br[45] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_48 
+ bl[46] br[46] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_49 
+ bl[47] br[47] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_50 
+ bl[48] br[48] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_51 
+ bl[49] br[49] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_52 
+ bl[50] br[50] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_53 
+ bl[51] br[51] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_54 
+ bl[52] br[52] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_55 
+ bl[53] br[53] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_56 
+ bl[54] br[54] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_57 
+ bl[55] br[55] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_58 
+ bl[56] br[56] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_59 
+ bl[57] br[57] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_60 
+ bl[58] br[58] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_61 
+ bl[59] br[59] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_62 
+ bl[60] br[60] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_63 
+ bl[61] br[61] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_64 
+ bl[62] br[62] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_65 
+ bl[63] br[63] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_66 
+ bl[64] br[64] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_67 
+ bl[65] br[65] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_68 
+ bl[66] br[66] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_69 
+ bl[67] br[67] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_70 
+ bl[68] br[68] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_71 
+ bl[69] br[69] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_72 
+ bl[70] br[70] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_73 
+ bl[71] br[71] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_74 
+ bl[72] br[72] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_75 
+ bl[73] br[73] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_76 
+ bl[74] br[74] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_77 
+ bl[75] br[75] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_78 
+ bl[76] br[76] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_79 
+ bl[77] br[77] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_80 
+ bl[78] br[78] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_81 
+ bl[79] br[79] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_82 
+ bl[80] br[80] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_83 
+ bl[81] br[81] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_84 
+ bl[82] br[82] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_85 
+ bl[83] br[83] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_86 
+ bl[84] br[84] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_87 
+ bl[85] br[85] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_88 
+ bl[86] br[86] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_89 
+ bl[87] br[87] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_90 
+ bl[88] br[88] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_91 
+ bl[89] br[89] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_92 
+ bl[90] br[90] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_93 
+ bl[91] br[91] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_94 
+ bl[92] br[92] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_95 
+ bl[93] br[93] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_96 
+ bl[94] br[94] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_97 
+ bl[95] br[95] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_98 
+ bl[96] br[96] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_99 
+ bl[97] br[97] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_100 
+ bl[98] br[98] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_101 
+ bl[99] br[99] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_102 
+ bl[100] br[100] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_103 
+ bl[101] br[101] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_104 
+ bl[102] br[102] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_105 
+ bl[103] br[103] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_106 
+ bl[104] br[104] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_107 
+ bl[105] br[105] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_108 
+ bl[106] br[106] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_109 
+ bl[107] br[107] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_110 
+ bl[108] br[108] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_111 
+ bl[109] br[109] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_112 
+ bl[110] br[110] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_113 
+ bl[111] br[111] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_114 
+ bl[112] br[112] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_115 
+ bl[113] br[113] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_116 
+ bl[114] br[114] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_117 
+ bl[115] br[115] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_118 
+ bl[116] br[116] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_119 
+ bl[117] br[117] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_120 
+ bl[118] br[118] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_121 
+ bl[119] br[119] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_122 
+ bl[120] br[120] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_123 
+ bl[121] br[121] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_124 
+ bl[122] br[122] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_125 
+ bl[123] br[123] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_126 
+ bl[124] br[124] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_127 
+ bl[125] br[125] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_128 
+ bl[126] br[126] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_129 
+ bl[127] br[127] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_130 
+ bl[128] br[128] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_131 
+ bl[129] br[129] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_132 
+ bl[130] br[130] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_133 
+ bl[131] br[131] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_134 
+ bl[132] br[132] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_135 
+ bl[133] br[133] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_136 
+ bl[134] br[134] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_137 
+ bl[135] br[135] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_138 
+ bl[136] br[136] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_139 
+ bl[137] br[137] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_140 
+ bl[138] br[138] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_141 
+ bl[139] br[139] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_142 
+ bl[140] br[140] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_143 
+ bl[141] br[141] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_144 
+ bl[142] br[142] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_145 
+ bl[143] br[143] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_146 
+ bl[144] br[144] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_147 
+ bl[145] br[145] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_148 
+ bl[146] br[146] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_149 
+ bl[147] br[147] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_150 
+ bl[148] br[148] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_151 
+ bl[149] br[149] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_152 
+ bl[150] br[150] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_153 
+ bl[151] br[151] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_154 
+ bl[152] br[152] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_155 
+ bl[153] br[153] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_156 
+ bl[154] br[154] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_157 
+ bl[155] br[155] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_158 
+ bl[156] br[156] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_159 
+ bl[157] br[157] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_160 
+ bl[158] br[158] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_161 
+ bl[159] br[159] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_162 
+ bl[160] br[160] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_163 
+ bl[161] br[161] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_164 
+ bl[162] br[162] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_165 
+ bl[163] br[163] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_166 
+ bl[164] br[164] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_167 
+ bl[165] br[165] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_168 
+ bl[166] br[166] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_169 
+ bl[167] br[167] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_170 
+ bl[168] br[168] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_171 
+ bl[169] br[169] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_172 
+ bl[170] br[170] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_173 
+ bl[171] br[171] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_174 
+ bl[172] br[172] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_175 
+ bl[173] br[173] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_176 
+ bl[174] br[174] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_177 
+ bl[175] br[175] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_178 
+ bl[176] br[176] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_179 
+ bl[177] br[177] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_180 
+ bl[178] br[178] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_181 
+ bl[179] br[179] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_182 
+ bl[180] br[180] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_183 
+ bl[181] br[181] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_184 
+ bl[182] br[182] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_185 
+ bl[183] br[183] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_186 
+ bl[184] br[184] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_187 
+ bl[185] br[185] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_188 
+ bl[186] br[186] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_189 
+ bl[187] br[187] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_190 
+ bl[188] br[188] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_191 
+ bl[189] br[189] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_192 
+ bl[190] br[190] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_193 
+ bl[191] br[191] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_194 
+ bl[192] br[192] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_195 
+ bl[193] br[193] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_196 
+ bl[194] br[194] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_197 
+ bl[195] br[195] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_198 
+ bl[196] br[196] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_199 
+ bl[197] br[197] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_200 
+ bl[198] br[198] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_201 
+ bl[199] br[199] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_202 
+ bl[200] br[200] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_203 
+ bl[201] br[201] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_204 
+ bl[202] br[202] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_205 
+ bl[203] br[203] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_206 
+ bl[204] br[204] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_207 
+ bl[205] br[205] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_208 
+ bl[206] br[206] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_209 
+ bl[207] br[207] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_210 
+ bl[208] br[208] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_211 
+ bl[209] br[209] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_212 
+ bl[210] br[210] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_213 
+ bl[211] br[211] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_214 
+ bl[212] br[212] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_215 
+ bl[213] br[213] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_216 
+ bl[214] br[214] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_217 
+ bl[215] br[215] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_218 
+ bl[216] br[216] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_219 
+ bl[217] br[217] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_220 
+ bl[218] br[218] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_221 
+ bl[219] br[219] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_222 
+ bl[220] br[220] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_223 
+ bl[221] br[221] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_224 
+ bl[222] br[222] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_225 
+ bl[223] br[223] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_226 
+ bl[224] br[224] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_227 
+ bl[225] br[225] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_228 
+ bl[226] br[226] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_229 
+ bl[227] br[227] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_230 
+ bl[228] br[228] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_231 
+ bl[229] br[229] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_232 
+ bl[230] br[230] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_233 
+ bl[231] br[231] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_234 
+ bl[232] br[232] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_235 
+ bl[233] br[233] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_236 
+ bl[234] br[234] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_237 
+ bl[235] br[235] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_238 
+ bl[236] br[236] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_239 
+ bl[237] br[237] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_240 
+ bl[238] br[238] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_241 
+ bl[239] br[239] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_242 
+ bl[240] br[240] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_243 
+ bl[241] br[241] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_244 
+ bl[242] br[242] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_245 
+ bl[243] br[243] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_246 
+ bl[244] br[244] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_247 
+ bl[245] br[245] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_248 
+ bl[246] br[246] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_249 
+ bl[247] br[247] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_250 
+ bl[248] br[248] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_251 
+ bl[249] br[249] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_252 
+ bl[250] br[250] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_253 
+ bl[251] br[251] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_254 
+ bl[252] br[252] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_255 
+ bl[253] br[253] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_256 
+ bl[254] br[254] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_257 
+ bl[255] br[255] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_258 
+ vdd vdd vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_259 
+ vdd vdd vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_0 
+ vdd vdd vss vdd vpb vnb wl[69] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_71_1 
+ rbl rbr vss vdd vpb vnb wl[69] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_71_2 
+ bl[0] br[0] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_3 
+ bl[1] br[1] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_4 
+ bl[2] br[2] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_5 
+ bl[3] br[3] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_6 
+ bl[4] br[4] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_7 
+ bl[5] br[5] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_8 
+ bl[6] br[6] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_9 
+ bl[7] br[7] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_10 
+ bl[8] br[8] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_11 
+ bl[9] br[9] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_12 
+ bl[10] br[10] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_13 
+ bl[11] br[11] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_14 
+ bl[12] br[12] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_15 
+ bl[13] br[13] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_16 
+ bl[14] br[14] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_17 
+ bl[15] br[15] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_18 
+ bl[16] br[16] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_19 
+ bl[17] br[17] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_20 
+ bl[18] br[18] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_21 
+ bl[19] br[19] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_22 
+ bl[20] br[20] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_23 
+ bl[21] br[21] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_24 
+ bl[22] br[22] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_25 
+ bl[23] br[23] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_26 
+ bl[24] br[24] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_27 
+ bl[25] br[25] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_28 
+ bl[26] br[26] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_29 
+ bl[27] br[27] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_30 
+ bl[28] br[28] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_31 
+ bl[29] br[29] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_32 
+ bl[30] br[30] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_33 
+ bl[31] br[31] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_34 
+ bl[32] br[32] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_35 
+ bl[33] br[33] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_36 
+ bl[34] br[34] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_37 
+ bl[35] br[35] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_38 
+ bl[36] br[36] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_39 
+ bl[37] br[37] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_40 
+ bl[38] br[38] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_41 
+ bl[39] br[39] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_42 
+ bl[40] br[40] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_43 
+ bl[41] br[41] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_44 
+ bl[42] br[42] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_45 
+ bl[43] br[43] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_46 
+ bl[44] br[44] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_47 
+ bl[45] br[45] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_48 
+ bl[46] br[46] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_49 
+ bl[47] br[47] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_50 
+ bl[48] br[48] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_51 
+ bl[49] br[49] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_52 
+ bl[50] br[50] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_53 
+ bl[51] br[51] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_54 
+ bl[52] br[52] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_55 
+ bl[53] br[53] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_56 
+ bl[54] br[54] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_57 
+ bl[55] br[55] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_58 
+ bl[56] br[56] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_59 
+ bl[57] br[57] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_60 
+ bl[58] br[58] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_61 
+ bl[59] br[59] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_62 
+ bl[60] br[60] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_63 
+ bl[61] br[61] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_64 
+ bl[62] br[62] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_65 
+ bl[63] br[63] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_66 
+ bl[64] br[64] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_67 
+ bl[65] br[65] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_68 
+ bl[66] br[66] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_69 
+ bl[67] br[67] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_70 
+ bl[68] br[68] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_71 
+ bl[69] br[69] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_72 
+ bl[70] br[70] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_73 
+ bl[71] br[71] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_74 
+ bl[72] br[72] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_75 
+ bl[73] br[73] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_76 
+ bl[74] br[74] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_77 
+ bl[75] br[75] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_78 
+ bl[76] br[76] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_79 
+ bl[77] br[77] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_80 
+ bl[78] br[78] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_81 
+ bl[79] br[79] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_82 
+ bl[80] br[80] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_83 
+ bl[81] br[81] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_84 
+ bl[82] br[82] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_85 
+ bl[83] br[83] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_86 
+ bl[84] br[84] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_87 
+ bl[85] br[85] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_88 
+ bl[86] br[86] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_89 
+ bl[87] br[87] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_90 
+ bl[88] br[88] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_91 
+ bl[89] br[89] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_92 
+ bl[90] br[90] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_93 
+ bl[91] br[91] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_94 
+ bl[92] br[92] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_95 
+ bl[93] br[93] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_96 
+ bl[94] br[94] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_97 
+ bl[95] br[95] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_98 
+ bl[96] br[96] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_99 
+ bl[97] br[97] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_100 
+ bl[98] br[98] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_101 
+ bl[99] br[99] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_102 
+ bl[100] br[100] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_103 
+ bl[101] br[101] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_104 
+ bl[102] br[102] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_105 
+ bl[103] br[103] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_106 
+ bl[104] br[104] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_107 
+ bl[105] br[105] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_108 
+ bl[106] br[106] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_109 
+ bl[107] br[107] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_110 
+ bl[108] br[108] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_111 
+ bl[109] br[109] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_112 
+ bl[110] br[110] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_113 
+ bl[111] br[111] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_114 
+ bl[112] br[112] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_115 
+ bl[113] br[113] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_116 
+ bl[114] br[114] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_117 
+ bl[115] br[115] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_118 
+ bl[116] br[116] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_119 
+ bl[117] br[117] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_120 
+ bl[118] br[118] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_121 
+ bl[119] br[119] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_122 
+ bl[120] br[120] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_123 
+ bl[121] br[121] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_124 
+ bl[122] br[122] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_125 
+ bl[123] br[123] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_126 
+ bl[124] br[124] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_127 
+ bl[125] br[125] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_128 
+ bl[126] br[126] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_129 
+ bl[127] br[127] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_130 
+ bl[128] br[128] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_131 
+ bl[129] br[129] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_132 
+ bl[130] br[130] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_133 
+ bl[131] br[131] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_134 
+ bl[132] br[132] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_135 
+ bl[133] br[133] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_136 
+ bl[134] br[134] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_137 
+ bl[135] br[135] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_138 
+ bl[136] br[136] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_139 
+ bl[137] br[137] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_140 
+ bl[138] br[138] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_141 
+ bl[139] br[139] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_142 
+ bl[140] br[140] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_143 
+ bl[141] br[141] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_144 
+ bl[142] br[142] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_145 
+ bl[143] br[143] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_146 
+ bl[144] br[144] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_147 
+ bl[145] br[145] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_148 
+ bl[146] br[146] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_149 
+ bl[147] br[147] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_150 
+ bl[148] br[148] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_151 
+ bl[149] br[149] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_152 
+ bl[150] br[150] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_153 
+ bl[151] br[151] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_154 
+ bl[152] br[152] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_155 
+ bl[153] br[153] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_156 
+ bl[154] br[154] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_157 
+ bl[155] br[155] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_158 
+ bl[156] br[156] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_159 
+ bl[157] br[157] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_160 
+ bl[158] br[158] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_161 
+ bl[159] br[159] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_162 
+ bl[160] br[160] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_163 
+ bl[161] br[161] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_164 
+ bl[162] br[162] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_165 
+ bl[163] br[163] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_166 
+ bl[164] br[164] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_167 
+ bl[165] br[165] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_168 
+ bl[166] br[166] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_169 
+ bl[167] br[167] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_170 
+ bl[168] br[168] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_171 
+ bl[169] br[169] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_172 
+ bl[170] br[170] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_173 
+ bl[171] br[171] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_174 
+ bl[172] br[172] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_175 
+ bl[173] br[173] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_176 
+ bl[174] br[174] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_177 
+ bl[175] br[175] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_178 
+ bl[176] br[176] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_179 
+ bl[177] br[177] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_180 
+ bl[178] br[178] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_181 
+ bl[179] br[179] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_182 
+ bl[180] br[180] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_183 
+ bl[181] br[181] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_184 
+ bl[182] br[182] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_185 
+ bl[183] br[183] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_186 
+ bl[184] br[184] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_187 
+ bl[185] br[185] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_188 
+ bl[186] br[186] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_189 
+ bl[187] br[187] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_190 
+ bl[188] br[188] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_191 
+ bl[189] br[189] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_192 
+ bl[190] br[190] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_193 
+ bl[191] br[191] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_194 
+ bl[192] br[192] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_195 
+ bl[193] br[193] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_196 
+ bl[194] br[194] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_197 
+ bl[195] br[195] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_198 
+ bl[196] br[196] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_199 
+ bl[197] br[197] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_200 
+ bl[198] br[198] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_201 
+ bl[199] br[199] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_202 
+ bl[200] br[200] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_203 
+ bl[201] br[201] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_204 
+ bl[202] br[202] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_205 
+ bl[203] br[203] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_206 
+ bl[204] br[204] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_207 
+ bl[205] br[205] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_208 
+ bl[206] br[206] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_209 
+ bl[207] br[207] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_210 
+ bl[208] br[208] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_211 
+ bl[209] br[209] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_212 
+ bl[210] br[210] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_213 
+ bl[211] br[211] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_214 
+ bl[212] br[212] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_215 
+ bl[213] br[213] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_216 
+ bl[214] br[214] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_217 
+ bl[215] br[215] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_218 
+ bl[216] br[216] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_219 
+ bl[217] br[217] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_220 
+ bl[218] br[218] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_221 
+ bl[219] br[219] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_222 
+ bl[220] br[220] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_223 
+ bl[221] br[221] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_224 
+ bl[222] br[222] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_225 
+ bl[223] br[223] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_226 
+ bl[224] br[224] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_227 
+ bl[225] br[225] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_228 
+ bl[226] br[226] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_229 
+ bl[227] br[227] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_230 
+ bl[228] br[228] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_231 
+ bl[229] br[229] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_232 
+ bl[230] br[230] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_233 
+ bl[231] br[231] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_234 
+ bl[232] br[232] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_235 
+ bl[233] br[233] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_236 
+ bl[234] br[234] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_237 
+ bl[235] br[235] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_238 
+ bl[236] br[236] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_239 
+ bl[237] br[237] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_240 
+ bl[238] br[238] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_241 
+ bl[239] br[239] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_242 
+ bl[240] br[240] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_243 
+ bl[241] br[241] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_244 
+ bl[242] br[242] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_245 
+ bl[243] br[243] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_246 
+ bl[244] br[244] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_247 
+ bl[245] br[245] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_248 
+ bl[246] br[246] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_249 
+ bl[247] br[247] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_250 
+ bl[248] br[248] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_251 
+ bl[249] br[249] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_252 
+ bl[250] br[250] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_253 
+ bl[251] br[251] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_254 
+ bl[252] br[252] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_255 
+ bl[253] br[253] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_256 
+ bl[254] br[254] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_257 
+ bl[255] br[255] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_258 
+ vdd vdd vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_259 
+ vdd vdd vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_0 
+ vdd vdd vss vdd vpb vnb wl[70] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_72_1 
+ rbl rbr vss vdd vpb vnb wl[70] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_72_2 
+ bl[0] br[0] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_3 
+ bl[1] br[1] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_4 
+ bl[2] br[2] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_5 
+ bl[3] br[3] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_6 
+ bl[4] br[4] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_7 
+ bl[5] br[5] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_8 
+ bl[6] br[6] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_9 
+ bl[7] br[7] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_10 
+ bl[8] br[8] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_11 
+ bl[9] br[9] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_12 
+ bl[10] br[10] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_13 
+ bl[11] br[11] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_14 
+ bl[12] br[12] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_15 
+ bl[13] br[13] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_16 
+ bl[14] br[14] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_17 
+ bl[15] br[15] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_18 
+ bl[16] br[16] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_19 
+ bl[17] br[17] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_20 
+ bl[18] br[18] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_21 
+ bl[19] br[19] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_22 
+ bl[20] br[20] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_23 
+ bl[21] br[21] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_24 
+ bl[22] br[22] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_25 
+ bl[23] br[23] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_26 
+ bl[24] br[24] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_27 
+ bl[25] br[25] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_28 
+ bl[26] br[26] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_29 
+ bl[27] br[27] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_30 
+ bl[28] br[28] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_31 
+ bl[29] br[29] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_32 
+ bl[30] br[30] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_33 
+ bl[31] br[31] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_34 
+ bl[32] br[32] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_35 
+ bl[33] br[33] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_36 
+ bl[34] br[34] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_37 
+ bl[35] br[35] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_38 
+ bl[36] br[36] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_39 
+ bl[37] br[37] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_40 
+ bl[38] br[38] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_41 
+ bl[39] br[39] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_42 
+ bl[40] br[40] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_43 
+ bl[41] br[41] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_44 
+ bl[42] br[42] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_45 
+ bl[43] br[43] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_46 
+ bl[44] br[44] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_47 
+ bl[45] br[45] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_48 
+ bl[46] br[46] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_49 
+ bl[47] br[47] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_50 
+ bl[48] br[48] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_51 
+ bl[49] br[49] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_52 
+ bl[50] br[50] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_53 
+ bl[51] br[51] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_54 
+ bl[52] br[52] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_55 
+ bl[53] br[53] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_56 
+ bl[54] br[54] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_57 
+ bl[55] br[55] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_58 
+ bl[56] br[56] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_59 
+ bl[57] br[57] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_60 
+ bl[58] br[58] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_61 
+ bl[59] br[59] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_62 
+ bl[60] br[60] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_63 
+ bl[61] br[61] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_64 
+ bl[62] br[62] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_65 
+ bl[63] br[63] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_66 
+ bl[64] br[64] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_67 
+ bl[65] br[65] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_68 
+ bl[66] br[66] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_69 
+ bl[67] br[67] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_70 
+ bl[68] br[68] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_71 
+ bl[69] br[69] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_72 
+ bl[70] br[70] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_73 
+ bl[71] br[71] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_74 
+ bl[72] br[72] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_75 
+ bl[73] br[73] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_76 
+ bl[74] br[74] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_77 
+ bl[75] br[75] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_78 
+ bl[76] br[76] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_79 
+ bl[77] br[77] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_80 
+ bl[78] br[78] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_81 
+ bl[79] br[79] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_82 
+ bl[80] br[80] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_83 
+ bl[81] br[81] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_84 
+ bl[82] br[82] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_85 
+ bl[83] br[83] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_86 
+ bl[84] br[84] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_87 
+ bl[85] br[85] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_88 
+ bl[86] br[86] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_89 
+ bl[87] br[87] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_90 
+ bl[88] br[88] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_91 
+ bl[89] br[89] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_92 
+ bl[90] br[90] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_93 
+ bl[91] br[91] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_94 
+ bl[92] br[92] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_95 
+ bl[93] br[93] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_96 
+ bl[94] br[94] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_97 
+ bl[95] br[95] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_98 
+ bl[96] br[96] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_99 
+ bl[97] br[97] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_100 
+ bl[98] br[98] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_101 
+ bl[99] br[99] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_102 
+ bl[100] br[100] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_103 
+ bl[101] br[101] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_104 
+ bl[102] br[102] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_105 
+ bl[103] br[103] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_106 
+ bl[104] br[104] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_107 
+ bl[105] br[105] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_108 
+ bl[106] br[106] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_109 
+ bl[107] br[107] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_110 
+ bl[108] br[108] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_111 
+ bl[109] br[109] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_112 
+ bl[110] br[110] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_113 
+ bl[111] br[111] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_114 
+ bl[112] br[112] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_115 
+ bl[113] br[113] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_116 
+ bl[114] br[114] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_117 
+ bl[115] br[115] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_118 
+ bl[116] br[116] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_119 
+ bl[117] br[117] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_120 
+ bl[118] br[118] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_121 
+ bl[119] br[119] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_122 
+ bl[120] br[120] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_123 
+ bl[121] br[121] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_124 
+ bl[122] br[122] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_125 
+ bl[123] br[123] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_126 
+ bl[124] br[124] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_127 
+ bl[125] br[125] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_128 
+ bl[126] br[126] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_129 
+ bl[127] br[127] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_130 
+ bl[128] br[128] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_131 
+ bl[129] br[129] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_132 
+ bl[130] br[130] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_133 
+ bl[131] br[131] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_134 
+ bl[132] br[132] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_135 
+ bl[133] br[133] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_136 
+ bl[134] br[134] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_137 
+ bl[135] br[135] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_138 
+ bl[136] br[136] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_139 
+ bl[137] br[137] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_140 
+ bl[138] br[138] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_141 
+ bl[139] br[139] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_142 
+ bl[140] br[140] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_143 
+ bl[141] br[141] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_144 
+ bl[142] br[142] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_145 
+ bl[143] br[143] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_146 
+ bl[144] br[144] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_147 
+ bl[145] br[145] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_148 
+ bl[146] br[146] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_149 
+ bl[147] br[147] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_150 
+ bl[148] br[148] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_151 
+ bl[149] br[149] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_152 
+ bl[150] br[150] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_153 
+ bl[151] br[151] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_154 
+ bl[152] br[152] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_155 
+ bl[153] br[153] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_156 
+ bl[154] br[154] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_157 
+ bl[155] br[155] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_158 
+ bl[156] br[156] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_159 
+ bl[157] br[157] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_160 
+ bl[158] br[158] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_161 
+ bl[159] br[159] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_162 
+ bl[160] br[160] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_163 
+ bl[161] br[161] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_164 
+ bl[162] br[162] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_165 
+ bl[163] br[163] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_166 
+ bl[164] br[164] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_167 
+ bl[165] br[165] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_168 
+ bl[166] br[166] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_169 
+ bl[167] br[167] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_170 
+ bl[168] br[168] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_171 
+ bl[169] br[169] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_172 
+ bl[170] br[170] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_173 
+ bl[171] br[171] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_174 
+ bl[172] br[172] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_175 
+ bl[173] br[173] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_176 
+ bl[174] br[174] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_177 
+ bl[175] br[175] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_178 
+ bl[176] br[176] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_179 
+ bl[177] br[177] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_180 
+ bl[178] br[178] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_181 
+ bl[179] br[179] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_182 
+ bl[180] br[180] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_183 
+ bl[181] br[181] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_184 
+ bl[182] br[182] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_185 
+ bl[183] br[183] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_186 
+ bl[184] br[184] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_187 
+ bl[185] br[185] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_188 
+ bl[186] br[186] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_189 
+ bl[187] br[187] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_190 
+ bl[188] br[188] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_191 
+ bl[189] br[189] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_192 
+ bl[190] br[190] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_193 
+ bl[191] br[191] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_194 
+ bl[192] br[192] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_195 
+ bl[193] br[193] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_196 
+ bl[194] br[194] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_197 
+ bl[195] br[195] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_198 
+ bl[196] br[196] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_199 
+ bl[197] br[197] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_200 
+ bl[198] br[198] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_201 
+ bl[199] br[199] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_202 
+ bl[200] br[200] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_203 
+ bl[201] br[201] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_204 
+ bl[202] br[202] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_205 
+ bl[203] br[203] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_206 
+ bl[204] br[204] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_207 
+ bl[205] br[205] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_208 
+ bl[206] br[206] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_209 
+ bl[207] br[207] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_210 
+ bl[208] br[208] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_211 
+ bl[209] br[209] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_212 
+ bl[210] br[210] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_213 
+ bl[211] br[211] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_214 
+ bl[212] br[212] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_215 
+ bl[213] br[213] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_216 
+ bl[214] br[214] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_217 
+ bl[215] br[215] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_218 
+ bl[216] br[216] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_219 
+ bl[217] br[217] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_220 
+ bl[218] br[218] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_221 
+ bl[219] br[219] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_222 
+ bl[220] br[220] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_223 
+ bl[221] br[221] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_224 
+ bl[222] br[222] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_225 
+ bl[223] br[223] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_226 
+ bl[224] br[224] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_227 
+ bl[225] br[225] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_228 
+ bl[226] br[226] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_229 
+ bl[227] br[227] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_230 
+ bl[228] br[228] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_231 
+ bl[229] br[229] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_232 
+ bl[230] br[230] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_233 
+ bl[231] br[231] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_234 
+ bl[232] br[232] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_235 
+ bl[233] br[233] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_236 
+ bl[234] br[234] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_237 
+ bl[235] br[235] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_238 
+ bl[236] br[236] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_239 
+ bl[237] br[237] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_240 
+ bl[238] br[238] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_241 
+ bl[239] br[239] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_242 
+ bl[240] br[240] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_243 
+ bl[241] br[241] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_244 
+ bl[242] br[242] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_245 
+ bl[243] br[243] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_246 
+ bl[244] br[244] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_247 
+ bl[245] br[245] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_248 
+ bl[246] br[246] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_249 
+ bl[247] br[247] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_250 
+ bl[248] br[248] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_251 
+ bl[249] br[249] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_252 
+ bl[250] br[250] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_253 
+ bl[251] br[251] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_254 
+ bl[252] br[252] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_255 
+ bl[253] br[253] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_256 
+ bl[254] br[254] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_257 
+ bl[255] br[255] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_258 
+ vdd vdd vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_259 
+ vdd vdd vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_0 
+ vdd vdd vss vdd vpb vnb wl[71] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_73_1 
+ rbl rbr vss vdd vpb vnb wl[71] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_73_2 
+ bl[0] br[0] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_3 
+ bl[1] br[1] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_4 
+ bl[2] br[2] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_5 
+ bl[3] br[3] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_6 
+ bl[4] br[4] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_7 
+ bl[5] br[5] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_8 
+ bl[6] br[6] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_9 
+ bl[7] br[7] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_10 
+ bl[8] br[8] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_11 
+ bl[9] br[9] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_12 
+ bl[10] br[10] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_13 
+ bl[11] br[11] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_14 
+ bl[12] br[12] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_15 
+ bl[13] br[13] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_16 
+ bl[14] br[14] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_17 
+ bl[15] br[15] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_18 
+ bl[16] br[16] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_19 
+ bl[17] br[17] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_20 
+ bl[18] br[18] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_21 
+ bl[19] br[19] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_22 
+ bl[20] br[20] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_23 
+ bl[21] br[21] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_24 
+ bl[22] br[22] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_25 
+ bl[23] br[23] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_26 
+ bl[24] br[24] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_27 
+ bl[25] br[25] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_28 
+ bl[26] br[26] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_29 
+ bl[27] br[27] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_30 
+ bl[28] br[28] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_31 
+ bl[29] br[29] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_32 
+ bl[30] br[30] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_33 
+ bl[31] br[31] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_34 
+ bl[32] br[32] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_35 
+ bl[33] br[33] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_36 
+ bl[34] br[34] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_37 
+ bl[35] br[35] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_38 
+ bl[36] br[36] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_39 
+ bl[37] br[37] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_40 
+ bl[38] br[38] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_41 
+ bl[39] br[39] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_42 
+ bl[40] br[40] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_43 
+ bl[41] br[41] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_44 
+ bl[42] br[42] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_45 
+ bl[43] br[43] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_46 
+ bl[44] br[44] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_47 
+ bl[45] br[45] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_48 
+ bl[46] br[46] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_49 
+ bl[47] br[47] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_50 
+ bl[48] br[48] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_51 
+ bl[49] br[49] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_52 
+ bl[50] br[50] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_53 
+ bl[51] br[51] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_54 
+ bl[52] br[52] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_55 
+ bl[53] br[53] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_56 
+ bl[54] br[54] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_57 
+ bl[55] br[55] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_58 
+ bl[56] br[56] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_59 
+ bl[57] br[57] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_60 
+ bl[58] br[58] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_61 
+ bl[59] br[59] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_62 
+ bl[60] br[60] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_63 
+ bl[61] br[61] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_64 
+ bl[62] br[62] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_65 
+ bl[63] br[63] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_66 
+ bl[64] br[64] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_67 
+ bl[65] br[65] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_68 
+ bl[66] br[66] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_69 
+ bl[67] br[67] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_70 
+ bl[68] br[68] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_71 
+ bl[69] br[69] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_72 
+ bl[70] br[70] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_73 
+ bl[71] br[71] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_74 
+ bl[72] br[72] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_75 
+ bl[73] br[73] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_76 
+ bl[74] br[74] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_77 
+ bl[75] br[75] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_78 
+ bl[76] br[76] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_79 
+ bl[77] br[77] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_80 
+ bl[78] br[78] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_81 
+ bl[79] br[79] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_82 
+ bl[80] br[80] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_83 
+ bl[81] br[81] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_84 
+ bl[82] br[82] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_85 
+ bl[83] br[83] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_86 
+ bl[84] br[84] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_87 
+ bl[85] br[85] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_88 
+ bl[86] br[86] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_89 
+ bl[87] br[87] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_90 
+ bl[88] br[88] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_91 
+ bl[89] br[89] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_92 
+ bl[90] br[90] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_93 
+ bl[91] br[91] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_94 
+ bl[92] br[92] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_95 
+ bl[93] br[93] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_96 
+ bl[94] br[94] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_97 
+ bl[95] br[95] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_98 
+ bl[96] br[96] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_99 
+ bl[97] br[97] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_100 
+ bl[98] br[98] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_101 
+ bl[99] br[99] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_102 
+ bl[100] br[100] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_103 
+ bl[101] br[101] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_104 
+ bl[102] br[102] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_105 
+ bl[103] br[103] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_106 
+ bl[104] br[104] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_107 
+ bl[105] br[105] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_108 
+ bl[106] br[106] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_109 
+ bl[107] br[107] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_110 
+ bl[108] br[108] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_111 
+ bl[109] br[109] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_112 
+ bl[110] br[110] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_113 
+ bl[111] br[111] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_114 
+ bl[112] br[112] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_115 
+ bl[113] br[113] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_116 
+ bl[114] br[114] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_117 
+ bl[115] br[115] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_118 
+ bl[116] br[116] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_119 
+ bl[117] br[117] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_120 
+ bl[118] br[118] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_121 
+ bl[119] br[119] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_122 
+ bl[120] br[120] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_123 
+ bl[121] br[121] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_124 
+ bl[122] br[122] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_125 
+ bl[123] br[123] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_126 
+ bl[124] br[124] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_127 
+ bl[125] br[125] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_128 
+ bl[126] br[126] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_129 
+ bl[127] br[127] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_130 
+ bl[128] br[128] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_131 
+ bl[129] br[129] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_132 
+ bl[130] br[130] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_133 
+ bl[131] br[131] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_134 
+ bl[132] br[132] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_135 
+ bl[133] br[133] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_136 
+ bl[134] br[134] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_137 
+ bl[135] br[135] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_138 
+ bl[136] br[136] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_139 
+ bl[137] br[137] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_140 
+ bl[138] br[138] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_141 
+ bl[139] br[139] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_142 
+ bl[140] br[140] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_143 
+ bl[141] br[141] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_144 
+ bl[142] br[142] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_145 
+ bl[143] br[143] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_146 
+ bl[144] br[144] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_147 
+ bl[145] br[145] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_148 
+ bl[146] br[146] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_149 
+ bl[147] br[147] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_150 
+ bl[148] br[148] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_151 
+ bl[149] br[149] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_152 
+ bl[150] br[150] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_153 
+ bl[151] br[151] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_154 
+ bl[152] br[152] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_155 
+ bl[153] br[153] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_156 
+ bl[154] br[154] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_157 
+ bl[155] br[155] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_158 
+ bl[156] br[156] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_159 
+ bl[157] br[157] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_160 
+ bl[158] br[158] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_161 
+ bl[159] br[159] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_162 
+ bl[160] br[160] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_163 
+ bl[161] br[161] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_164 
+ bl[162] br[162] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_165 
+ bl[163] br[163] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_166 
+ bl[164] br[164] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_167 
+ bl[165] br[165] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_168 
+ bl[166] br[166] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_169 
+ bl[167] br[167] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_170 
+ bl[168] br[168] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_171 
+ bl[169] br[169] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_172 
+ bl[170] br[170] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_173 
+ bl[171] br[171] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_174 
+ bl[172] br[172] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_175 
+ bl[173] br[173] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_176 
+ bl[174] br[174] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_177 
+ bl[175] br[175] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_178 
+ bl[176] br[176] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_179 
+ bl[177] br[177] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_180 
+ bl[178] br[178] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_181 
+ bl[179] br[179] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_182 
+ bl[180] br[180] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_183 
+ bl[181] br[181] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_184 
+ bl[182] br[182] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_185 
+ bl[183] br[183] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_186 
+ bl[184] br[184] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_187 
+ bl[185] br[185] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_188 
+ bl[186] br[186] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_189 
+ bl[187] br[187] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_190 
+ bl[188] br[188] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_191 
+ bl[189] br[189] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_192 
+ bl[190] br[190] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_193 
+ bl[191] br[191] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_194 
+ bl[192] br[192] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_195 
+ bl[193] br[193] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_196 
+ bl[194] br[194] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_197 
+ bl[195] br[195] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_198 
+ bl[196] br[196] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_199 
+ bl[197] br[197] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_200 
+ bl[198] br[198] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_201 
+ bl[199] br[199] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_202 
+ bl[200] br[200] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_203 
+ bl[201] br[201] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_204 
+ bl[202] br[202] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_205 
+ bl[203] br[203] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_206 
+ bl[204] br[204] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_207 
+ bl[205] br[205] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_208 
+ bl[206] br[206] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_209 
+ bl[207] br[207] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_210 
+ bl[208] br[208] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_211 
+ bl[209] br[209] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_212 
+ bl[210] br[210] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_213 
+ bl[211] br[211] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_214 
+ bl[212] br[212] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_215 
+ bl[213] br[213] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_216 
+ bl[214] br[214] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_217 
+ bl[215] br[215] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_218 
+ bl[216] br[216] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_219 
+ bl[217] br[217] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_220 
+ bl[218] br[218] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_221 
+ bl[219] br[219] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_222 
+ bl[220] br[220] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_223 
+ bl[221] br[221] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_224 
+ bl[222] br[222] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_225 
+ bl[223] br[223] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_226 
+ bl[224] br[224] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_227 
+ bl[225] br[225] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_228 
+ bl[226] br[226] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_229 
+ bl[227] br[227] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_230 
+ bl[228] br[228] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_231 
+ bl[229] br[229] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_232 
+ bl[230] br[230] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_233 
+ bl[231] br[231] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_234 
+ bl[232] br[232] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_235 
+ bl[233] br[233] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_236 
+ bl[234] br[234] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_237 
+ bl[235] br[235] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_238 
+ bl[236] br[236] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_239 
+ bl[237] br[237] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_240 
+ bl[238] br[238] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_241 
+ bl[239] br[239] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_242 
+ bl[240] br[240] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_243 
+ bl[241] br[241] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_244 
+ bl[242] br[242] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_245 
+ bl[243] br[243] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_246 
+ bl[244] br[244] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_247 
+ bl[245] br[245] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_248 
+ bl[246] br[246] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_249 
+ bl[247] br[247] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_250 
+ bl[248] br[248] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_251 
+ bl[249] br[249] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_252 
+ bl[250] br[250] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_253 
+ bl[251] br[251] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_254 
+ bl[252] br[252] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_255 
+ bl[253] br[253] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_256 
+ bl[254] br[254] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_257 
+ bl[255] br[255] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_258 
+ vdd vdd vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_259 
+ vdd vdd vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_0 
+ vdd vdd vss vdd vpb vnb wl[72] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_74_1 
+ rbl rbr vss vdd vpb vnb wl[72] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_74_2 
+ bl[0] br[0] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_3 
+ bl[1] br[1] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_4 
+ bl[2] br[2] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_5 
+ bl[3] br[3] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_6 
+ bl[4] br[4] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_7 
+ bl[5] br[5] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_8 
+ bl[6] br[6] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_9 
+ bl[7] br[7] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_10 
+ bl[8] br[8] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_11 
+ bl[9] br[9] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_12 
+ bl[10] br[10] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_13 
+ bl[11] br[11] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_14 
+ bl[12] br[12] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_15 
+ bl[13] br[13] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_16 
+ bl[14] br[14] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_17 
+ bl[15] br[15] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_18 
+ bl[16] br[16] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_19 
+ bl[17] br[17] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_20 
+ bl[18] br[18] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_21 
+ bl[19] br[19] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_22 
+ bl[20] br[20] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_23 
+ bl[21] br[21] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_24 
+ bl[22] br[22] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_25 
+ bl[23] br[23] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_26 
+ bl[24] br[24] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_27 
+ bl[25] br[25] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_28 
+ bl[26] br[26] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_29 
+ bl[27] br[27] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_30 
+ bl[28] br[28] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_31 
+ bl[29] br[29] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_32 
+ bl[30] br[30] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_33 
+ bl[31] br[31] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_34 
+ bl[32] br[32] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_35 
+ bl[33] br[33] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_36 
+ bl[34] br[34] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_37 
+ bl[35] br[35] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_38 
+ bl[36] br[36] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_39 
+ bl[37] br[37] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_40 
+ bl[38] br[38] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_41 
+ bl[39] br[39] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_42 
+ bl[40] br[40] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_43 
+ bl[41] br[41] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_44 
+ bl[42] br[42] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_45 
+ bl[43] br[43] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_46 
+ bl[44] br[44] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_47 
+ bl[45] br[45] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_48 
+ bl[46] br[46] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_49 
+ bl[47] br[47] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_50 
+ bl[48] br[48] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_51 
+ bl[49] br[49] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_52 
+ bl[50] br[50] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_53 
+ bl[51] br[51] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_54 
+ bl[52] br[52] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_55 
+ bl[53] br[53] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_56 
+ bl[54] br[54] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_57 
+ bl[55] br[55] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_58 
+ bl[56] br[56] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_59 
+ bl[57] br[57] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_60 
+ bl[58] br[58] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_61 
+ bl[59] br[59] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_62 
+ bl[60] br[60] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_63 
+ bl[61] br[61] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_64 
+ bl[62] br[62] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_65 
+ bl[63] br[63] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_66 
+ bl[64] br[64] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_67 
+ bl[65] br[65] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_68 
+ bl[66] br[66] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_69 
+ bl[67] br[67] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_70 
+ bl[68] br[68] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_71 
+ bl[69] br[69] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_72 
+ bl[70] br[70] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_73 
+ bl[71] br[71] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_74 
+ bl[72] br[72] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_75 
+ bl[73] br[73] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_76 
+ bl[74] br[74] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_77 
+ bl[75] br[75] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_78 
+ bl[76] br[76] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_79 
+ bl[77] br[77] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_80 
+ bl[78] br[78] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_81 
+ bl[79] br[79] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_82 
+ bl[80] br[80] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_83 
+ bl[81] br[81] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_84 
+ bl[82] br[82] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_85 
+ bl[83] br[83] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_86 
+ bl[84] br[84] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_87 
+ bl[85] br[85] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_88 
+ bl[86] br[86] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_89 
+ bl[87] br[87] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_90 
+ bl[88] br[88] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_91 
+ bl[89] br[89] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_92 
+ bl[90] br[90] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_93 
+ bl[91] br[91] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_94 
+ bl[92] br[92] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_95 
+ bl[93] br[93] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_96 
+ bl[94] br[94] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_97 
+ bl[95] br[95] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_98 
+ bl[96] br[96] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_99 
+ bl[97] br[97] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_100 
+ bl[98] br[98] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_101 
+ bl[99] br[99] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_102 
+ bl[100] br[100] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_103 
+ bl[101] br[101] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_104 
+ bl[102] br[102] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_105 
+ bl[103] br[103] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_106 
+ bl[104] br[104] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_107 
+ bl[105] br[105] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_108 
+ bl[106] br[106] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_109 
+ bl[107] br[107] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_110 
+ bl[108] br[108] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_111 
+ bl[109] br[109] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_112 
+ bl[110] br[110] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_113 
+ bl[111] br[111] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_114 
+ bl[112] br[112] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_115 
+ bl[113] br[113] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_116 
+ bl[114] br[114] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_117 
+ bl[115] br[115] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_118 
+ bl[116] br[116] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_119 
+ bl[117] br[117] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_120 
+ bl[118] br[118] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_121 
+ bl[119] br[119] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_122 
+ bl[120] br[120] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_123 
+ bl[121] br[121] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_124 
+ bl[122] br[122] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_125 
+ bl[123] br[123] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_126 
+ bl[124] br[124] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_127 
+ bl[125] br[125] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_128 
+ bl[126] br[126] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_129 
+ bl[127] br[127] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_130 
+ bl[128] br[128] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_131 
+ bl[129] br[129] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_132 
+ bl[130] br[130] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_133 
+ bl[131] br[131] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_134 
+ bl[132] br[132] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_135 
+ bl[133] br[133] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_136 
+ bl[134] br[134] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_137 
+ bl[135] br[135] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_138 
+ bl[136] br[136] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_139 
+ bl[137] br[137] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_140 
+ bl[138] br[138] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_141 
+ bl[139] br[139] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_142 
+ bl[140] br[140] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_143 
+ bl[141] br[141] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_144 
+ bl[142] br[142] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_145 
+ bl[143] br[143] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_146 
+ bl[144] br[144] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_147 
+ bl[145] br[145] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_148 
+ bl[146] br[146] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_149 
+ bl[147] br[147] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_150 
+ bl[148] br[148] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_151 
+ bl[149] br[149] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_152 
+ bl[150] br[150] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_153 
+ bl[151] br[151] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_154 
+ bl[152] br[152] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_155 
+ bl[153] br[153] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_156 
+ bl[154] br[154] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_157 
+ bl[155] br[155] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_158 
+ bl[156] br[156] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_159 
+ bl[157] br[157] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_160 
+ bl[158] br[158] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_161 
+ bl[159] br[159] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_162 
+ bl[160] br[160] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_163 
+ bl[161] br[161] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_164 
+ bl[162] br[162] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_165 
+ bl[163] br[163] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_166 
+ bl[164] br[164] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_167 
+ bl[165] br[165] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_168 
+ bl[166] br[166] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_169 
+ bl[167] br[167] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_170 
+ bl[168] br[168] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_171 
+ bl[169] br[169] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_172 
+ bl[170] br[170] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_173 
+ bl[171] br[171] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_174 
+ bl[172] br[172] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_175 
+ bl[173] br[173] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_176 
+ bl[174] br[174] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_177 
+ bl[175] br[175] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_178 
+ bl[176] br[176] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_179 
+ bl[177] br[177] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_180 
+ bl[178] br[178] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_181 
+ bl[179] br[179] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_182 
+ bl[180] br[180] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_183 
+ bl[181] br[181] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_184 
+ bl[182] br[182] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_185 
+ bl[183] br[183] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_186 
+ bl[184] br[184] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_187 
+ bl[185] br[185] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_188 
+ bl[186] br[186] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_189 
+ bl[187] br[187] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_190 
+ bl[188] br[188] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_191 
+ bl[189] br[189] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_192 
+ bl[190] br[190] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_193 
+ bl[191] br[191] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_194 
+ bl[192] br[192] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_195 
+ bl[193] br[193] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_196 
+ bl[194] br[194] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_197 
+ bl[195] br[195] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_198 
+ bl[196] br[196] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_199 
+ bl[197] br[197] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_200 
+ bl[198] br[198] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_201 
+ bl[199] br[199] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_202 
+ bl[200] br[200] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_203 
+ bl[201] br[201] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_204 
+ bl[202] br[202] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_205 
+ bl[203] br[203] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_206 
+ bl[204] br[204] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_207 
+ bl[205] br[205] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_208 
+ bl[206] br[206] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_209 
+ bl[207] br[207] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_210 
+ bl[208] br[208] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_211 
+ bl[209] br[209] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_212 
+ bl[210] br[210] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_213 
+ bl[211] br[211] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_214 
+ bl[212] br[212] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_215 
+ bl[213] br[213] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_216 
+ bl[214] br[214] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_217 
+ bl[215] br[215] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_218 
+ bl[216] br[216] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_219 
+ bl[217] br[217] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_220 
+ bl[218] br[218] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_221 
+ bl[219] br[219] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_222 
+ bl[220] br[220] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_223 
+ bl[221] br[221] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_224 
+ bl[222] br[222] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_225 
+ bl[223] br[223] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_226 
+ bl[224] br[224] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_227 
+ bl[225] br[225] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_228 
+ bl[226] br[226] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_229 
+ bl[227] br[227] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_230 
+ bl[228] br[228] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_231 
+ bl[229] br[229] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_232 
+ bl[230] br[230] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_233 
+ bl[231] br[231] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_234 
+ bl[232] br[232] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_235 
+ bl[233] br[233] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_236 
+ bl[234] br[234] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_237 
+ bl[235] br[235] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_238 
+ bl[236] br[236] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_239 
+ bl[237] br[237] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_240 
+ bl[238] br[238] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_241 
+ bl[239] br[239] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_242 
+ bl[240] br[240] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_243 
+ bl[241] br[241] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_244 
+ bl[242] br[242] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_245 
+ bl[243] br[243] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_246 
+ bl[244] br[244] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_247 
+ bl[245] br[245] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_248 
+ bl[246] br[246] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_249 
+ bl[247] br[247] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_250 
+ bl[248] br[248] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_251 
+ bl[249] br[249] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_252 
+ bl[250] br[250] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_253 
+ bl[251] br[251] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_254 
+ bl[252] br[252] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_255 
+ bl[253] br[253] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_256 
+ bl[254] br[254] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_257 
+ bl[255] br[255] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_258 
+ vdd vdd vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_259 
+ vdd vdd vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_0 
+ vdd vdd vss vdd vpb vnb wl[73] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_75_1 
+ rbl rbr vss vdd vpb vnb wl[73] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_75_2 
+ bl[0] br[0] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_3 
+ bl[1] br[1] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_4 
+ bl[2] br[2] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_5 
+ bl[3] br[3] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_6 
+ bl[4] br[4] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_7 
+ bl[5] br[5] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_8 
+ bl[6] br[6] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_9 
+ bl[7] br[7] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_10 
+ bl[8] br[8] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_11 
+ bl[9] br[9] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_12 
+ bl[10] br[10] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_13 
+ bl[11] br[11] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_14 
+ bl[12] br[12] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_15 
+ bl[13] br[13] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_16 
+ bl[14] br[14] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_17 
+ bl[15] br[15] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_18 
+ bl[16] br[16] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_19 
+ bl[17] br[17] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_20 
+ bl[18] br[18] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_21 
+ bl[19] br[19] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_22 
+ bl[20] br[20] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_23 
+ bl[21] br[21] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_24 
+ bl[22] br[22] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_25 
+ bl[23] br[23] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_26 
+ bl[24] br[24] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_27 
+ bl[25] br[25] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_28 
+ bl[26] br[26] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_29 
+ bl[27] br[27] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_30 
+ bl[28] br[28] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_31 
+ bl[29] br[29] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_32 
+ bl[30] br[30] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_33 
+ bl[31] br[31] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_34 
+ bl[32] br[32] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_35 
+ bl[33] br[33] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_36 
+ bl[34] br[34] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_37 
+ bl[35] br[35] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_38 
+ bl[36] br[36] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_39 
+ bl[37] br[37] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_40 
+ bl[38] br[38] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_41 
+ bl[39] br[39] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_42 
+ bl[40] br[40] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_43 
+ bl[41] br[41] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_44 
+ bl[42] br[42] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_45 
+ bl[43] br[43] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_46 
+ bl[44] br[44] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_47 
+ bl[45] br[45] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_48 
+ bl[46] br[46] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_49 
+ bl[47] br[47] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_50 
+ bl[48] br[48] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_51 
+ bl[49] br[49] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_52 
+ bl[50] br[50] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_53 
+ bl[51] br[51] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_54 
+ bl[52] br[52] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_55 
+ bl[53] br[53] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_56 
+ bl[54] br[54] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_57 
+ bl[55] br[55] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_58 
+ bl[56] br[56] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_59 
+ bl[57] br[57] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_60 
+ bl[58] br[58] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_61 
+ bl[59] br[59] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_62 
+ bl[60] br[60] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_63 
+ bl[61] br[61] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_64 
+ bl[62] br[62] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_65 
+ bl[63] br[63] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_66 
+ bl[64] br[64] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_67 
+ bl[65] br[65] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_68 
+ bl[66] br[66] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_69 
+ bl[67] br[67] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_70 
+ bl[68] br[68] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_71 
+ bl[69] br[69] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_72 
+ bl[70] br[70] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_73 
+ bl[71] br[71] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_74 
+ bl[72] br[72] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_75 
+ bl[73] br[73] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_76 
+ bl[74] br[74] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_77 
+ bl[75] br[75] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_78 
+ bl[76] br[76] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_79 
+ bl[77] br[77] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_80 
+ bl[78] br[78] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_81 
+ bl[79] br[79] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_82 
+ bl[80] br[80] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_83 
+ bl[81] br[81] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_84 
+ bl[82] br[82] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_85 
+ bl[83] br[83] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_86 
+ bl[84] br[84] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_87 
+ bl[85] br[85] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_88 
+ bl[86] br[86] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_89 
+ bl[87] br[87] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_90 
+ bl[88] br[88] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_91 
+ bl[89] br[89] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_92 
+ bl[90] br[90] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_93 
+ bl[91] br[91] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_94 
+ bl[92] br[92] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_95 
+ bl[93] br[93] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_96 
+ bl[94] br[94] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_97 
+ bl[95] br[95] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_98 
+ bl[96] br[96] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_99 
+ bl[97] br[97] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_100 
+ bl[98] br[98] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_101 
+ bl[99] br[99] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_102 
+ bl[100] br[100] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_103 
+ bl[101] br[101] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_104 
+ bl[102] br[102] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_105 
+ bl[103] br[103] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_106 
+ bl[104] br[104] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_107 
+ bl[105] br[105] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_108 
+ bl[106] br[106] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_109 
+ bl[107] br[107] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_110 
+ bl[108] br[108] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_111 
+ bl[109] br[109] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_112 
+ bl[110] br[110] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_113 
+ bl[111] br[111] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_114 
+ bl[112] br[112] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_115 
+ bl[113] br[113] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_116 
+ bl[114] br[114] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_117 
+ bl[115] br[115] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_118 
+ bl[116] br[116] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_119 
+ bl[117] br[117] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_120 
+ bl[118] br[118] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_121 
+ bl[119] br[119] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_122 
+ bl[120] br[120] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_123 
+ bl[121] br[121] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_124 
+ bl[122] br[122] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_125 
+ bl[123] br[123] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_126 
+ bl[124] br[124] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_127 
+ bl[125] br[125] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_128 
+ bl[126] br[126] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_129 
+ bl[127] br[127] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_130 
+ bl[128] br[128] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_131 
+ bl[129] br[129] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_132 
+ bl[130] br[130] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_133 
+ bl[131] br[131] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_134 
+ bl[132] br[132] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_135 
+ bl[133] br[133] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_136 
+ bl[134] br[134] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_137 
+ bl[135] br[135] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_138 
+ bl[136] br[136] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_139 
+ bl[137] br[137] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_140 
+ bl[138] br[138] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_141 
+ bl[139] br[139] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_142 
+ bl[140] br[140] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_143 
+ bl[141] br[141] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_144 
+ bl[142] br[142] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_145 
+ bl[143] br[143] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_146 
+ bl[144] br[144] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_147 
+ bl[145] br[145] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_148 
+ bl[146] br[146] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_149 
+ bl[147] br[147] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_150 
+ bl[148] br[148] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_151 
+ bl[149] br[149] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_152 
+ bl[150] br[150] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_153 
+ bl[151] br[151] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_154 
+ bl[152] br[152] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_155 
+ bl[153] br[153] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_156 
+ bl[154] br[154] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_157 
+ bl[155] br[155] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_158 
+ bl[156] br[156] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_159 
+ bl[157] br[157] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_160 
+ bl[158] br[158] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_161 
+ bl[159] br[159] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_162 
+ bl[160] br[160] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_163 
+ bl[161] br[161] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_164 
+ bl[162] br[162] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_165 
+ bl[163] br[163] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_166 
+ bl[164] br[164] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_167 
+ bl[165] br[165] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_168 
+ bl[166] br[166] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_169 
+ bl[167] br[167] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_170 
+ bl[168] br[168] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_171 
+ bl[169] br[169] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_172 
+ bl[170] br[170] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_173 
+ bl[171] br[171] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_174 
+ bl[172] br[172] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_175 
+ bl[173] br[173] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_176 
+ bl[174] br[174] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_177 
+ bl[175] br[175] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_178 
+ bl[176] br[176] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_179 
+ bl[177] br[177] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_180 
+ bl[178] br[178] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_181 
+ bl[179] br[179] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_182 
+ bl[180] br[180] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_183 
+ bl[181] br[181] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_184 
+ bl[182] br[182] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_185 
+ bl[183] br[183] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_186 
+ bl[184] br[184] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_187 
+ bl[185] br[185] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_188 
+ bl[186] br[186] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_189 
+ bl[187] br[187] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_190 
+ bl[188] br[188] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_191 
+ bl[189] br[189] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_192 
+ bl[190] br[190] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_193 
+ bl[191] br[191] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_194 
+ bl[192] br[192] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_195 
+ bl[193] br[193] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_196 
+ bl[194] br[194] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_197 
+ bl[195] br[195] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_198 
+ bl[196] br[196] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_199 
+ bl[197] br[197] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_200 
+ bl[198] br[198] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_201 
+ bl[199] br[199] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_202 
+ bl[200] br[200] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_203 
+ bl[201] br[201] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_204 
+ bl[202] br[202] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_205 
+ bl[203] br[203] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_206 
+ bl[204] br[204] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_207 
+ bl[205] br[205] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_208 
+ bl[206] br[206] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_209 
+ bl[207] br[207] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_210 
+ bl[208] br[208] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_211 
+ bl[209] br[209] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_212 
+ bl[210] br[210] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_213 
+ bl[211] br[211] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_214 
+ bl[212] br[212] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_215 
+ bl[213] br[213] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_216 
+ bl[214] br[214] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_217 
+ bl[215] br[215] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_218 
+ bl[216] br[216] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_219 
+ bl[217] br[217] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_220 
+ bl[218] br[218] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_221 
+ bl[219] br[219] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_222 
+ bl[220] br[220] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_223 
+ bl[221] br[221] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_224 
+ bl[222] br[222] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_225 
+ bl[223] br[223] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_226 
+ bl[224] br[224] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_227 
+ bl[225] br[225] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_228 
+ bl[226] br[226] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_229 
+ bl[227] br[227] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_230 
+ bl[228] br[228] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_231 
+ bl[229] br[229] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_232 
+ bl[230] br[230] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_233 
+ bl[231] br[231] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_234 
+ bl[232] br[232] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_235 
+ bl[233] br[233] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_236 
+ bl[234] br[234] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_237 
+ bl[235] br[235] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_238 
+ bl[236] br[236] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_239 
+ bl[237] br[237] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_240 
+ bl[238] br[238] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_241 
+ bl[239] br[239] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_242 
+ bl[240] br[240] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_243 
+ bl[241] br[241] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_244 
+ bl[242] br[242] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_245 
+ bl[243] br[243] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_246 
+ bl[244] br[244] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_247 
+ bl[245] br[245] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_248 
+ bl[246] br[246] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_249 
+ bl[247] br[247] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_250 
+ bl[248] br[248] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_251 
+ bl[249] br[249] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_252 
+ bl[250] br[250] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_253 
+ bl[251] br[251] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_254 
+ bl[252] br[252] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_255 
+ bl[253] br[253] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_256 
+ bl[254] br[254] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_257 
+ bl[255] br[255] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_258 
+ vdd vdd vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_259 
+ vdd vdd vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_0 
+ vdd vdd vss vdd vpb vnb wl[74] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_76_1 
+ rbl rbr vss vdd vpb vnb wl[74] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_76_2 
+ bl[0] br[0] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_3 
+ bl[1] br[1] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_4 
+ bl[2] br[2] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_5 
+ bl[3] br[3] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_6 
+ bl[4] br[4] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_7 
+ bl[5] br[5] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_8 
+ bl[6] br[6] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_9 
+ bl[7] br[7] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_10 
+ bl[8] br[8] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_11 
+ bl[9] br[9] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_12 
+ bl[10] br[10] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_13 
+ bl[11] br[11] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_14 
+ bl[12] br[12] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_15 
+ bl[13] br[13] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_16 
+ bl[14] br[14] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_17 
+ bl[15] br[15] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_18 
+ bl[16] br[16] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_19 
+ bl[17] br[17] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_20 
+ bl[18] br[18] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_21 
+ bl[19] br[19] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_22 
+ bl[20] br[20] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_23 
+ bl[21] br[21] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_24 
+ bl[22] br[22] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_25 
+ bl[23] br[23] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_26 
+ bl[24] br[24] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_27 
+ bl[25] br[25] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_28 
+ bl[26] br[26] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_29 
+ bl[27] br[27] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_30 
+ bl[28] br[28] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_31 
+ bl[29] br[29] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_32 
+ bl[30] br[30] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_33 
+ bl[31] br[31] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_34 
+ bl[32] br[32] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_35 
+ bl[33] br[33] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_36 
+ bl[34] br[34] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_37 
+ bl[35] br[35] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_38 
+ bl[36] br[36] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_39 
+ bl[37] br[37] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_40 
+ bl[38] br[38] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_41 
+ bl[39] br[39] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_42 
+ bl[40] br[40] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_43 
+ bl[41] br[41] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_44 
+ bl[42] br[42] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_45 
+ bl[43] br[43] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_46 
+ bl[44] br[44] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_47 
+ bl[45] br[45] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_48 
+ bl[46] br[46] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_49 
+ bl[47] br[47] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_50 
+ bl[48] br[48] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_51 
+ bl[49] br[49] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_52 
+ bl[50] br[50] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_53 
+ bl[51] br[51] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_54 
+ bl[52] br[52] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_55 
+ bl[53] br[53] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_56 
+ bl[54] br[54] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_57 
+ bl[55] br[55] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_58 
+ bl[56] br[56] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_59 
+ bl[57] br[57] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_60 
+ bl[58] br[58] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_61 
+ bl[59] br[59] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_62 
+ bl[60] br[60] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_63 
+ bl[61] br[61] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_64 
+ bl[62] br[62] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_65 
+ bl[63] br[63] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_66 
+ bl[64] br[64] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_67 
+ bl[65] br[65] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_68 
+ bl[66] br[66] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_69 
+ bl[67] br[67] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_70 
+ bl[68] br[68] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_71 
+ bl[69] br[69] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_72 
+ bl[70] br[70] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_73 
+ bl[71] br[71] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_74 
+ bl[72] br[72] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_75 
+ bl[73] br[73] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_76 
+ bl[74] br[74] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_77 
+ bl[75] br[75] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_78 
+ bl[76] br[76] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_79 
+ bl[77] br[77] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_80 
+ bl[78] br[78] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_81 
+ bl[79] br[79] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_82 
+ bl[80] br[80] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_83 
+ bl[81] br[81] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_84 
+ bl[82] br[82] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_85 
+ bl[83] br[83] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_86 
+ bl[84] br[84] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_87 
+ bl[85] br[85] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_88 
+ bl[86] br[86] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_89 
+ bl[87] br[87] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_90 
+ bl[88] br[88] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_91 
+ bl[89] br[89] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_92 
+ bl[90] br[90] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_93 
+ bl[91] br[91] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_94 
+ bl[92] br[92] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_95 
+ bl[93] br[93] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_96 
+ bl[94] br[94] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_97 
+ bl[95] br[95] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_98 
+ bl[96] br[96] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_99 
+ bl[97] br[97] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_100 
+ bl[98] br[98] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_101 
+ bl[99] br[99] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_102 
+ bl[100] br[100] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_103 
+ bl[101] br[101] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_104 
+ bl[102] br[102] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_105 
+ bl[103] br[103] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_106 
+ bl[104] br[104] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_107 
+ bl[105] br[105] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_108 
+ bl[106] br[106] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_109 
+ bl[107] br[107] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_110 
+ bl[108] br[108] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_111 
+ bl[109] br[109] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_112 
+ bl[110] br[110] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_113 
+ bl[111] br[111] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_114 
+ bl[112] br[112] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_115 
+ bl[113] br[113] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_116 
+ bl[114] br[114] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_117 
+ bl[115] br[115] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_118 
+ bl[116] br[116] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_119 
+ bl[117] br[117] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_120 
+ bl[118] br[118] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_121 
+ bl[119] br[119] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_122 
+ bl[120] br[120] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_123 
+ bl[121] br[121] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_124 
+ bl[122] br[122] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_125 
+ bl[123] br[123] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_126 
+ bl[124] br[124] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_127 
+ bl[125] br[125] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_128 
+ bl[126] br[126] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_129 
+ bl[127] br[127] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_130 
+ bl[128] br[128] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_131 
+ bl[129] br[129] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_132 
+ bl[130] br[130] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_133 
+ bl[131] br[131] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_134 
+ bl[132] br[132] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_135 
+ bl[133] br[133] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_136 
+ bl[134] br[134] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_137 
+ bl[135] br[135] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_138 
+ bl[136] br[136] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_139 
+ bl[137] br[137] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_140 
+ bl[138] br[138] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_141 
+ bl[139] br[139] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_142 
+ bl[140] br[140] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_143 
+ bl[141] br[141] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_144 
+ bl[142] br[142] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_145 
+ bl[143] br[143] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_146 
+ bl[144] br[144] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_147 
+ bl[145] br[145] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_148 
+ bl[146] br[146] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_149 
+ bl[147] br[147] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_150 
+ bl[148] br[148] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_151 
+ bl[149] br[149] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_152 
+ bl[150] br[150] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_153 
+ bl[151] br[151] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_154 
+ bl[152] br[152] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_155 
+ bl[153] br[153] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_156 
+ bl[154] br[154] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_157 
+ bl[155] br[155] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_158 
+ bl[156] br[156] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_159 
+ bl[157] br[157] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_160 
+ bl[158] br[158] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_161 
+ bl[159] br[159] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_162 
+ bl[160] br[160] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_163 
+ bl[161] br[161] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_164 
+ bl[162] br[162] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_165 
+ bl[163] br[163] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_166 
+ bl[164] br[164] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_167 
+ bl[165] br[165] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_168 
+ bl[166] br[166] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_169 
+ bl[167] br[167] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_170 
+ bl[168] br[168] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_171 
+ bl[169] br[169] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_172 
+ bl[170] br[170] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_173 
+ bl[171] br[171] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_174 
+ bl[172] br[172] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_175 
+ bl[173] br[173] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_176 
+ bl[174] br[174] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_177 
+ bl[175] br[175] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_178 
+ bl[176] br[176] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_179 
+ bl[177] br[177] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_180 
+ bl[178] br[178] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_181 
+ bl[179] br[179] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_182 
+ bl[180] br[180] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_183 
+ bl[181] br[181] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_184 
+ bl[182] br[182] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_185 
+ bl[183] br[183] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_186 
+ bl[184] br[184] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_187 
+ bl[185] br[185] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_188 
+ bl[186] br[186] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_189 
+ bl[187] br[187] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_190 
+ bl[188] br[188] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_191 
+ bl[189] br[189] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_192 
+ bl[190] br[190] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_193 
+ bl[191] br[191] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_194 
+ bl[192] br[192] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_195 
+ bl[193] br[193] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_196 
+ bl[194] br[194] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_197 
+ bl[195] br[195] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_198 
+ bl[196] br[196] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_199 
+ bl[197] br[197] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_200 
+ bl[198] br[198] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_201 
+ bl[199] br[199] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_202 
+ bl[200] br[200] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_203 
+ bl[201] br[201] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_204 
+ bl[202] br[202] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_205 
+ bl[203] br[203] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_206 
+ bl[204] br[204] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_207 
+ bl[205] br[205] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_208 
+ bl[206] br[206] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_209 
+ bl[207] br[207] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_210 
+ bl[208] br[208] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_211 
+ bl[209] br[209] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_212 
+ bl[210] br[210] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_213 
+ bl[211] br[211] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_214 
+ bl[212] br[212] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_215 
+ bl[213] br[213] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_216 
+ bl[214] br[214] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_217 
+ bl[215] br[215] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_218 
+ bl[216] br[216] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_219 
+ bl[217] br[217] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_220 
+ bl[218] br[218] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_221 
+ bl[219] br[219] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_222 
+ bl[220] br[220] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_223 
+ bl[221] br[221] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_224 
+ bl[222] br[222] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_225 
+ bl[223] br[223] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_226 
+ bl[224] br[224] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_227 
+ bl[225] br[225] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_228 
+ bl[226] br[226] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_229 
+ bl[227] br[227] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_230 
+ bl[228] br[228] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_231 
+ bl[229] br[229] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_232 
+ bl[230] br[230] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_233 
+ bl[231] br[231] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_234 
+ bl[232] br[232] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_235 
+ bl[233] br[233] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_236 
+ bl[234] br[234] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_237 
+ bl[235] br[235] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_238 
+ bl[236] br[236] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_239 
+ bl[237] br[237] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_240 
+ bl[238] br[238] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_241 
+ bl[239] br[239] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_242 
+ bl[240] br[240] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_243 
+ bl[241] br[241] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_244 
+ bl[242] br[242] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_245 
+ bl[243] br[243] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_246 
+ bl[244] br[244] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_247 
+ bl[245] br[245] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_248 
+ bl[246] br[246] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_249 
+ bl[247] br[247] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_250 
+ bl[248] br[248] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_251 
+ bl[249] br[249] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_252 
+ bl[250] br[250] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_253 
+ bl[251] br[251] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_254 
+ bl[252] br[252] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_255 
+ bl[253] br[253] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_256 
+ bl[254] br[254] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_257 
+ bl[255] br[255] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_258 
+ vdd vdd vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_259 
+ vdd vdd vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_0 
+ vdd vdd vss vdd vpb vnb wl[75] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_77_1 
+ rbl rbr vss vdd vpb vnb wl[75] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_77_2 
+ bl[0] br[0] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_3 
+ bl[1] br[1] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_4 
+ bl[2] br[2] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_5 
+ bl[3] br[3] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_6 
+ bl[4] br[4] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_7 
+ bl[5] br[5] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_8 
+ bl[6] br[6] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_9 
+ bl[7] br[7] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_10 
+ bl[8] br[8] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_11 
+ bl[9] br[9] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_12 
+ bl[10] br[10] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_13 
+ bl[11] br[11] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_14 
+ bl[12] br[12] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_15 
+ bl[13] br[13] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_16 
+ bl[14] br[14] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_17 
+ bl[15] br[15] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_18 
+ bl[16] br[16] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_19 
+ bl[17] br[17] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_20 
+ bl[18] br[18] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_21 
+ bl[19] br[19] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_22 
+ bl[20] br[20] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_23 
+ bl[21] br[21] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_24 
+ bl[22] br[22] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_25 
+ bl[23] br[23] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_26 
+ bl[24] br[24] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_27 
+ bl[25] br[25] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_28 
+ bl[26] br[26] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_29 
+ bl[27] br[27] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_30 
+ bl[28] br[28] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_31 
+ bl[29] br[29] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_32 
+ bl[30] br[30] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_33 
+ bl[31] br[31] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_34 
+ bl[32] br[32] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_35 
+ bl[33] br[33] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_36 
+ bl[34] br[34] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_37 
+ bl[35] br[35] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_38 
+ bl[36] br[36] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_39 
+ bl[37] br[37] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_40 
+ bl[38] br[38] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_41 
+ bl[39] br[39] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_42 
+ bl[40] br[40] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_43 
+ bl[41] br[41] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_44 
+ bl[42] br[42] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_45 
+ bl[43] br[43] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_46 
+ bl[44] br[44] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_47 
+ bl[45] br[45] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_48 
+ bl[46] br[46] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_49 
+ bl[47] br[47] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_50 
+ bl[48] br[48] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_51 
+ bl[49] br[49] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_52 
+ bl[50] br[50] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_53 
+ bl[51] br[51] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_54 
+ bl[52] br[52] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_55 
+ bl[53] br[53] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_56 
+ bl[54] br[54] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_57 
+ bl[55] br[55] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_58 
+ bl[56] br[56] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_59 
+ bl[57] br[57] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_60 
+ bl[58] br[58] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_61 
+ bl[59] br[59] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_62 
+ bl[60] br[60] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_63 
+ bl[61] br[61] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_64 
+ bl[62] br[62] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_65 
+ bl[63] br[63] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_66 
+ bl[64] br[64] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_67 
+ bl[65] br[65] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_68 
+ bl[66] br[66] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_69 
+ bl[67] br[67] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_70 
+ bl[68] br[68] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_71 
+ bl[69] br[69] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_72 
+ bl[70] br[70] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_73 
+ bl[71] br[71] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_74 
+ bl[72] br[72] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_75 
+ bl[73] br[73] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_76 
+ bl[74] br[74] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_77 
+ bl[75] br[75] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_78 
+ bl[76] br[76] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_79 
+ bl[77] br[77] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_80 
+ bl[78] br[78] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_81 
+ bl[79] br[79] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_82 
+ bl[80] br[80] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_83 
+ bl[81] br[81] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_84 
+ bl[82] br[82] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_85 
+ bl[83] br[83] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_86 
+ bl[84] br[84] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_87 
+ bl[85] br[85] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_88 
+ bl[86] br[86] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_89 
+ bl[87] br[87] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_90 
+ bl[88] br[88] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_91 
+ bl[89] br[89] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_92 
+ bl[90] br[90] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_93 
+ bl[91] br[91] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_94 
+ bl[92] br[92] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_95 
+ bl[93] br[93] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_96 
+ bl[94] br[94] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_97 
+ bl[95] br[95] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_98 
+ bl[96] br[96] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_99 
+ bl[97] br[97] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_100 
+ bl[98] br[98] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_101 
+ bl[99] br[99] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_102 
+ bl[100] br[100] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_103 
+ bl[101] br[101] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_104 
+ bl[102] br[102] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_105 
+ bl[103] br[103] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_106 
+ bl[104] br[104] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_107 
+ bl[105] br[105] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_108 
+ bl[106] br[106] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_109 
+ bl[107] br[107] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_110 
+ bl[108] br[108] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_111 
+ bl[109] br[109] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_112 
+ bl[110] br[110] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_113 
+ bl[111] br[111] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_114 
+ bl[112] br[112] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_115 
+ bl[113] br[113] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_116 
+ bl[114] br[114] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_117 
+ bl[115] br[115] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_118 
+ bl[116] br[116] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_119 
+ bl[117] br[117] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_120 
+ bl[118] br[118] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_121 
+ bl[119] br[119] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_122 
+ bl[120] br[120] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_123 
+ bl[121] br[121] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_124 
+ bl[122] br[122] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_125 
+ bl[123] br[123] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_126 
+ bl[124] br[124] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_127 
+ bl[125] br[125] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_128 
+ bl[126] br[126] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_129 
+ bl[127] br[127] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_130 
+ bl[128] br[128] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_131 
+ bl[129] br[129] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_132 
+ bl[130] br[130] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_133 
+ bl[131] br[131] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_134 
+ bl[132] br[132] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_135 
+ bl[133] br[133] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_136 
+ bl[134] br[134] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_137 
+ bl[135] br[135] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_138 
+ bl[136] br[136] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_139 
+ bl[137] br[137] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_140 
+ bl[138] br[138] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_141 
+ bl[139] br[139] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_142 
+ bl[140] br[140] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_143 
+ bl[141] br[141] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_144 
+ bl[142] br[142] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_145 
+ bl[143] br[143] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_146 
+ bl[144] br[144] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_147 
+ bl[145] br[145] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_148 
+ bl[146] br[146] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_149 
+ bl[147] br[147] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_150 
+ bl[148] br[148] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_151 
+ bl[149] br[149] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_152 
+ bl[150] br[150] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_153 
+ bl[151] br[151] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_154 
+ bl[152] br[152] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_155 
+ bl[153] br[153] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_156 
+ bl[154] br[154] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_157 
+ bl[155] br[155] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_158 
+ bl[156] br[156] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_159 
+ bl[157] br[157] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_160 
+ bl[158] br[158] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_161 
+ bl[159] br[159] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_162 
+ bl[160] br[160] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_163 
+ bl[161] br[161] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_164 
+ bl[162] br[162] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_165 
+ bl[163] br[163] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_166 
+ bl[164] br[164] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_167 
+ bl[165] br[165] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_168 
+ bl[166] br[166] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_169 
+ bl[167] br[167] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_170 
+ bl[168] br[168] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_171 
+ bl[169] br[169] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_172 
+ bl[170] br[170] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_173 
+ bl[171] br[171] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_174 
+ bl[172] br[172] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_175 
+ bl[173] br[173] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_176 
+ bl[174] br[174] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_177 
+ bl[175] br[175] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_178 
+ bl[176] br[176] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_179 
+ bl[177] br[177] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_180 
+ bl[178] br[178] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_181 
+ bl[179] br[179] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_182 
+ bl[180] br[180] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_183 
+ bl[181] br[181] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_184 
+ bl[182] br[182] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_185 
+ bl[183] br[183] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_186 
+ bl[184] br[184] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_187 
+ bl[185] br[185] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_188 
+ bl[186] br[186] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_189 
+ bl[187] br[187] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_190 
+ bl[188] br[188] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_191 
+ bl[189] br[189] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_192 
+ bl[190] br[190] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_193 
+ bl[191] br[191] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_194 
+ bl[192] br[192] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_195 
+ bl[193] br[193] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_196 
+ bl[194] br[194] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_197 
+ bl[195] br[195] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_198 
+ bl[196] br[196] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_199 
+ bl[197] br[197] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_200 
+ bl[198] br[198] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_201 
+ bl[199] br[199] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_202 
+ bl[200] br[200] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_203 
+ bl[201] br[201] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_204 
+ bl[202] br[202] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_205 
+ bl[203] br[203] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_206 
+ bl[204] br[204] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_207 
+ bl[205] br[205] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_208 
+ bl[206] br[206] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_209 
+ bl[207] br[207] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_210 
+ bl[208] br[208] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_211 
+ bl[209] br[209] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_212 
+ bl[210] br[210] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_213 
+ bl[211] br[211] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_214 
+ bl[212] br[212] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_215 
+ bl[213] br[213] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_216 
+ bl[214] br[214] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_217 
+ bl[215] br[215] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_218 
+ bl[216] br[216] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_219 
+ bl[217] br[217] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_220 
+ bl[218] br[218] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_221 
+ bl[219] br[219] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_222 
+ bl[220] br[220] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_223 
+ bl[221] br[221] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_224 
+ bl[222] br[222] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_225 
+ bl[223] br[223] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_226 
+ bl[224] br[224] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_227 
+ bl[225] br[225] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_228 
+ bl[226] br[226] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_229 
+ bl[227] br[227] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_230 
+ bl[228] br[228] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_231 
+ bl[229] br[229] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_232 
+ bl[230] br[230] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_233 
+ bl[231] br[231] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_234 
+ bl[232] br[232] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_235 
+ bl[233] br[233] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_236 
+ bl[234] br[234] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_237 
+ bl[235] br[235] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_238 
+ bl[236] br[236] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_239 
+ bl[237] br[237] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_240 
+ bl[238] br[238] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_241 
+ bl[239] br[239] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_242 
+ bl[240] br[240] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_243 
+ bl[241] br[241] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_244 
+ bl[242] br[242] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_245 
+ bl[243] br[243] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_246 
+ bl[244] br[244] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_247 
+ bl[245] br[245] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_248 
+ bl[246] br[246] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_249 
+ bl[247] br[247] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_250 
+ bl[248] br[248] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_251 
+ bl[249] br[249] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_252 
+ bl[250] br[250] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_253 
+ bl[251] br[251] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_254 
+ bl[252] br[252] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_255 
+ bl[253] br[253] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_256 
+ bl[254] br[254] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_257 
+ bl[255] br[255] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_258 
+ vdd vdd vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_259 
+ vdd vdd vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_0 
+ vdd vdd vss vdd vpb vnb wl[76] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_78_1 
+ rbl rbr vss vdd vpb vnb wl[76] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_78_2 
+ bl[0] br[0] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_3 
+ bl[1] br[1] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_4 
+ bl[2] br[2] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_5 
+ bl[3] br[3] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_6 
+ bl[4] br[4] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_7 
+ bl[5] br[5] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_8 
+ bl[6] br[6] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_9 
+ bl[7] br[7] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_10 
+ bl[8] br[8] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_11 
+ bl[9] br[9] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_12 
+ bl[10] br[10] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_13 
+ bl[11] br[11] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_14 
+ bl[12] br[12] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_15 
+ bl[13] br[13] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_16 
+ bl[14] br[14] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_17 
+ bl[15] br[15] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_18 
+ bl[16] br[16] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_19 
+ bl[17] br[17] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_20 
+ bl[18] br[18] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_21 
+ bl[19] br[19] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_22 
+ bl[20] br[20] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_23 
+ bl[21] br[21] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_24 
+ bl[22] br[22] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_25 
+ bl[23] br[23] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_26 
+ bl[24] br[24] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_27 
+ bl[25] br[25] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_28 
+ bl[26] br[26] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_29 
+ bl[27] br[27] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_30 
+ bl[28] br[28] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_31 
+ bl[29] br[29] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_32 
+ bl[30] br[30] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_33 
+ bl[31] br[31] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_34 
+ bl[32] br[32] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_35 
+ bl[33] br[33] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_36 
+ bl[34] br[34] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_37 
+ bl[35] br[35] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_38 
+ bl[36] br[36] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_39 
+ bl[37] br[37] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_40 
+ bl[38] br[38] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_41 
+ bl[39] br[39] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_42 
+ bl[40] br[40] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_43 
+ bl[41] br[41] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_44 
+ bl[42] br[42] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_45 
+ bl[43] br[43] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_46 
+ bl[44] br[44] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_47 
+ bl[45] br[45] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_48 
+ bl[46] br[46] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_49 
+ bl[47] br[47] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_50 
+ bl[48] br[48] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_51 
+ bl[49] br[49] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_52 
+ bl[50] br[50] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_53 
+ bl[51] br[51] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_54 
+ bl[52] br[52] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_55 
+ bl[53] br[53] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_56 
+ bl[54] br[54] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_57 
+ bl[55] br[55] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_58 
+ bl[56] br[56] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_59 
+ bl[57] br[57] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_60 
+ bl[58] br[58] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_61 
+ bl[59] br[59] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_62 
+ bl[60] br[60] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_63 
+ bl[61] br[61] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_64 
+ bl[62] br[62] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_65 
+ bl[63] br[63] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_66 
+ bl[64] br[64] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_67 
+ bl[65] br[65] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_68 
+ bl[66] br[66] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_69 
+ bl[67] br[67] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_70 
+ bl[68] br[68] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_71 
+ bl[69] br[69] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_72 
+ bl[70] br[70] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_73 
+ bl[71] br[71] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_74 
+ bl[72] br[72] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_75 
+ bl[73] br[73] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_76 
+ bl[74] br[74] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_77 
+ bl[75] br[75] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_78 
+ bl[76] br[76] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_79 
+ bl[77] br[77] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_80 
+ bl[78] br[78] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_81 
+ bl[79] br[79] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_82 
+ bl[80] br[80] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_83 
+ bl[81] br[81] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_84 
+ bl[82] br[82] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_85 
+ bl[83] br[83] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_86 
+ bl[84] br[84] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_87 
+ bl[85] br[85] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_88 
+ bl[86] br[86] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_89 
+ bl[87] br[87] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_90 
+ bl[88] br[88] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_91 
+ bl[89] br[89] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_92 
+ bl[90] br[90] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_93 
+ bl[91] br[91] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_94 
+ bl[92] br[92] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_95 
+ bl[93] br[93] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_96 
+ bl[94] br[94] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_97 
+ bl[95] br[95] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_98 
+ bl[96] br[96] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_99 
+ bl[97] br[97] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_100 
+ bl[98] br[98] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_101 
+ bl[99] br[99] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_102 
+ bl[100] br[100] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_103 
+ bl[101] br[101] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_104 
+ bl[102] br[102] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_105 
+ bl[103] br[103] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_106 
+ bl[104] br[104] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_107 
+ bl[105] br[105] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_108 
+ bl[106] br[106] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_109 
+ bl[107] br[107] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_110 
+ bl[108] br[108] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_111 
+ bl[109] br[109] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_112 
+ bl[110] br[110] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_113 
+ bl[111] br[111] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_114 
+ bl[112] br[112] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_115 
+ bl[113] br[113] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_116 
+ bl[114] br[114] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_117 
+ bl[115] br[115] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_118 
+ bl[116] br[116] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_119 
+ bl[117] br[117] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_120 
+ bl[118] br[118] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_121 
+ bl[119] br[119] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_122 
+ bl[120] br[120] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_123 
+ bl[121] br[121] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_124 
+ bl[122] br[122] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_125 
+ bl[123] br[123] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_126 
+ bl[124] br[124] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_127 
+ bl[125] br[125] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_128 
+ bl[126] br[126] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_129 
+ bl[127] br[127] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_130 
+ bl[128] br[128] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_131 
+ bl[129] br[129] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_132 
+ bl[130] br[130] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_133 
+ bl[131] br[131] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_134 
+ bl[132] br[132] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_135 
+ bl[133] br[133] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_136 
+ bl[134] br[134] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_137 
+ bl[135] br[135] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_138 
+ bl[136] br[136] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_139 
+ bl[137] br[137] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_140 
+ bl[138] br[138] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_141 
+ bl[139] br[139] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_142 
+ bl[140] br[140] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_143 
+ bl[141] br[141] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_144 
+ bl[142] br[142] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_145 
+ bl[143] br[143] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_146 
+ bl[144] br[144] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_147 
+ bl[145] br[145] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_148 
+ bl[146] br[146] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_149 
+ bl[147] br[147] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_150 
+ bl[148] br[148] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_151 
+ bl[149] br[149] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_152 
+ bl[150] br[150] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_153 
+ bl[151] br[151] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_154 
+ bl[152] br[152] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_155 
+ bl[153] br[153] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_156 
+ bl[154] br[154] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_157 
+ bl[155] br[155] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_158 
+ bl[156] br[156] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_159 
+ bl[157] br[157] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_160 
+ bl[158] br[158] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_161 
+ bl[159] br[159] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_162 
+ bl[160] br[160] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_163 
+ bl[161] br[161] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_164 
+ bl[162] br[162] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_165 
+ bl[163] br[163] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_166 
+ bl[164] br[164] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_167 
+ bl[165] br[165] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_168 
+ bl[166] br[166] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_169 
+ bl[167] br[167] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_170 
+ bl[168] br[168] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_171 
+ bl[169] br[169] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_172 
+ bl[170] br[170] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_173 
+ bl[171] br[171] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_174 
+ bl[172] br[172] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_175 
+ bl[173] br[173] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_176 
+ bl[174] br[174] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_177 
+ bl[175] br[175] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_178 
+ bl[176] br[176] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_179 
+ bl[177] br[177] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_180 
+ bl[178] br[178] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_181 
+ bl[179] br[179] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_182 
+ bl[180] br[180] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_183 
+ bl[181] br[181] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_184 
+ bl[182] br[182] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_185 
+ bl[183] br[183] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_186 
+ bl[184] br[184] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_187 
+ bl[185] br[185] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_188 
+ bl[186] br[186] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_189 
+ bl[187] br[187] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_190 
+ bl[188] br[188] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_191 
+ bl[189] br[189] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_192 
+ bl[190] br[190] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_193 
+ bl[191] br[191] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_194 
+ bl[192] br[192] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_195 
+ bl[193] br[193] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_196 
+ bl[194] br[194] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_197 
+ bl[195] br[195] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_198 
+ bl[196] br[196] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_199 
+ bl[197] br[197] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_200 
+ bl[198] br[198] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_201 
+ bl[199] br[199] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_202 
+ bl[200] br[200] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_203 
+ bl[201] br[201] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_204 
+ bl[202] br[202] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_205 
+ bl[203] br[203] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_206 
+ bl[204] br[204] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_207 
+ bl[205] br[205] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_208 
+ bl[206] br[206] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_209 
+ bl[207] br[207] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_210 
+ bl[208] br[208] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_211 
+ bl[209] br[209] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_212 
+ bl[210] br[210] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_213 
+ bl[211] br[211] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_214 
+ bl[212] br[212] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_215 
+ bl[213] br[213] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_216 
+ bl[214] br[214] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_217 
+ bl[215] br[215] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_218 
+ bl[216] br[216] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_219 
+ bl[217] br[217] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_220 
+ bl[218] br[218] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_221 
+ bl[219] br[219] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_222 
+ bl[220] br[220] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_223 
+ bl[221] br[221] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_224 
+ bl[222] br[222] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_225 
+ bl[223] br[223] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_226 
+ bl[224] br[224] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_227 
+ bl[225] br[225] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_228 
+ bl[226] br[226] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_229 
+ bl[227] br[227] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_230 
+ bl[228] br[228] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_231 
+ bl[229] br[229] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_232 
+ bl[230] br[230] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_233 
+ bl[231] br[231] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_234 
+ bl[232] br[232] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_235 
+ bl[233] br[233] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_236 
+ bl[234] br[234] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_237 
+ bl[235] br[235] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_238 
+ bl[236] br[236] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_239 
+ bl[237] br[237] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_240 
+ bl[238] br[238] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_241 
+ bl[239] br[239] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_242 
+ bl[240] br[240] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_243 
+ bl[241] br[241] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_244 
+ bl[242] br[242] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_245 
+ bl[243] br[243] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_246 
+ bl[244] br[244] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_247 
+ bl[245] br[245] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_248 
+ bl[246] br[246] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_249 
+ bl[247] br[247] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_250 
+ bl[248] br[248] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_251 
+ bl[249] br[249] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_252 
+ bl[250] br[250] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_253 
+ bl[251] br[251] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_254 
+ bl[252] br[252] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_255 
+ bl[253] br[253] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_256 
+ bl[254] br[254] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_257 
+ bl[255] br[255] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_258 
+ vdd vdd vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_259 
+ vdd vdd vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_0 
+ vdd vdd vss vdd vpb vnb wl[77] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_79_1 
+ rbl rbr vss vdd vpb vnb wl[77] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_79_2 
+ bl[0] br[0] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_3 
+ bl[1] br[1] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_4 
+ bl[2] br[2] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_5 
+ bl[3] br[3] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_6 
+ bl[4] br[4] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_7 
+ bl[5] br[5] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_8 
+ bl[6] br[6] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_9 
+ bl[7] br[7] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_10 
+ bl[8] br[8] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_11 
+ bl[9] br[9] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_12 
+ bl[10] br[10] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_13 
+ bl[11] br[11] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_14 
+ bl[12] br[12] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_15 
+ bl[13] br[13] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_16 
+ bl[14] br[14] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_17 
+ bl[15] br[15] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_18 
+ bl[16] br[16] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_19 
+ bl[17] br[17] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_20 
+ bl[18] br[18] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_21 
+ bl[19] br[19] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_22 
+ bl[20] br[20] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_23 
+ bl[21] br[21] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_24 
+ bl[22] br[22] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_25 
+ bl[23] br[23] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_26 
+ bl[24] br[24] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_27 
+ bl[25] br[25] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_28 
+ bl[26] br[26] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_29 
+ bl[27] br[27] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_30 
+ bl[28] br[28] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_31 
+ bl[29] br[29] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_32 
+ bl[30] br[30] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_33 
+ bl[31] br[31] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_34 
+ bl[32] br[32] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_35 
+ bl[33] br[33] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_36 
+ bl[34] br[34] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_37 
+ bl[35] br[35] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_38 
+ bl[36] br[36] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_39 
+ bl[37] br[37] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_40 
+ bl[38] br[38] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_41 
+ bl[39] br[39] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_42 
+ bl[40] br[40] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_43 
+ bl[41] br[41] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_44 
+ bl[42] br[42] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_45 
+ bl[43] br[43] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_46 
+ bl[44] br[44] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_47 
+ bl[45] br[45] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_48 
+ bl[46] br[46] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_49 
+ bl[47] br[47] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_50 
+ bl[48] br[48] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_51 
+ bl[49] br[49] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_52 
+ bl[50] br[50] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_53 
+ bl[51] br[51] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_54 
+ bl[52] br[52] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_55 
+ bl[53] br[53] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_56 
+ bl[54] br[54] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_57 
+ bl[55] br[55] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_58 
+ bl[56] br[56] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_59 
+ bl[57] br[57] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_60 
+ bl[58] br[58] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_61 
+ bl[59] br[59] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_62 
+ bl[60] br[60] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_63 
+ bl[61] br[61] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_64 
+ bl[62] br[62] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_65 
+ bl[63] br[63] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_66 
+ bl[64] br[64] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_67 
+ bl[65] br[65] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_68 
+ bl[66] br[66] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_69 
+ bl[67] br[67] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_70 
+ bl[68] br[68] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_71 
+ bl[69] br[69] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_72 
+ bl[70] br[70] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_73 
+ bl[71] br[71] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_74 
+ bl[72] br[72] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_75 
+ bl[73] br[73] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_76 
+ bl[74] br[74] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_77 
+ bl[75] br[75] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_78 
+ bl[76] br[76] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_79 
+ bl[77] br[77] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_80 
+ bl[78] br[78] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_81 
+ bl[79] br[79] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_82 
+ bl[80] br[80] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_83 
+ bl[81] br[81] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_84 
+ bl[82] br[82] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_85 
+ bl[83] br[83] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_86 
+ bl[84] br[84] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_87 
+ bl[85] br[85] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_88 
+ bl[86] br[86] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_89 
+ bl[87] br[87] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_90 
+ bl[88] br[88] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_91 
+ bl[89] br[89] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_92 
+ bl[90] br[90] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_93 
+ bl[91] br[91] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_94 
+ bl[92] br[92] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_95 
+ bl[93] br[93] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_96 
+ bl[94] br[94] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_97 
+ bl[95] br[95] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_98 
+ bl[96] br[96] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_99 
+ bl[97] br[97] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_100 
+ bl[98] br[98] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_101 
+ bl[99] br[99] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_102 
+ bl[100] br[100] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_103 
+ bl[101] br[101] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_104 
+ bl[102] br[102] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_105 
+ bl[103] br[103] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_106 
+ bl[104] br[104] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_107 
+ bl[105] br[105] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_108 
+ bl[106] br[106] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_109 
+ bl[107] br[107] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_110 
+ bl[108] br[108] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_111 
+ bl[109] br[109] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_112 
+ bl[110] br[110] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_113 
+ bl[111] br[111] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_114 
+ bl[112] br[112] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_115 
+ bl[113] br[113] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_116 
+ bl[114] br[114] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_117 
+ bl[115] br[115] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_118 
+ bl[116] br[116] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_119 
+ bl[117] br[117] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_120 
+ bl[118] br[118] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_121 
+ bl[119] br[119] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_122 
+ bl[120] br[120] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_123 
+ bl[121] br[121] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_124 
+ bl[122] br[122] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_125 
+ bl[123] br[123] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_126 
+ bl[124] br[124] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_127 
+ bl[125] br[125] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_128 
+ bl[126] br[126] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_129 
+ bl[127] br[127] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_130 
+ bl[128] br[128] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_131 
+ bl[129] br[129] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_132 
+ bl[130] br[130] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_133 
+ bl[131] br[131] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_134 
+ bl[132] br[132] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_135 
+ bl[133] br[133] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_136 
+ bl[134] br[134] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_137 
+ bl[135] br[135] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_138 
+ bl[136] br[136] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_139 
+ bl[137] br[137] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_140 
+ bl[138] br[138] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_141 
+ bl[139] br[139] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_142 
+ bl[140] br[140] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_143 
+ bl[141] br[141] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_144 
+ bl[142] br[142] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_145 
+ bl[143] br[143] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_146 
+ bl[144] br[144] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_147 
+ bl[145] br[145] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_148 
+ bl[146] br[146] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_149 
+ bl[147] br[147] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_150 
+ bl[148] br[148] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_151 
+ bl[149] br[149] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_152 
+ bl[150] br[150] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_153 
+ bl[151] br[151] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_154 
+ bl[152] br[152] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_155 
+ bl[153] br[153] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_156 
+ bl[154] br[154] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_157 
+ bl[155] br[155] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_158 
+ bl[156] br[156] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_159 
+ bl[157] br[157] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_160 
+ bl[158] br[158] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_161 
+ bl[159] br[159] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_162 
+ bl[160] br[160] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_163 
+ bl[161] br[161] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_164 
+ bl[162] br[162] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_165 
+ bl[163] br[163] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_166 
+ bl[164] br[164] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_167 
+ bl[165] br[165] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_168 
+ bl[166] br[166] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_169 
+ bl[167] br[167] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_170 
+ bl[168] br[168] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_171 
+ bl[169] br[169] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_172 
+ bl[170] br[170] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_173 
+ bl[171] br[171] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_174 
+ bl[172] br[172] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_175 
+ bl[173] br[173] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_176 
+ bl[174] br[174] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_177 
+ bl[175] br[175] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_178 
+ bl[176] br[176] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_179 
+ bl[177] br[177] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_180 
+ bl[178] br[178] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_181 
+ bl[179] br[179] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_182 
+ bl[180] br[180] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_183 
+ bl[181] br[181] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_184 
+ bl[182] br[182] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_185 
+ bl[183] br[183] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_186 
+ bl[184] br[184] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_187 
+ bl[185] br[185] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_188 
+ bl[186] br[186] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_189 
+ bl[187] br[187] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_190 
+ bl[188] br[188] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_191 
+ bl[189] br[189] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_192 
+ bl[190] br[190] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_193 
+ bl[191] br[191] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_194 
+ bl[192] br[192] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_195 
+ bl[193] br[193] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_196 
+ bl[194] br[194] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_197 
+ bl[195] br[195] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_198 
+ bl[196] br[196] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_199 
+ bl[197] br[197] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_200 
+ bl[198] br[198] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_201 
+ bl[199] br[199] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_202 
+ bl[200] br[200] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_203 
+ bl[201] br[201] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_204 
+ bl[202] br[202] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_205 
+ bl[203] br[203] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_206 
+ bl[204] br[204] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_207 
+ bl[205] br[205] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_208 
+ bl[206] br[206] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_209 
+ bl[207] br[207] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_210 
+ bl[208] br[208] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_211 
+ bl[209] br[209] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_212 
+ bl[210] br[210] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_213 
+ bl[211] br[211] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_214 
+ bl[212] br[212] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_215 
+ bl[213] br[213] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_216 
+ bl[214] br[214] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_217 
+ bl[215] br[215] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_218 
+ bl[216] br[216] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_219 
+ bl[217] br[217] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_220 
+ bl[218] br[218] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_221 
+ bl[219] br[219] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_222 
+ bl[220] br[220] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_223 
+ bl[221] br[221] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_224 
+ bl[222] br[222] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_225 
+ bl[223] br[223] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_226 
+ bl[224] br[224] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_227 
+ bl[225] br[225] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_228 
+ bl[226] br[226] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_229 
+ bl[227] br[227] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_230 
+ bl[228] br[228] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_231 
+ bl[229] br[229] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_232 
+ bl[230] br[230] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_233 
+ bl[231] br[231] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_234 
+ bl[232] br[232] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_235 
+ bl[233] br[233] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_236 
+ bl[234] br[234] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_237 
+ bl[235] br[235] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_238 
+ bl[236] br[236] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_239 
+ bl[237] br[237] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_240 
+ bl[238] br[238] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_241 
+ bl[239] br[239] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_242 
+ bl[240] br[240] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_243 
+ bl[241] br[241] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_244 
+ bl[242] br[242] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_245 
+ bl[243] br[243] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_246 
+ bl[244] br[244] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_247 
+ bl[245] br[245] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_248 
+ bl[246] br[246] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_249 
+ bl[247] br[247] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_250 
+ bl[248] br[248] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_251 
+ bl[249] br[249] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_252 
+ bl[250] br[250] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_253 
+ bl[251] br[251] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_254 
+ bl[252] br[252] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_255 
+ bl[253] br[253] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_256 
+ bl[254] br[254] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_257 
+ bl[255] br[255] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_258 
+ vdd vdd vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_259 
+ vdd vdd vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_0 
+ vdd vdd vss vdd vpb vnb wl[78] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_80_1 
+ rbl rbr vss vdd vpb vnb wl[78] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_80_2 
+ bl[0] br[0] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_3 
+ bl[1] br[1] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_4 
+ bl[2] br[2] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_5 
+ bl[3] br[3] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_6 
+ bl[4] br[4] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_7 
+ bl[5] br[5] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_8 
+ bl[6] br[6] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_9 
+ bl[7] br[7] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_10 
+ bl[8] br[8] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_11 
+ bl[9] br[9] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_12 
+ bl[10] br[10] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_13 
+ bl[11] br[11] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_14 
+ bl[12] br[12] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_15 
+ bl[13] br[13] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_16 
+ bl[14] br[14] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_17 
+ bl[15] br[15] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_18 
+ bl[16] br[16] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_19 
+ bl[17] br[17] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_20 
+ bl[18] br[18] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_21 
+ bl[19] br[19] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_22 
+ bl[20] br[20] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_23 
+ bl[21] br[21] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_24 
+ bl[22] br[22] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_25 
+ bl[23] br[23] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_26 
+ bl[24] br[24] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_27 
+ bl[25] br[25] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_28 
+ bl[26] br[26] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_29 
+ bl[27] br[27] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_30 
+ bl[28] br[28] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_31 
+ bl[29] br[29] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_32 
+ bl[30] br[30] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_33 
+ bl[31] br[31] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_34 
+ bl[32] br[32] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_35 
+ bl[33] br[33] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_36 
+ bl[34] br[34] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_37 
+ bl[35] br[35] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_38 
+ bl[36] br[36] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_39 
+ bl[37] br[37] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_40 
+ bl[38] br[38] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_41 
+ bl[39] br[39] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_42 
+ bl[40] br[40] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_43 
+ bl[41] br[41] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_44 
+ bl[42] br[42] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_45 
+ bl[43] br[43] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_46 
+ bl[44] br[44] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_47 
+ bl[45] br[45] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_48 
+ bl[46] br[46] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_49 
+ bl[47] br[47] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_50 
+ bl[48] br[48] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_51 
+ bl[49] br[49] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_52 
+ bl[50] br[50] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_53 
+ bl[51] br[51] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_54 
+ bl[52] br[52] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_55 
+ bl[53] br[53] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_56 
+ bl[54] br[54] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_57 
+ bl[55] br[55] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_58 
+ bl[56] br[56] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_59 
+ bl[57] br[57] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_60 
+ bl[58] br[58] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_61 
+ bl[59] br[59] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_62 
+ bl[60] br[60] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_63 
+ bl[61] br[61] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_64 
+ bl[62] br[62] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_65 
+ bl[63] br[63] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_66 
+ bl[64] br[64] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_67 
+ bl[65] br[65] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_68 
+ bl[66] br[66] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_69 
+ bl[67] br[67] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_70 
+ bl[68] br[68] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_71 
+ bl[69] br[69] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_72 
+ bl[70] br[70] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_73 
+ bl[71] br[71] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_74 
+ bl[72] br[72] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_75 
+ bl[73] br[73] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_76 
+ bl[74] br[74] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_77 
+ bl[75] br[75] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_78 
+ bl[76] br[76] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_79 
+ bl[77] br[77] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_80 
+ bl[78] br[78] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_81 
+ bl[79] br[79] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_82 
+ bl[80] br[80] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_83 
+ bl[81] br[81] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_84 
+ bl[82] br[82] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_85 
+ bl[83] br[83] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_86 
+ bl[84] br[84] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_87 
+ bl[85] br[85] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_88 
+ bl[86] br[86] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_89 
+ bl[87] br[87] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_90 
+ bl[88] br[88] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_91 
+ bl[89] br[89] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_92 
+ bl[90] br[90] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_93 
+ bl[91] br[91] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_94 
+ bl[92] br[92] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_95 
+ bl[93] br[93] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_96 
+ bl[94] br[94] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_97 
+ bl[95] br[95] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_98 
+ bl[96] br[96] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_99 
+ bl[97] br[97] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_100 
+ bl[98] br[98] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_101 
+ bl[99] br[99] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_102 
+ bl[100] br[100] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_103 
+ bl[101] br[101] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_104 
+ bl[102] br[102] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_105 
+ bl[103] br[103] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_106 
+ bl[104] br[104] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_107 
+ bl[105] br[105] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_108 
+ bl[106] br[106] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_109 
+ bl[107] br[107] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_110 
+ bl[108] br[108] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_111 
+ bl[109] br[109] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_112 
+ bl[110] br[110] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_113 
+ bl[111] br[111] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_114 
+ bl[112] br[112] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_115 
+ bl[113] br[113] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_116 
+ bl[114] br[114] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_117 
+ bl[115] br[115] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_118 
+ bl[116] br[116] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_119 
+ bl[117] br[117] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_120 
+ bl[118] br[118] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_121 
+ bl[119] br[119] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_122 
+ bl[120] br[120] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_123 
+ bl[121] br[121] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_124 
+ bl[122] br[122] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_125 
+ bl[123] br[123] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_126 
+ bl[124] br[124] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_127 
+ bl[125] br[125] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_128 
+ bl[126] br[126] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_129 
+ bl[127] br[127] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_130 
+ bl[128] br[128] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_131 
+ bl[129] br[129] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_132 
+ bl[130] br[130] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_133 
+ bl[131] br[131] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_134 
+ bl[132] br[132] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_135 
+ bl[133] br[133] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_136 
+ bl[134] br[134] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_137 
+ bl[135] br[135] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_138 
+ bl[136] br[136] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_139 
+ bl[137] br[137] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_140 
+ bl[138] br[138] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_141 
+ bl[139] br[139] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_142 
+ bl[140] br[140] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_143 
+ bl[141] br[141] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_144 
+ bl[142] br[142] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_145 
+ bl[143] br[143] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_146 
+ bl[144] br[144] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_147 
+ bl[145] br[145] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_148 
+ bl[146] br[146] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_149 
+ bl[147] br[147] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_150 
+ bl[148] br[148] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_151 
+ bl[149] br[149] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_152 
+ bl[150] br[150] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_153 
+ bl[151] br[151] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_154 
+ bl[152] br[152] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_155 
+ bl[153] br[153] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_156 
+ bl[154] br[154] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_157 
+ bl[155] br[155] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_158 
+ bl[156] br[156] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_159 
+ bl[157] br[157] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_160 
+ bl[158] br[158] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_161 
+ bl[159] br[159] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_162 
+ bl[160] br[160] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_163 
+ bl[161] br[161] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_164 
+ bl[162] br[162] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_165 
+ bl[163] br[163] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_166 
+ bl[164] br[164] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_167 
+ bl[165] br[165] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_168 
+ bl[166] br[166] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_169 
+ bl[167] br[167] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_170 
+ bl[168] br[168] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_171 
+ bl[169] br[169] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_172 
+ bl[170] br[170] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_173 
+ bl[171] br[171] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_174 
+ bl[172] br[172] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_175 
+ bl[173] br[173] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_176 
+ bl[174] br[174] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_177 
+ bl[175] br[175] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_178 
+ bl[176] br[176] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_179 
+ bl[177] br[177] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_180 
+ bl[178] br[178] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_181 
+ bl[179] br[179] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_182 
+ bl[180] br[180] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_183 
+ bl[181] br[181] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_184 
+ bl[182] br[182] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_185 
+ bl[183] br[183] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_186 
+ bl[184] br[184] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_187 
+ bl[185] br[185] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_188 
+ bl[186] br[186] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_189 
+ bl[187] br[187] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_190 
+ bl[188] br[188] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_191 
+ bl[189] br[189] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_192 
+ bl[190] br[190] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_193 
+ bl[191] br[191] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_194 
+ bl[192] br[192] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_195 
+ bl[193] br[193] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_196 
+ bl[194] br[194] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_197 
+ bl[195] br[195] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_198 
+ bl[196] br[196] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_199 
+ bl[197] br[197] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_200 
+ bl[198] br[198] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_201 
+ bl[199] br[199] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_202 
+ bl[200] br[200] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_203 
+ bl[201] br[201] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_204 
+ bl[202] br[202] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_205 
+ bl[203] br[203] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_206 
+ bl[204] br[204] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_207 
+ bl[205] br[205] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_208 
+ bl[206] br[206] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_209 
+ bl[207] br[207] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_210 
+ bl[208] br[208] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_211 
+ bl[209] br[209] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_212 
+ bl[210] br[210] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_213 
+ bl[211] br[211] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_214 
+ bl[212] br[212] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_215 
+ bl[213] br[213] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_216 
+ bl[214] br[214] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_217 
+ bl[215] br[215] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_218 
+ bl[216] br[216] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_219 
+ bl[217] br[217] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_220 
+ bl[218] br[218] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_221 
+ bl[219] br[219] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_222 
+ bl[220] br[220] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_223 
+ bl[221] br[221] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_224 
+ bl[222] br[222] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_225 
+ bl[223] br[223] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_226 
+ bl[224] br[224] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_227 
+ bl[225] br[225] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_228 
+ bl[226] br[226] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_229 
+ bl[227] br[227] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_230 
+ bl[228] br[228] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_231 
+ bl[229] br[229] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_232 
+ bl[230] br[230] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_233 
+ bl[231] br[231] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_234 
+ bl[232] br[232] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_235 
+ bl[233] br[233] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_236 
+ bl[234] br[234] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_237 
+ bl[235] br[235] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_238 
+ bl[236] br[236] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_239 
+ bl[237] br[237] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_240 
+ bl[238] br[238] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_241 
+ bl[239] br[239] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_242 
+ bl[240] br[240] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_243 
+ bl[241] br[241] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_244 
+ bl[242] br[242] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_245 
+ bl[243] br[243] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_246 
+ bl[244] br[244] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_247 
+ bl[245] br[245] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_248 
+ bl[246] br[246] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_249 
+ bl[247] br[247] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_250 
+ bl[248] br[248] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_251 
+ bl[249] br[249] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_252 
+ bl[250] br[250] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_253 
+ bl[251] br[251] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_254 
+ bl[252] br[252] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_255 
+ bl[253] br[253] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_256 
+ bl[254] br[254] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_257 
+ bl[255] br[255] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_258 
+ vdd vdd vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_259 
+ vdd vdd vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_0 
+ vdd vdd vss vdd vpb vnb wl[79] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_81_1 
+ rbl rbr vss vdd vpb vnb wl[79] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_81_2 
+ bl[0] br[0] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_3 
+ bl[1] br[1] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_4 
+ bl[2] br[2] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_5 
+ bl[3] br[3] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_6 
+ bl[4] br[4] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_7 
+ bl[5] br[5] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_8 
+ bl[6] br[6] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_9 
+ bl[7] br[7] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_10 
+ bl[8] br[8] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_11 
+ bl[9] br[9] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_12 
+ bl[10] br[10] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_13 
+ bl[11] br[11] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_14 
+ bl[12] br[12] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_15 
+ bl[13] br[13] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_16 
+ bl[14] br[14] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_17 
+ bl[15] br[15] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_18 
+ bl[16] br[16] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_19 
+ bl[17] br[17] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_20 
+ bl[18] br[18] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_21 
+ bl[19] br[19] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_22 
+ bl[20] br[20] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_23 
+ bl[21] br[21] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_24 
+ bl[22] br[22] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_25 
+ bl[23] br[23] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_26 
+ bl[24] br[24] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_27 
+ bl[25] br[25] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_28 
+ bl[26] br[26] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_29 
+ bl[27] br[27] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_30 
+ bl[28] br[28] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_31 
+ bl[29] br[29] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_32 
+ bl[30] br[30] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_33 
+ bl[31] br[31] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_34 
+ bl[32] br[32] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_35 
+ bl[33] br[33] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_36 
+ bl[34] br[34] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_37 
+ bl[35] br[35] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_38 
+ bl[36] br[36] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_39 
+ bl[37] br[37] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_40 
+ bl[38] br[38] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_41 
+ bl[39] br[39] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_42 
+ bl[40] br[40] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_43 
+ bl[41] br[41] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_44 
+ bl[42] br[42] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_45 
+ bl[43] br[43] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_46 
+ bl[44] br[44] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_47 
+ bl[45] br[45] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_48 
+ bl[46] br[46] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_49 
+ bl[47] br[47] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_50 
+ bl[48] br[48] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_51 
+ bl[49] br[49] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_52 
+ bl[50] br[50] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_53 
+ bl[51] br[51] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_54 
+ bl[52] br[52] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_55 
+ bl[53] br[53] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_56 
+ bl[54] br[54] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_57 
+ bl[55] br[55] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_58 
+ bl[56] br[56] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_59 
+ bl[57] br[57] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_60 
+ bl[58] br[58] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_61 
+ bl[59] br[59] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_62 
+ bl[60] br[60] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_63 
+ bl[61] br[61] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_64 
+ bl[62] br[62] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_65 
+ bl[63] br[63] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_66 
+ bl[64] br[64] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_67 
+ bl[65] br[65] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_68 
+ bl[66] br[66] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_69 
+ bl[67] br[67] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_70 
+ bl[68] br[68] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_71 
+ bl[69] br[69] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_72 
+ bl[70] br[70] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_73 
+ bl[71] br[71] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_74 
+ bl[72] br[72] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_75 
+ bl[73] br[73] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_76 
+ bl[74] br[74] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_77 
+ bl[75] br[75] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_78 
+ bl[76] br[76] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_79 
+ bl[77] br[77] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_80 
+ bl[78] br[78] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_81 
+ bl[79] br[79] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_82 
+ bl[80] br[80] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_83 
+ bl[81] br[81] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_84 
+ bl[82] br[82] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_85 
+ bl[83] br[83] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_86 
+ bl[84] br[84] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_87 
+ bl[85] br[85] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_88 
+ bl[86] br[86] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_89 
+ bl[87] br[87] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_90 
+ bl[88] br[88] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_91 
+ bl[89] br[89] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_92 
+ bl[90] br[90] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_93 
+ bl[91] br[91] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_94 
+ bl[92] br[92] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_95 
+ bl[93] br[93] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_96 
+ bl[94] br[94] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_97 
+ bl[95] br[95] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_98 
+ bl[96] br[96] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_99 
+ bl[97] br[97] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_100 
+ bl[98] br[98] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_101 
+ bl[99] br[99] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_102 
+ bl[100] br[100] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_103 
+ bl[101] br[101] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_104 
+ bl[102] br[102] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_105 
+ bl[103] br[103] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_106 
+ bl[104] br[104] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_107 
+ bl[105] br[105] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_108 
+ bl[106] br[106] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_109 
+ bl[107] br[107] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_110 
+ bl[108] br[108] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_111 
+ bl[109] br[109] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_112 
+ bl[110] br[110] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_113 
+ bl[111] br[111] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_114 
+ bl[112] br[112] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_115 
+ bl[113] br[113] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_116 
+ bl[114] br[114] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_117 
+ bl[115] br[115] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_118 
+ bl[116] br[116] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_119 
+ bl[117] br[117] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_120 
+ bl[118] br[118] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_121 
+ bl[119] br[119] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_122 
+ bl[120] br[120] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_123 
+ bl[121] br[121] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_124 
+ bl[122] br[122] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_125 
+ bl[123] br[123] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_126 
+ bl[124] br[124] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_127 
+ bl[125] br[125] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_128 
+ bl[126] br[126] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_129 
+ bl[127] br[127] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_130 
+ bl[128] br[128] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_131 
+ bl[129] br[129] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_132 
+ bl[130] br[130] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_133 
+ bl[131] br[131] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_134 
+ bl[132] br[132] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_135 
+ bl[133] br[133] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_136 
+ bl[134] br[134] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_137 
+ bl[135] br[135] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_138 
+ bl[136] br[136] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_139 
+ bl[137] br[137] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_140 
+ bl[138] br[138] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_141 
+ bl[139] br[139] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_142 
+ bl[140] br[140] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_143 
+ bl[141] br[141] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_144 
+ bl[142] br[142] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_145 
+ bl[143] br[143] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_146 
+ bl[144] br[144] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_147 
+ bl[145] br[145] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_148 
+ bl[146] br[146] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_149 
+ bl[147] br[147] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_150 
+ bl[148] br[148] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_151 
+ bl[149] br[149] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_152 
+ bl[150] br[150] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_153 
+ bl[151] br[151] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_154 
+ bl[152] br[152] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_155 
+ bl[153] br[153] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_156 
+ bl[154] br[154] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_157 
+ bl[155] br[155] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_158 
+ bl[156] br[156] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_159 
+ bl[157] br[157] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_160 
+ bl[158] br[158] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_161 
+ bl[159] br[159] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_162 
+ bl[160] br[160] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_163 
+ bl[161] br[161] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_164 
+ bl[162] br[162] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_165 
+ bl[163] br[163] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_166 
+ bl[164] br[164] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_167 
+ bl[165] br[165] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_168 
+ bl[166] br[166] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_169 
+ bl[167] br[167] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_170 
+ bl[168] br[168] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_171 
+ bl[169] br[169] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_172 
+ bl[170] br[170] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_173 
+ bl[171] br[171] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_174 
+ bl[172] br[172] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_175 
+ bl[173] br[173] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_176 
+ bl[174] br[174] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_177 
+ bl[175] br[175] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_178 
+ bl[176] br[176] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_179 
+ bl[177] br[177] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_180 
+ bl[178] br[178] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_181 
+ bl[179] br[179] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_182 
+ bl[180] br[180] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_183 
+ bl[181] br[181] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_184 
+ bl[182] br[182] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_185 
+ bl[183] br[183] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_186 
+ bl[184] br[184] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_187 
+ bl[185] br[185] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_188 
+ bl[186] br[186] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_189 
+ bl[187] br[187] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_190 
+ bl[188] br[188] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_191 
+ bl[189] br[189] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_192 
+ bl[190] br[190] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_193 
+ bl[191] br[191] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_194 
+ bl[192] br[192] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_195 
+ bl[193] br[193] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_196 
+ bl[194] br[194] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_197 
+ bl[195] br[195] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_198 
+ bl[196] br[196] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_199 
+ bl[197] br[197] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_200 
+ bl[198] br[198] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_201 
+ bl[199] br[199] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_202 
+ bl[200] br[200] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_203 
+ bl[201] br[201] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_204 
+ bl[202] br[202] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_205 
+ bl[203] br[203] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_206 
+ bl[204] br[204] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_207 
+ bl[205] br[205] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_208 
+ bl[206] br[206] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_209 
+ bl[207] br[207] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_210 
+ bl[208] br[208] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_211 
+ bl[209] br[209] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_212 
+ bl[210] br[210] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_213 
+ bl[211] br[211] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_214 
+ bl[212] br[212] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_215 
+ bl[213] br[213] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_216 
+ bl[214] br[214] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_217 
+ bl[215] br[215] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_218 
+ bl[216] br[216] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_219 
+ bl[217] br[217] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_220 
+ bl[218] br[218] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_221 
+ bl[219] br[219] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_222 
+ bl[220] br[220] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_223 
+ bl[221] br[221] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_224 
+ bl[222] br[222] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_225 
+ bl[223] br[223] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_226 
+ bl[224] br[224] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_227 
+ bl[225] br[225] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_228 
+ bl[226] br[226] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_229 
+ bl[227] br[227] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_230 
+ bl[228] br[228] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_231 
+ bl[229] br[229] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_232 
+ bl[230] br[230] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_233 
+ bl[231] br[231] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_234 
+ bl[232] br[232] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_235 
+ bl[233] br[233] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_236 
+ bl[234] br[234] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_237 
+ bl[235] br[235] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_238 
+ bl[236] br[236] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_239 
+ bl[237] br[237] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_240 
+ bl[238] br[238] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_241 
+ bl[239] br[239] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_242 
+ bl[240] br[240] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_243 
+ bl[241] br[241] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_244 
+ bl[242] br[242] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_245 
+ bl[243] br[243] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_246 
+ bl[244] br[244] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_247 
+ bl[245] br[245] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_248 
+ bl[246] br[246] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_249 
+ bl[247] br[247] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_250 
+ bl[248] br[248] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_251 
+ bl[249] br[249] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_252 
+ bl[250] br[250] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_253 
+ bl[251] br[251] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_254 
+ bl[252] br[252] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_255 
+ bl[253] br[253] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_256 
+ bl[254] br[254] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_257 
+ bl[255] br[255] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_258 
+ vdd vdd vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_259 
+ vdd vdd vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_0 
+ vdd vdd vss vdd vpb vnb wl[80] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_82_1 
+ rbl rbr vss vdd vpb vnb wl[80] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_82_2 
+ bl[0] br[0] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_3 
+ bl[1] br[1] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_4 
+ bl[2] br[2] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_5 
+ bl[3] br[3] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_6 
+ bl[4] br[4] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_7 
+ bl[5] br[5] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_8 
+ bl[6] br[6] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_9 
+ bl[7] br[7] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_10 
+ bl[8] br[8] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_11 
+ bl[9] br[9] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_12 
+ bl[10] br[10] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_13 
+ bl[11] br[11] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_14 
+ bl[12] br[12] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_15 
+ bl[13] br[13] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_16 
+ bl[14] br[14] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_17 
+ bl[15] br[15] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_18 
+ bl[16] br[16] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_19 
+ bl[17] br[17] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_20 
+ bl[18] br[18] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_21 
+ bl[19] br[19] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_22 
+ bl[20] br[20] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_23 
+ bl[21] br[21] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_24 
+ bl[22] br[22] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_25 
+ bl[23] br[23] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_26 
+ bl[24] br[24] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_27 
+ bl[25] br[25] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_28 
+ bl[26] br[26] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_29 
+ bl[27] br[27] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_30 
+ bl[28] br[28] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_31 
+ bl[29] br[29] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_32 
+ bl[30] br[30] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_33 
+ bl[31] br[31] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_34 
+ bl[32] br[32] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_35 
+ bl[33] br[33] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_36 
+ bl[34] br[34] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_37 
+ bl[35] br[35] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_38 
+ bl[36] br[36] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_39 
+ bl[37] br[37] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_40 
+ bl[38] br[38] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_41 
+ bl[39] br[39] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_42 
+ bl[40] br[40] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_43 
+ bl[41] br[41] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_44 
+ bl[42] br[42] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_45 
+ bl[43] br[43] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_46 
+ bl[44] br[44] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_47 
+ bl[45] br[45] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_48 
+ bl[46] br[46] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_49 
+ bl[47] br[47] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_50 
+ bl[48] br[48] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_51 
+ bl[49] br[49] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_52 
+ bl[50] br[50] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_53 
+ bl[51] br[51] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_54 
+ bl[52] br[52] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_55 
+ bl[53] br[53] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_56 
+ bl[54] br[54] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_57 
+ bl[55] br[55] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_58 
+ bl[56] br[56] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_59 
+ bl[57] br[57] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_60 
+ bl[58] br[58] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_61 
+ bl[59] br[59] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_62 
+ bl[60] br[60] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_63 
+ bl[61] br[61] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_64 
+ bl[62] br[62] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_65 
+ bl[63] br[63] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_66 
+ bl[64] br[64] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_67 
+ bl[65] br[65] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_68 
+ bl[66] br[66] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_69 
+ bl[67] br[67] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_70 
+ bl[68] br[68] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_71 
+ bl[69] br[69] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_72 
+ bl[70] br[70] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_73 
+ bl[71] br[71] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_74 
+ bl[72] br[72] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_75 
+ bl[73] br[73] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_76 
+ bl[74] br[74] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_77 
+ bl[75] br[75] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_78 
+ bl[76] br[76] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_79 
+ bl[77] br[77] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_80 
+ bl[78] br[78] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_81 
+ bl[79] br[79] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_82 
+ bl[80] br[80] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_83 
+ bl[81] br[81] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_84 
+ bl[82] br[82] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_85 
+ bl[83] br[83] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_86 
+ bl[84] br[84] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_87 
+ bl[85] br[85] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_88 
+ bl[86] br[86] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_89 
+ bl[87] br[87] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_90 
+ bl[88] br[88] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_91 
+ bl[89] br[89] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_92 
+ bl[90] br[90] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_93 
+ bl[91] br[91] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_94 
+ bl[92] br[92] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_95 
+ bl[93] br[93] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_96 
+ bl[94] br[94] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_97 
+ bl[95] br[95] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_98 
+ bl[96] br[96] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_99 
+ bl[97] br[97] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_100 
+ bl[98] br[98] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_101 
+ bl[99] br[99] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_102 
+ bl[100] br[100] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_103 
+ bl[101] br[101] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_104 
+ bl[102] br[102] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_105 
+ bl[103] br[103] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_106 
+ bl[104] br[104] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_107 
+ bl[105] br[105] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_108 
+ bl[106] br[106] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_109 
+ bl[107] br[107] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_110 
+ bl[108] br[108] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_111 
+ bl[109] br[109] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_112 
+ bl[110] br[110] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_113 
+ bl[111] br[111] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_114 
+ bl[112] br[112] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_115 
+ bl[113] br[113] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_116 
+ bl[114] br[114] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_117 
+ bl[115] br[115] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_118 
+ bl[116] br[116] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_119 
+ bl[117] br[117] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_120 
+ bl[118] br[118] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_121 
+ bl[119] br[119] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_122 
+ bl[120] br[120] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_123 
+ bl[121] br[121] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_124 
+ bl[122] br[122] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_125 
+ bl[123] br[123] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_126 
+ bl[124] br[124] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_127 
+ bl[125] br[125] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_128 
+ bl[126] br[126] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_129 
+ bl[127] br[127] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_130 
+ bl[128] br[128] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_131 
+ bl[129] br[129] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_132 
+ bl[130] br[130] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_133 
+ bl[131] br[131] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_134 
+ bl[132] br[132] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_135 
+ bl[133] br[133] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_136 
+ bl[134] br[134] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_137 
+ bl[135] br[135] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_138 
+ bl[136] br[136] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_139 
+ bl[137] br[137] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_140 
+ bl[138] br[138] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_141 
+ bl[139] br[139] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_142 
+ bl[140] br[140] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_143 
+ bl[141] br[141] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_144 
+ bl[142] br[142] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_145 
+ bl[143] br[143] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_146 
+ bl[144] br[144] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_147 
+ bl[145] br[145] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_148 
+ bl[146] br[146] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_149 
+ bl[147] br[147] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_150 
+ bl[148] br[148] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_151 
+ bl[149] br[149] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_152 
+ bl[150] br[150] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_153 
+ bl[151] br[151] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_154 
+ bl[152] br[152] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_155 
+ bl[153] br[153] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_156 
+ bl[154] br[154] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_157 
+ bl[155] br[155] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_158 
+ bl[156] br[156] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_159 
+ bl[157] br[157] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_160 
+ bl[158] br[158] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_161 
+ bl[159] br[159] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_162 
+ bl[160] br[160] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_163 
+ bl[161] br[161] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_164 
+ bl[162] br[162] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_165 
+ bl[163] br[163] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_166 
+ bl[164] br[164] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_167 
+ bl[165] br[165] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_168 
+ bl[166] br[166] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_169 
+ bl[167] br[167] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_170 
+ bl[168] br[168] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_171 
+ bl[169] br[169] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_172 
+ bl[170] br[170] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_173 
+ bl[171] br[171] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_174 
+ bl[172] br[172] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_175 
+ bl[173] br[173] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_176 
+ bl[174] br[174] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_177 
+ bl[175] br[175] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_178 
+ bl[176] br[176] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_179 
+ bl[177] br[177] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_180 
+ bl[178] br[178] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_181 
+ bl[179] br[179] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_182 
+ bl[180] br[180] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_183 
+ bl[181] br[181] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_184 
+ bl[182] br[182] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_185 
+ bl[183] br[183] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_186 
+ bl[184] br[184] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_187 
+ bl[185] br[185] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_188 
+ bl[186] br[186] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_189 
+ bl[187] br[187] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_190 
+ bl[188] br[188] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_191 
+ bl[189] br[189] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_192 
+ bl[190] br[190] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_193 
+ bl[191] br[191] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_194 
+ bl[192] br[192] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_195 
+ bl[193] br[193] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_196 
+ bl[194] br[194] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_197 
+ bl[195] br[195] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_198 
+ bl[196] br[196] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_199 
+ bl[197] br[197] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_200 
+ bl[198] br[198] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_201 
+ bl[199] br[199] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_202 
+ bl[200] br[200] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_203 
+ bl[201] br[201] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_204 
+ bl[202] br[202] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_205 
+ bl[203] br[203] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_206 
+ bl[204] br[204] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_207 
+ bl[205] br[205] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_208 
+ bl[206] br[206] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_209 
+ bl[207] br[207] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_210 
+ bl[208] br[208] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_211 
+ bl[209] br[209] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_212 
+ bl[210] br[210] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_213 
+ bl[211] br[211] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_214 
+ bl[212] br[212] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_215 
+ bl[213] br[213] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_216 
+ bl[214] br[214] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_217 
+ bl[215] br[215] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_218 
+ bl[216] br[216] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_219 
+ bl[217] br[217] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_220 
+ bl[218] br[218] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_221 
+ bl[219] br[219] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_222 
+ bl[220] br[220] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_223 
+ bl[221] br[221] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_224 
+ bl[222] br[222] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_225 
+ bl[223] br[223] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_226 
+ bl[224] br[224] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_227 
+ bl[225] br[225] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_228 
+ bl[226] br[226] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_229 
+ bl[227] br[227] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_230 
+ bl[228] br[228] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_231 
+ bl[229] br[229] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_232 
+ bl[230] br[230] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_233 
+ bl[231] br[231] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_234 
+ bl[232] br[232] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_235 
+ bl[233] br[233] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_236 
+ bl[234] br[234] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_237 
+ bl[235] br[235] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_238 
+ bl[236] br[236] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_239 
+ bl[237] br[237] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_240 
+ bl[238] br[238] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_241 
+ bl[239] br[239] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_242 
+ bl[240] br[240] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_243 
+ bl[241] br[241] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_244 
+ bl[242] br[242] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_245 
+ bl[243] br[243] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_246 
+ bl[244] br[244] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_247 
+ bl[245] br[245] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_248 
+ bl[246] br[246] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_249 
+ bl[247] br[247] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_250 
+ bl[248] br[248] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_251 
+ bl[249] br[249] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_252 
+ bl[250] br[250] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_253 
+ bl[251] br[251] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_254 
+ bl[252] br[252] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_255 
+ bl[253] br[253] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_256 
+ bl[254] br[254] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_257 
+ bl[255] br[255] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_258 
+ vdd vdd vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_259 
+ vdd vdd vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_0 
+ vdd vdd vss vdd vpb vnb wl[81] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_83_1 
+ rbl rbr vss vdd vpb vnb wl[81] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_83_2 
+ bl[0] br[0] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_3 
+ bl[1] br[1] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_4 
+ bl[2] br[2] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_5 
+ bl[3] br[3] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_6 
+ bl[4] br[4] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_7 
+ bl[5] br[5] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_8 
+ bl[6] br[6] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_9 
+ bl[7] br[7] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_10 
+ bl[8] br[8] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_11 
+ bl[9] br[9] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_12 
+ bl[10] br[10] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_13 
+ bl[11] br[11] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_14 
+ bl[12] br[12] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_15 
+ bl[13] br[13] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_16 
+ bl[14] br[14] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_17 
+ bl[15] br[15] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_18 
+ bl[16] br[16] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_19 
+ bl[17] br[17] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_20 
+ bl[18] br[18] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_21 
+ bl[19] br[19] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_22 
+ bl[20] br[20] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_23 
+ bl[21] br[21] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_24 
+ bl[22] br[22] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_25 
+ bl[23] br[23] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_26 
+ bl[24] br[24] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_27 
+ bl[25] br[25] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_28 
+ bl[26] br[26] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_29 
+ bl[27] br[27] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_30 
+ bl[28] br[28] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_31 
+ bl[29] br[29] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_32 
+ bl[30] br[30] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_33 
+ bl[31] br[31] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_34 
+ bl[32] br[32] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_35 
+ bl[33] br[33] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_36 
+ bl[34] br[34] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_37 
+ bl[35] br[35] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_38 
+ bl[36] br[36] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_39 
+ bl[37] br[37] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_40 
+ bl[38] br[38] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_41 
+ bl[39] br[39] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_42 
+ bl[40] br[40] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_43 
+ bl[41] br[41] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_44 
+ bl[42] br[42] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_45 
+ bl[43] br[43] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_46 
+ bl[44] br[44] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_47 
+ bl[45] br[45] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_48 
+ bl[46] br[46] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_49 
+ bl[47] br[47] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_50 
+ bl[48] br[48] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_51 
+ bl[49] br[49] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_52 
+ bl[50] br[50] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_53 
+ bl[51] br[51] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_54 
+ bl[52] br[52] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_55 
+ bl[53] br[53] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_56 
+ bl[54] br[54] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_57 
+ bl[55] br[55] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_58 
+ bl[56] br[56] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_59 
+ bl[57] br[57] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_60 
+ bl[58] br[58] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_61 
+ bl[59] br[59] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_62 
+ bl[60] br[60] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_63 
+ bl[61] br[61] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_64 
+ bl[62] br[62] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_65 
+ bl[63] br[63] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_66 
+ bl[64] br[64] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_67 
+ bl[65] br[65] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_68 
+ bl[66] br[66] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_69 
+ bl[67] br[67] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_70 
+ bl[68] br[68] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_71 
+ bl[69] br[69] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_72 
+ bl[70] br[70] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_73 
+ bl[71] br[71] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_74 
+ bl[72] br[72] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_75 
+ bl[73] br[73] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_76 
+ bl[74] br[74] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_77 
+ bl[75] br[75] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_78 
+ bl[76] br[76] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_79 
+ bl[77] br[77] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_80 
+ bl[78] br[78] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_81 
+ bl[79] br[79] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_82 
+ bl[80] br[80] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_83 
+ bl[81] br[81] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_84 
+ bl[82] br[82] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_85 
+ bl[83] br[83] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_86 
+ bl[84] br[84] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_87 
+ bl[85] br[85] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_88 
+ bl[86] br[86] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_89 
+ bl[87] br[87] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_90 
+ bl[88] br[88] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_91 
+ bl[89] br[89] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_92 
+ bl[90] br[90] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_93 
+ bl[91] br[91] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_94 
+ bl[92] br[92] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_95 
+ bl[93] br[93] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_96 
+ bl[94] br[94] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_97 
+ bl[95] br[95] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_98 
+ bl[96] br[96] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_99 
+ bl[97] br[97] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_100 
+ bl[98] br[98] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_101 
+ bl[99] br[99] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_102 
+ bl[100] br[100] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_103 
+ bl[101] br[101] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_104 
+ bl[102] br[102] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_105 
+ bl[103] br[103] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_106 
+ bl[104] br[104] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_107 
+ bl[105] br[105] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_108 
+ bl[106] br[106] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_109 
+ bl[107] br[107] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_110 
+ bl[108] br[108] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_111 
+ bl[109] br[109] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_112 
+ bl[110] br[110] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_113 
+ bl[111] br[111] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_114 
+ bl[112] br[112] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_115 
+ bl[113] br[113] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_116 
+ bl[114] br[114] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_117 
+ bl[115] br[115] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_118 
+ bl[116] br[116] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_119 
+ bl[117] br[117] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_120 
+ bl[118] br[118] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_121 
+ bl[119] br[119] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_122 
+ bl[120] br[120] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_123 
+ bl[121] br[121] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_124 
+ bl[122] br[122] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_125 
+ bl[123] br[123] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_126 
+ bl[124] br[124] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_127 
+ bl[125] br[125] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_128 
+ bl[126] br[126] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_129 
+ bl[127] br[127] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_130 
+ bl[128] br[128] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_131 
+ bl[129] br[129] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_132 
+ bl[130] br[130] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_133 
+ bl[131] br[131] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_134 
+ bl[132] br[132] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_135 
+ bl[133] br[133] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_136 
+ bl[134] br[134] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_137 
+ bl[135] br[135] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_138 
+ bl[136] br[136] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_139 
+ bl[137] br[137] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_140 
+ bl[138] br[138] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_141 
+ bl[139] br[139] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_142 
+ bl[140] br[140] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_143 
+ bl[141] br[141] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_144 
+ bl[142] br[142] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_145 
+ bl[143] br[143] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_146 
+ bl[144] br[144] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_147 
+ bl[145] br[145] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_148 
+ bl[146] br[146] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_149 
+ bl[147] br[147] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_150 
+ bl[148] br[148] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_151 
+ bl[149] br[149] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_152 
+ bl[150] br[150] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_153 
+ bl[151] br[151] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_154 
+ bl[152] br[152] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_155 
+ bl[153] br[153] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_156 
+ bl[154] br[154] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_157 
+ bl[155] br[155] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_158 
+ bl[156] br[156] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_159 
+ bl[157] br[157] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_160 
+ bl[158] br[158] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_161 
+ bl[159] br[159] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_162 
+ bl[160] br[160] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_163 
+ bl[161] br[161] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_164 
+ bl[162] br[162] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_165 
+ bl[163] br[163] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_166 
+ bl[164] br[164] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_167 
+ bl[165] br[165] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_168 
+ bl[166] br[166] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_169 
+ bl[167] br[167] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_170 
+ bl[168] br[168] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_171 
+ bl[169] br[169] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_172 
+ bl[170] br[170] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_173 
+ bl[171] br[171] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_174 
+ bl[172] br[172] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_175 
+ bl[173] br[173] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_176 
+ bl[174] br[174] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_177 
+ bl[175] br[175] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_178 
+ bl[176] br[176] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_179 
+ bl[177] br[177] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_180 
+ bl[178] br[178] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_181 
+ bl[179] br[179] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_182 
+ bl[180] br[180] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_183 
+ bl[181] br[181] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_184 
+ bl[182] br[182] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_185 
+ bl[183] br[183] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_186 
+ bl[184] br[184] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_187 
+ bl[185] br[185] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_188 
+ bl[186] br[186] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_189 
+ bl[187] br[187] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_190 
+ bl[188] br[188] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_191 
+ bl[189] br[189] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_192 
+ bl[190] br[190] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_193 
+ bl[191] br[191] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_194 
+ bl[192] br[192] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_195 
+ bl[193] br[193] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_196 
+ bl[194] br[194] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_197 
+ bl[195] br[195] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_198 
+ bl[196] br[196] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_199 
+ bl[197] br[197] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_200 
+ bl[198] br[198] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_201 
+ bl[199] br[199] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_202 
+ bl[200] br[200] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_203 
+ bl[201] br[201] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_204 
+ bl[202] br[202] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_205 
+ bl[203] br[203] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_206 
+ bl[204] br[204] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_207 
+ bl[205] br[205] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_208 
+ bl[206] br[206] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_209 
+ bl[207] br[207] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_210 
+ bl[208] br[208] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_211 
+ bl[209] br[209] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_212 
+ bl[210] br[210] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_213 
+ bl[211] br[211] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_214 
+ bl[212] br[212] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_215 
+ bl[213] br[213] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_216 
+ bl[214] br[214] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_217 
+ bl[215] br[215] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_218 
+ bl[216] br[216] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_219 
+ bl[217] br[217] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_220 
+ bl[218] br[218] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_221 
+ bl[219] br[219] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_222 
+ bl[220] br[220] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_223 
+ bl[221] br[221] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_224 
+ bl[222] br[222] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_225 
+ bl[223] br[223] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_226 
+ bl[224] br[224] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_227 
+ bl[225] br[225] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_228 
+ bl[226] br[226] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_229 
+ bl[227] br[227] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_230 
+ bl[228] br[228] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_231 
+ bl[229] br[229] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_232 
+ bl[230] br[230] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_233 
+ bl[231] br[231] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_234 
+ bl[232] br[232] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_235 
+ bl[233] br[233] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_236 
+ bl[234] br[234] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_237 
+ bl[235] br[235] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_238 
+ bl[236] br[236] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_239 
+ bl[237] br[237] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_240 
+ bl[238] br[238] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_241 
+ bl[239] br[239] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_242 
+ bl[240] br[240] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_243 
+ bl[241] br[241] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_244 
+ bl[242] br[242] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_245 
+ bl[243] br[243] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_246 
+ bl[244] br[244] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_247 
+ bl[245] br[245] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_248 
+ bl[246] br[246] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_249 
+ bl[247] br[247] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_250 
+ bl[248] br[248] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_251 
+ bl[249] br[249] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_252 
+ bl[250] br[250] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_253 
+ bl[251] br[251] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_254 
+ bl[252] br[252] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_255 
+ bl[253] br[253] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_256 
+ bl[254] br[254] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_257 
+ bl[255] br[255] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_258 
+ vdd vdd vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_259 
+ vdd vdd vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_0 
+ vdd vdd vss vdd vpb vnb wl[82] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_84_1 
+ rbl rbr vss vdd vpb vnb wl[82] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_84_2 
+ bl[0] br[0] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_3 
+ bl[1] br[1] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_4 
+ bl[2] br[2] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_5 
+ bl[3] br[3] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_6 
+ bl[4] br[4] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_7 
+ bl[5] br[5] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_8 
+ bl[6] br[6] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_9 
+ bl[7] br[7] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_10 
+ bl[8] br[8] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_11 
+ bl[9] br[9] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_12 
+ bl[10] br[10] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_13 
+ bl[11] br[11] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_14 
+ bl[12] br[12] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_15 
+ bl[13] br[13] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_16 
+ bl[14] br[14] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_17 
+ bl[15] br[15] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_18 
+ bl[16] br[16] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_19 
+ bl[17] br[17] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_20 
+ bl[18] br[18] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_21 
+ bl[19] br[19] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_22 
+ bl[20] br[20] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_23 
+ bl[21] br[21] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_24 
+ bl[22] br[22] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_25 
+ bl[23] br[23] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_26 
+ bl[24] br[24] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_27 
+ bl[25] br[25] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_28 
+ bl[26] br[26] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_29 
+ bl[27] br[27] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_30 
+ bl[28] br[28] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_31 
+ bl[29] br[29] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_32 
+ bl[30] br[30] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_33 
+ bl[31] br[31] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_34 
+ bl[32] br[32] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_35 
+ bl[33] br[33] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_36 
+ bl[34] br[34] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_37 
+ bl[35] br[35] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_38 
+ bl[36] br[36] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_39 
+ bl[37] br[37] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_40 
+ bl[38] br[38] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_41 
+ bl[39] br[39] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_42 
+ bl[40] br[40] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_43 
+ bl[41] br[41] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_44 
+ bl[42] br[42] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_45 
+ bl[43] br[43] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_46 
+ bl[44] br[44] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_47 
+ bl[45] br[45] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_48 
+ bl[46] br[46] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_49 
+ bl[47] br[47] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_50 
+ bl[48] br[48] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_51 
+ bl[49] br[49] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_52 
+ bl[50] br[50] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_53 
+ bl[51] br[51] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_54 
+ bl[52] br[52] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_55 
+ bl[53] br[53] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_56 
+ bl[54] br[54] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_57 
+ bl[55] br[55] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_58 
+ bl[56] br[56] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_59 
+ bl[57] br[57] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_60 
+ bl[58] br[58] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_61 
+ bl[59] br[59] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_62 
+ bl[60] br[60] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_63 
+ bl[61] br[61] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_64 
+ bl[62] br[62] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_65 
+ bl[63] br[63] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_66 
+ bl[64] br[64] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_67 
+ bl[65] br[65] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_68 
+ bl[66] br[66] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_69 
+ bl[67] br[67] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_70 
+ bl[68] br[68] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_71 
+ bl[69] br[69] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_72 
+ bl[70] br[70] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_73 
+ bl[71] br[71] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_74 
+ bl[72] br[72] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_75 
+ bl[73] br[73] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_76 
+ bl[74] br[74] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_77 
+ bl[75] br[75] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_78 
+ bl[76] br[76] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_79 
+ bl[77] br[77] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_80 
+ bl[78] br[78] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_81 
+ bl[79] br[79] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_82 
+ bl[80] br[80] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_83 
+ bl[81] br[81] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_84 
+ bl[82] br[82] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_85 
+ bl[83] br[83] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_86 
+ bl[84] br[84] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_87 
+ bl[85] br[85] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_88 
+ bl[86] br[86] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_89 
+ bl[87] br[87] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_90 
+ bl[88] br[88] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_91 
+ bl[89] br[89] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_92 
+ bl[90] br[90] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_93 
+ bl[91] br[91] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_94 
+ bl[92] br[92] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_95 
+ bl[93] br[93] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_96 
+ bl[94] br[94] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_97 
+ bl[95] br[95] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_98 
+ bl[96] br[96] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_99 
+ bl[97] br[97] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_100 
+ bl[98] br[98] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_101 
+ bl[99] br[99] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_102 
+ bl[100] br[100] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_103 
+ bl[101] br[101] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_104 
+ bl[102] br[102] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_105 
+ bl[103] br[103] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_106 
+ bl[104] br[104] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_107 
+ bl[105] br[105] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_108 
+ bl[106] br[106] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_109 
+ bl[107] br[107] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_110 
+ bl[108] br[108] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_111 
+ bl[109] br[109] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_112 
+ bl[110] br[110] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_113 
+ bl[111] br[111] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_114 
+ bl[112] br[112] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_115 
+ bl[113] br[113] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_116 
+ bl[114] br[114] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_117 
+ bl[115] br[115] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_118 
+ bl[116] br[116] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_119 
+ bl[117] br[117] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_120 
+ bl[118] br[118] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_121 
+ bl[119] br[119] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_122 
+ bl[120] br[120] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_123 
+ bl[121] br[121] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_124 
+ bl[122] br[122] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_125 
+ bl[123] br[123] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_126 
+ bl[124] br[124] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_127 
+ bl[125] br[125] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_128 
+ bl[126] br[126] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_129 
+ bl[127] br[127] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_130 
+ bl[128] br[128] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_131 
+ bl[129] br[129] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_132 
+ bl[130] br[130] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_133 
+ bl[131] br[131] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_134 
+ bl[132] br[132] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_135 
+ bl[133] br[133] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_136 
+ bl[134] br[134] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_137 
+ bl[135] br[135] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_138 
+ bl[136] br[136] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_139 
+ bl[137] br[137] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_140 
+ bl[138] br[138] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_141 
+ bl[139] br[139] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_142 
+ bl[140] br[140] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_143 
+ bl[141] br[141] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_144 
+ bl[142] br[142] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_145 
+ bl[143] br[143] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_146 
+ bl[144] br[144] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_147 
+ bl[145] br[145] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_148 
+ bl[146] br[146] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_149 
+ bl[147] br[147] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_150 
+ bl[148] br[148] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_151 
+ bl[149] br[149] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_152 
+ bl[150] br[150] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_153 
+ bl[151] br[151] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_154 
+ bl[152] br[152] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_155 
+ bl[153] br[153] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_156 
+ bl[154] br[154] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_157 
+ bl[155] br[155] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_158 
+ bl[156] br[156] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_159 
+ bl[157] br[157] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_160 
+ bl[158] br[158] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_161 
+ bl[159] br[159] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_162 
+ bl[160] br[160] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_163 
+ bl[161] br[161] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_164 
+ bl[162] br[162] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_165 
+ bl[163] br[163] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_166 
+ bl[164] br[164] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_167 
+ bl[165] br[165] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_168 
+ bl[166] br[166] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_169 
+ bl[167] br[167] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_170 
+ bl[168] br[168] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_171 
+ bl[169] br[169] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_172 
+ bl[170] br[170] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_173 
+ bl[171] br[171] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_174 
+ bl[172] br[172] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_175 
+ bl[173] br[173] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_176 
+ bl[174] br[174] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_177 
+ bl[175] br[175] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_178 
+ bl[176] br[176] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_179 
+ bl[177] br[177] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_180 
+ bl[178] br[178] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_181 
+ bl[179] br[179] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_182 
+ bl[180] br[180] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_183 
+ bl[181] br[181] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_184 
+ bl[182] br[182] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_185 
+ bl[183] br[183] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_186 
+ bl[184] br[184] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_187 
+ bl[185] br[185] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_188 
+ bl[186] br[186] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_189 
+ bl[187] br[187] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_190 
+ bl[188] br[188] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_191 
+ bl[189] br[189] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_192 
+ bl[190] br[190] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_193 
+ bl[191] br[191] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_194 
+ bl[192] br[192] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_195 
+ bl[193] br[193] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_196 
+ bl[194] br[194] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_197 
+ bl[195] br[195] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_198 
+ bl[196] br[196] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_199 
+ bl[197] br[197] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_200 
+ bl[198] br[198] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_201 
+ bl[199] br[199] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_202 
+ bl[200] br[200] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_203 
+ bl[201] br[201] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_204 
+ bl[202] br[202] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_205 
+ bl[203] br[203] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_206 
+ bl[204] br[204] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_207 
+ bl[205] br[205] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_208 
+ bl[206] br[206] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_209 
+ bl[207] br[207] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_210 
+ bl[208] br[208] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_211 
+ bl[209] br[209] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_212 
+ bl[210] br[210] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_213 
+ bl[211] br[211] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_214 
+ bl[212] br[212] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_215 
+ bl[213] br[213] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_216 
+ bl[214] br[214] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_217 
+ bl[215] br[215] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_218 
+ bl[216] br[216] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_219 
+ bl[217] br[217] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_220 
+ bl[218] br[218] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_221 
+ bl[219] br[219] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_222 
+ bl[220] br[220] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_223 
+ bl[221] br[221] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_224 
+ bl[222] br[222] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_225 
+ bl[223] br[223] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_226 
+ bl[224] br[224] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_227 
+ bl[225] br[225] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_228 
+ bl[226] br[226] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_229 
+ bl[227] br[227] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_230 
+ bl[228] br[228] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_231 
+ bl[229] br[229] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_232 
+ bl[230] br[230] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_233 
+ bl[231] br[231] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_234 
+ bl[232] br[232] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_235 
+ bl[233] br[233] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_236 
+ bl[234] br[234] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_237 
+ bl[235] br[235] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_238 
+ bl[236] br[236] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_239 
+ bl[237] br[237] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_240 
+ bl[238] br[238] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_241 
+ bl[239] br[239] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_242 
+ bl[240] br[240] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_243 
+ bl[241] br[241] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_244 
+ bl[242] br[242] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_245 
+ bl[243] br[243] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_246 
+ bl[244] br[244] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_247 
+ bl[245] br[245] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_248 
+ bl[246] br[246] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_249 
+ bl[247] br[247] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_250 
+ bl[248] br[248] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_251 
+ bl[249] br[249] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_252 
+ bl[250] br[250] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_253 
+ bl[251] br[251] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_254 
+ bl[252] br[252] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_255 
+ bl[253] br[253] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_256 
+ bl[254] br[254] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_257 
+ bl[255] br[255] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_258 
+ vdd vdd vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_259 
+ vdd vdd vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_0 
+ vdd vdd vss vdd vpb vnb wl[83] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_85_1 
+ rbl rbr vss vdd vpb vnb wl[83] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_85_2 
+ bl[0] br[0] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_3 
+ bl[1] br[1] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_4 
+ bl[2] br[2] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_5 
+ bl[3] br[3] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_6 
+ bl[4] br[4] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_7 
+ bl[5] br[5] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_8 
+ bl[6] br[6] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_9 
+ bl[7] br[7] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_10 
+ bl[8] br[8] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_11 
+ bl[9] br[9] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_12 
+ bl[10] br[10] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_13 
+ bl[11] br[11] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_14 
+ bl[12] br[12] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_15 
+ bl[13] br[13] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_16 
+ bl[14] br[14] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_17 
+ bl[15] br[15] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_18 
+ bl[16] br[16] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_19 
+ bl[17] br[17] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_20 
+ bl[18] br[18] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_21 
+ bl[19] br[19] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_22 
+ bl[20] br[20] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_23 
+ bl[21] br[21] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_24 
+ bl[22] br[22] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_25 
+ bl[23] br[23] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_26 
+ bl[24] br[24] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_27 
+ bl[25] br[25] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_28 
+ bl[26] br[26] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_29 
+ bl[27] br[27] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_30 
+ bl[28] br[28] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_31 
+ bl[29] br[29] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_32 
+ bl[30] br[30] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_33 
+ bl[31] br[31] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_34 
+ bl[32] br[32] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_35 
+ bl[33] br[33] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_36 
+ bl[34] br[34] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_37 
+ bl[35] br[35] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_38 
+ bl[36] br[36] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_39 
+ bl[37] br[37] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_40 
+ bl[38] br[38] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_41 
+ bl[39] br[39] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_42 
+ bl[40] br[40] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_43 
+ bl[41] br[41] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_44 
+ bl[42] br[42] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_45 
+ bl[43] br[43] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_46 
+ bl[44] br[44] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_47 
+ bl[45] br[45] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_48 
+ bl[46] br[46] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_49 
+ bl[47] br[47] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_50 
+ bl[48] br[48] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_51 
+ bl[49] br[49] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_52 
+ bl[50] br[50] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_53 
+ bl[51] br[51] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_54 
+ bl[52] br[52] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_55 
+ bl[53] br[53] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_56 
+ bl[54] br[54] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_57 
+ bl[55] br[55] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_58 
+ bl[56] br[56] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_59 
+ bl[57] br[57] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_60 
+ bl[58] br[58] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_61 
+ bl[59] br[59] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_62 
+ bl[60] br[60] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_63 
+ bl[61] br[61] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_64 
+ bl[62] br[62] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_65 
+ bl[63] br[63] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_66 
+ bl[64] br[64] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_67 
+ bl[65] br[65] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_68 
+ bl[66] br[66] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_69 
+ bl[67] br[67] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_70 
+ bl[68] br[68] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_71 
+ bl[69] br[69] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_72 
+ bl[70] br[70] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_73 
+ bl[71] br[71] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_74 
+ bl[72] br[72] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_75 
+ bl[73] br[73] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_76 
+ bl[74] br[74] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_77 
+ bl[75] br[75] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_78 
+ bl[76] br[76] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_79 
+ bl[77] br[77] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_80 
+ bl[78] br[78] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_81 
+ bl[79] br[79] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_82 
+ bl[80] br[80] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_83 
+ bl[81] br[81] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_84 
+ bl[82] br[82] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_85 
+ bl[83] br[83] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_86 
+ bl[84] br[84] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_87 
+ bl[85] br[85] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_88 
+ bl[86] br[86] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_89 
+ bl[87] br[87] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_90 
+ bl[88] br[88] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_91 
+ bl[89] br[89] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_92 
+ bl[90] br[90] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_93 
+ bl[91] br[91] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_94 
+ bl[92] br[92] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_95 
+ bl[93] br[93] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_96 
+ bl[94] br[94] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_97 
+ bl[95] br[95] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_98 
+ bl[96] br[96] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_99 
+ bl[97] br[97] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_100 
+ bl[98] br[98] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_101 
+ bl[99] br[99] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_102 
+ bl[100] br[100] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_103 
+ bl[101] br[101] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_104 
+ bl[102] br[102] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_105 
+ bl[103] br[103] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_106 
+ bl[104] br[104] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_107 
+ bl[105] br[105] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_108 
+ bl[106] br[106] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_109 
+ bl[107] br[107] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_110 
+ bl[108] br[108] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_111 
+ bl[109] br[109] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_112 
+ bl[110] br[110] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_113 
+ bl[111] br[111] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_114 
+ bl[112] br[112] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_115 
+ bl[113] br[113] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_116 
+ bl[114] br[114] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_117 
+ bl[115] br[115] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_118 
+ bl[116] br[116] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_119 
+ bl[117] br[117] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_120 
+ bl[118] br[118] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_121 
+ bl[119] br[119] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_122 
+ bl[120] br[120] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_123 
+ bl[121] br[121] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_124 
+ bl[122] br[122] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_125 
+ bl[123] br[123] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_126 
+ bl[124] br[124] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_127 
+ bl[125] br[125] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_128 
+ bl[126] br[126] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_129 
+ bl[127] br[127] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_130 
+ bl[128] br[128] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_131 
+ bl[129] br[129] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_132 
+ bl[130] br[130] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_133 
+ bl[131] br[131] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_134 
+ bl[132] br[132] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_135 
+ bl[133] br[133] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_136 
+ bl[134] br[134] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_137 
+ bl[135] br[135] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_138 
+ bl[136] br[136] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_139 
+ bl[137] br[137] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_140 
+ bl[138] br[138] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_141 
+ bl[139] br[139] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_142 
+ bl[140] br[140] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_143 
+ bl[141] br[141] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_144 
+ bl[142] br[142] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_145 
+ bl[143] br[143] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_146 
+ bl[144] br[144] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_147 
+ bl[145] br[145] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_148 
+ bl[146] br[146] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_149 
+ bl[147] br[147] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_150 
+ bl[148] br[148] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_151 
+ bl[149] br[149] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_152 
+ bl[150] br[150] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_153 
+ bl[151] br[151] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_154 
+ bl[152] br[152] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_155 
+ bl[153] br[153] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_156 
+ bl[154] br[154] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_157 
+ bl[155] br[155] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_158 
+ bl[156] br[156] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_159 
+ bl[157] br[157] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_160 
+ bl[158] br[158] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_161 
+ bl[159] br[159] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_162 
+ bl[160] br[160] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_163 
+ bl[161] br[161] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_164 
+ bl[162] br[162] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_165 
+ bl[163] br[163] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_166 
+ bl[164] br[164] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_167 
+ bl[165] br[165] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_168 
+ bl[166] br[166] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_169 
+ bl[167] br[167] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_170 
+ bl[168] br[168] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_171 
+ bl[169] br[169] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_172 
+ bl[170] br[170] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_173 
+ bl[171] br[171] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_174 
+ bl[172] br[172] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_175 
+ bl[173] br[173] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_176 
+ bl[174] br[174] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_177 
+ bl[175] br[175] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_178 
+ bl[176] br[176] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_179 
+ bl[177] br[177] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_180 
+ bl[178] br[178] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_181 
+ bl[179] br[179] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_182 
+ bl[180] br[180] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_183 
+ bl[181] br[181] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_184 
+ bl[182] br[182] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_185 
+ bl[183] br[183] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_186 
+ bl[184] br[184] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_187 
+ bl[185] br[185] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_188 
+ bl[186] br[186] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_189 
+ bl[187] br[187] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_190 
+ bl[188] br[188] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_191 
+ bl[189] br[189] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_192 
+ bl[190] br[190] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_193 
+ bl[191] br[191] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_194 
+ bl[192] br[192] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_195 
+ bl[193] br[193] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_196 
+ bl[194] br[194] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_197 
+ bl[195] br[195] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_198 
+ bl[196] br[196] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_199 
+ bl[197] br[197] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_200 
+ bl[198] br[198] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_201 
+ bl[199] br[199] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_202 
+ bl[200] br[200] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_203 
+ bl[201] br[201] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_204 
+ bl[202] br[202] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_205 
+ bl[203] br[203] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_206 
+ bl[204] br[204] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_207 
+ bl[205] br[205] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_208 
+ bl[206] br[206] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_209 
+ bl[207] br[207] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_210 
+ bl[208] br[208] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_211 
+ bl[209] br[209] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_212 
+ bl[210] br[210] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_213 
+ bl[211] br[211] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_214 
+ bl[212] br[212] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_215 
+ bl[213] br[213] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_216 
+ bl[214] br[214] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_217 
+ bl[215] br[215] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_218 
+ bl[216] br[216] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_219 
+ bl[217] br[217] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_220 
+ bl[218] br[218] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_221 
+ bl[219] br[219] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_222 
+ bl[220] br[220] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_223 
+ bl[221] br[221] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_224 
+ bl[222] br[222] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_225 
+ bl[223] br[223] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_226 
+ bl[224] br[224] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_227 
+ bl[225] br[225] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_228 
+ bl[226] br[226] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_229 
+ bl[227] br[227] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_230 
+ bl[228] br[228] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_231 
+ bl[229] br[229] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_232 
+ bl[230] br[230] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_233 
+ bl[231] br[231] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_234 
+ bl[232] br[232] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_235 
+ bl[233] br[233] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_236 
+ bl[234] br[234] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_237 
+ bl[235] br[235] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_238 
+ bl[236] br[236] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_239 
+ bl[237] br[237] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_240 
+ bl[238] br[238] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_241 
+ bl[239] br[239] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_242 
+ bl[240] br[240] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_243 
+ bl[241] br[241] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_244 
+ bl[242] br[242] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_245 
+ bl[243] br[243] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_246 
+ bl[244] br[244] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_247 
+ bl[245] br[245] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_248 
+ bl[246] br[246] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_249 
+ bl[247] br[247] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_250 
+ bl[248] br[248] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_251 
+ bl[249] br[249] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_252 
+ bl[250] br[250] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_253 
+ bl[251] br[251] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_254 
+ bl[252] br[252] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_255 
+ bl[253] br[253] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_256 
+ bl[254] br[254] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_257 
+ bl[255] br[255] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_258 
+ vdd vdd vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_259 
+ vdd vdd vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_0 
+ vdd vdd vss vdd vpb vnb wl[84] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_86_1 
+ rbl rbr vss vdd vpb vnb wl[84] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_86_2 
+ bl[0] br[0] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_3 
+ bl[1] br[1] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_4 
+ bl[2] br[2] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_5 
+ bl[3] br[3] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_6 
+ bl[4] br[4] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_7 
+ bl[5] br[5] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_8 
+ bl[6] br[6] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_9 
+ bl[7] br[7] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_10 
+ bl[8] br[8] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_11 
+ bl[9] br[9] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_12 
+ bl[10] br[10] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_13 
+ bl[11] br[11] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_14 
+ bl[12] br[12] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_15 
+ bl[13] br[13] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_16 
+ bl[14] br[14] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_17 
+ bl[15] br[15] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_18 
+ bl[16] br[16] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_19 
+ bl[17] br[17] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_20 
+ bl[18] br[18] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_21 
+ bl[19] br[19] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_22 
+ bl[20] br[20] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_23 
+ bl[21] br[21] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_24 
+ bl[22] br[22] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_25 
+ bl[23] br[23] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_26 
+ bl[24] br[24] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_27 
+ bl[25] br[25] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_28 
+ bl[26] br[26] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_29 
+ bl[27] br[27] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_30 
+ bl[28] br[28] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_31 
+ bl[29] br[29] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_32 
+ bl[30] br[30] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_33 
+ bl[31] br[31] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_34 
+ bl[32] br[32] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_35 
+ bl[33] br[33] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_36 
+ bl[34] br[34] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_37 
+ bl[35] br[35] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_38 
+ bl[36] br[36] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_39 
+ bl[37] br[37] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_40 
+ bl[38] br[38] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_41 
+ bl[39] br[39] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_42 
+ bl[40] br[40] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_43 
+ bl[41] br[41] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_44 
+ bl[42] br[42] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_45 
+ bl[43] br[43] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_46 
+ bl[44] br[44] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_47 
+ bl[45] br[45] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_48 
+ bl[46] br[46] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_49 
+ bl[47] br[47] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_50 
+ bl[48] br[48] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_51 
+ bl[49] br[49] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_52 
+ bl[50] br[50] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_53 
+ bl[51] br[51] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_54 
+ bl[52] br[52] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_55 
+ bl[53] br[53] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_56 
+ bl[54] br[54] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_57 
+ bl[55] br[55] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_58 
+ bl[56] br[56] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_59 
+ bl[57] br[57] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_60 
+ bl[58] br[58] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_61 
+ bl[59] br[59] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_62 
+ bl[60] br[60] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_63 
+ bl[61] br[61] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_64 
+ bl[62] br[62] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_65 
+ bl[63] br[63] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_66 
+ bl[64] br[64] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_67 
+ bl[65] br[65] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_68 
+ bl[66] br[66] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_69 
+ bl[67] br[67] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_70 
+ bl[68] br[68] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_71 
+ bl[69] br[69] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_72 
+ bl[70] br[70] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_73 
+ bl[71] br[71] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_74 
+ bl[72] br[72] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_75 
+ bl[73] br[73] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_76 
+ bl[74] br[74] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_77 
+ bl[75] br[75] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_78 
+ bl[76] br[76] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_79 
+ bl[77] br[77] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_80 
+ bl[78] br[78] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_81 
+ bl[79] br[79] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_82 
+ bl[80] br[80] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_83 
+ bl[81] br[81] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_84 
+ bl[82] br[82] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_85 
+ bl[83] br[83] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_86 
+ bl[84] br[84] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_87 
+ bl[85] br[85] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_88 
+ bl[86] br[86] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_89 
+ bl[87] br[87] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_90 
+ bl[88] br[88] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_91 
+ bl[89] br[89] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_92 
+ bl[90] br[90] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_93 
+ bl[91] br[91] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_94 
+ bl[92] br[92] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_95 
+ bl[93] br[93] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_96 
+ bl[94] br[94] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_97 
+ bl[95] br[95] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_98 
+ bl[96] br[96] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_99 
+ bl[97] br[97] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_100 
+ bl[98] br[98] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_101 
+ bl[99] br[99] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_102 
+ bl[100] br[100] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_103 
+ bl[101] br[101] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_104 
+ bl[102] br[102] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_105 
+ bl[103] br[103] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_106 
+ bl[104] br[104] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_107 
+ bl[105] br[105] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_108 
+ bl[106] br[106] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_109 
+ bl[107] br[107] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_110 
+ bl[108] br[108] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_111 
+ bl[109] br[109] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_112 
+ bl[110] br[110] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_113 
+ bl[111] br[111] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_114 
+ bl[112] br[112] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_115 
+ bl[113] br[113] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_116 
+ bl[114] br[114] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_117 
+ bl[115] br[115] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_118 
+ bl[116] br[116] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_119 
+ bl[117] br[117] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_120 
+ bl[118] br[118] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_121 
+ bl[119] br[119] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_122 
+ bl[120] br[120] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_123 
+ bl[121] br[121] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_124 
+ bl[122] br[122] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_125 
+ bl[123] br[123] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_126 
+ bl[124] br[124] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_127 
+ bl[125] br[125] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_128 
+ bl[126] br[126] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_129 
+ bl[127] br[127] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_130 
+ bl[128] br[128] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_131 
+ bl[129] br[129] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_132 
+ bl[130] br[130] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_133 
+ bl[131] br[131] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_134 
+ bl[132] br[132] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_135 
+ bl[133] br[133] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_136 
+ bl[134] br[134] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_137 
+ bl[135] br[135] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_138 
+ bl[136] br[136] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_139 
+ bl[137] br[137] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_140 
+ bl[138] br[138] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_141 
+ bl[139] br[139] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_142 
+ bl[140] br[140] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_143 
+ bl[141] br[141] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_144 
+ bl[142] br[142] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_145 
+ bl[143] br[143] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_146 
+ bl[144] br[144] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_147 
+ bl[145] br[145] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_148 
+ bl[146] br[146] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_149 
+ bl[147] br[147] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_150 
+ bl[148] br[148] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_151 
+ bl[149] br[149] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_152 
+ bl[150] br[150] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_153 
+ bl[151] br[151] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_154 
+ bl[152] br[152] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_155 
+ bl[153] br[153] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_156 
+ bl[154] br[154] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_157 
+ bl[155] br[155] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_158 
+ bl[156] br[156] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_159 
+ bl[157] br[157] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_160 
+ bl[158] br[158] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_161 
+ bl[159] br[159] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_162 
+ bl[160] br[160] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_163 
+ bl[161] br[161] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_164 
+ bl[162] br[162] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_165 
+ bl[163] br[163] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_166 
+ bl[164] br[164] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_167 
+ bl[165] br[165] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_168 
+ bl[166] br[166] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_169 
+ bl[167] br[167] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_170 
+ bl[168] br[168] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_171 
+ bl[169] br[169] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_172 
+ bl[170] br[170] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_173 
+ bl[171] br[171] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_174 
+ bl[172] br[172] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_175 
+ bl[173] br[173] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_176 
+ bl[174] br[174] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_177 
+ bl[175] br[175] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_178 
+ bl[176] br[176] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_179 
+ bl[177] br[177] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_180 
+ bl[178] br[178] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_181 
+ bl[179] br[179] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_182 
+ bl[180] br[180] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_183 
+ bl[181] br[181] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_184 
+ bl[182] br[182] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_185 
+ bl[183] br[183] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_186 
+ bl[184] br[184] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_187 
+ bl[185] br[185] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_188 
+ bl[186] br[186] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_189 
+ bl[187] br[187] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_190 
+ bl[188] br[188] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_191 
+ bl[189] br[189] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_192 
+ bl[190] br[190] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_193 
+ bl[191] br[191] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_194 
+ bl[192] br[192] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_195 
+ bl[193] br[193] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_196 
+ bl[194] br[194] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_197 
+ bl[195] br[195] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_198 
+ bl[196] br[196] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_199 
+ bl[197] br[197] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_200 
+ bl[198] br[198] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_201 
+ bl[199] br[199] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_202 
+ bl[200] br[200] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_203 
+ bl[201] br[201] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_204 
+ bl[202] br[202] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_205 
+ bl[203] br[203] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_206 
+ bl[204] br[204] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_207 
+ bl[205] br[205] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_208 
+ bl[206] br[206] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_209 
+ bl[207] br[207] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_210 
+ bl[208] br[208] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_211 
+ bl[209] br[209] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_212 
+ bl[210] br[210] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_213 
+ bl[211] br[211] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_214 
+ bl[212] br[212] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_215 
+ bl[213] br[213] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_216 
+ bl[214] br[214] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_217 
+ bl[215] br[215] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_218 
+ bl[216] br[216] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_219 
+ bl[217] br[217] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_220 
+ bl[218] br[218] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_221 
+ bl[219] br[219] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_222 
+ bl[220] br[220] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_223 
+ bl[221] br[221] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_224 
+ bl[222] br[222] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_225 
+ bl[223] br[223] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_226 
+ bl[224] br[224] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_227 
+ bl[225] br[225] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_228 
+ bl[226] br[226] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_229 
+ bl[227] br[227] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_230 
+ bl[228] br[228] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_231 
+ bl[229] br[229] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_232 
+ bl[230] br[230] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_233 
+ bl[231] br[231] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_234 
+ bl[232] br[232] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_235 
+ bl[233] br[233] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_236 
+ bl[234] br[234] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_237 
+ bl[235] br[235] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_238 
+ bl[236] br[236] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_239 
+ bl[237] br[237] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_240 
+ bl[238] br[238] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_241 
+ bl[239] br[239] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_242 
+ bl[240] br[240] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_243 
+ bl[241] br[241] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_244 
+ bl[242] br[242] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_245 
+ bl[243] br[243] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_246 
+ bl[244] br[244] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_247 
+ bl[245] br[245] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_248 
+ bl[246] br[246] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_249 
+ bl[247] br[247] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_250 
+ bl[248] br[248] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_251 
+ bl[249] br[249] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_252 
+ bl[250] br[250] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_253 
+ bl[251] br[251] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_254 
+ bl[252] br[252] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_255 
+ bl[253] br[253] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_256 
+ bl[254] br[254] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_257 
+ bl[255] br[255] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_258 
+ vdd vdd vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_259 
+ vdd vdd vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_0 
+ vdd vdd vss vdd vpb vnb wl[85] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_87_1 
+ rbl rbr vss vdd vpb vnb wl[85] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_87_2 
+ bl[0] br[0] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_3 
+ bl[1] br[1] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_4 
+ bl[2] br[2] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_5 
+ bl[3] br[3] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_6 
+ bl[4] br[4] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_7 
+ bl[5] br[5] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_8 
+ bl[6] br[6] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_9 
+ bl[7] br[7] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_10 
+ bl[8] br[8] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_11 
+ bl[9] br[9] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_12 
+ bl[10] br[10] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_13 
+ bl[11] br[11] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_14 
+ bl[12] br[12] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_15 
+ bl[13] br[13] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_16 
+ bl[14] br[14] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_17 
+ bl[15] br[15] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_18 
+ bl[16] br[16] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_19 
+ bl[17] br[17] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_20 
+ bl[18] br[18] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_21 
+ bl[19] br[19] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_22 
+ bl[20] br[20] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_23 
+ bl[21] br[21] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_24 
+ bl[22] br[22] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_25 
+ bl[23] br[23] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_26 
+ bl[24] br[24] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_27 
+ bl[25] br[25] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_28 
+ bl[26] br[26] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_29 
+ bl[27] br[27] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_30 
+ bl[28] br[28] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_31 
+ bl[29] br[29] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_32 
+ bl[30] br[30] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_33 
+ bl[31] br[31] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_34 
+ bl[32] br[32] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_35 
+ bl[33] br[33] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_36 
+ bl[34] br[34] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_37 
+ bl[35] br[35] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_38 
+ bl[36] br[36] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_39 
+ bl[37] br[37] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_40 
+ bl[38] br[38] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_41 
+ bl[39] br[39] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_42 
+ bl[40] br[40] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_43 
+ bl[41] br[41] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_44 
+ bl[42] br[42] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_45 
+ bl[43] br[43] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_46 
+ bl[44] br[44] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_47 
+ bl[45] br[45] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_48 
+ bl[46] br[46] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_49 
+ bl[47] br[47] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_50 
+ bl[48] br[48] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_51 
+ bl[49] br[49] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_52 
+ bl[50] br[50] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_53 
+ bl[51] br[51] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_54 
+ bl[52] br[52] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_55 
+ bl[53] br[53] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_56 
+ bl[54] br[54] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_57 
+ bl[55] br[55] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_58 
+ bl[56] br[56] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_59 
+ bl[57] br[57] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_60 
+ bl[58] br[58] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_61 
+ bl[59] br[59] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_62 
+ bl[60] br[60] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_63 
+ bl[61] br[61] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_64 
+ bl[62] br[62] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_65 
+ bl[63] br[63] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_66 
+ bl[64] br[64] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_67 
+ bl[65] br[65] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_68 
+ bl[66] br[66] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_69 
+ bl[67] br[67] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_70 
+ bl[68] br[68] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_71 
+ bl[69] br[69] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_72 
+ bl[70] br[70] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_73 
+ bl[71] br[71] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_74 
+ bl[72] br[72] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_75 
+ bl[73] br[73] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_76 
+ bl[74] br[74] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_77 
+ bl[75] br[75] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_78 
+ bl[76] br[76] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_79 
+ bl[77] br[77] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_80 
+ bl[78] br[78] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_81 
+ bl[79] br[79] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_82 
+ bl[80] br[80] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_83 
+ bl[81] br[81] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_84 
+ bl[82] br[82] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_85 
+ bl[83] br[83] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_86 
+ bl[84] br[84] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_87 
+ bl[85] br[85] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_88 
+ bl[86] br[86] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_89 
+ bl[87] br[87] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_90 
+ bl[88] br[88] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_91 
+ bl[89] br[89] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_92 
+ bl[90] br[90] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_93 
+ bl[91] br[91] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_94 
+ bl[92] br[92] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_95 
+ bl[93] br[93] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_96 
+ bl[94] br[94] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_97 
+ bl[95] br[95] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_98 
+ bl[96] br[96] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_99 
+ bl[97] br[97] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_100 
+ bl[98] br[98] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_101 
+ bl[99] br[99] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_102 
+ bl[100] br[100] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_103 
+ bl[101] br[101] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_104 
+ bl[102] br[102] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_105 
+ bl[103] br[103] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_106 
+ bl[104] br[104] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_107 
+ bl[105] br[105] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_108 
+ bl[106] br[106] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_109 
+ bl[107] br[107] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_110 
+ bl[108] br[108] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_111 
+ bl[109] br[109] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_112 
+ bl[110] br[110] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_113 
+ bl[111] br[111] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_114 
+ bl[112] br[112] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_115 
+ bl[113] br[113] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_116 
+ bl[114] br[114] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_117 
+ bl[115] br[115] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_118 
+ bl[116] br[116] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_119 
+ bl[117] br[117] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_120 
+ bl[118] br[118] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_121 
+ bl[119] br[119] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_122 
+ bl[120] br[120] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_123 
+ bl[121] br[121] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_124 
+ bl[122] br[122] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_125 
+ bl[123] br[123] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_126 
+ bl[124] br[124] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_127 
+ bl[125] br[125] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_128 
+ bl[126] br[126] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_129 
+ bl[127] br[127] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_130 
+ bl[128] br[128] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_131 
+ bl[129] br[129] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_132 
+ bl[130] br[130] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_133 
+ bl[131] br[131] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_134 
+ bl[132] br[132] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_135 
+ bl[133] br[133] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_136 
+ bl[134] br[134] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_137 
+ bl[135] br[135] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_138 
+ bl[136] br[136] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_139 
+ bl[137] br[137] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_140 
+ bl[138] br[138] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_141 
+ bl[139] br[139] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_142 
+ bl[140] br[140] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_143 
+ bl[141] br[141] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_144 
+ bl[142] br[142] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_145 
+ bl[143] br[143] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_146 
+ bl[144] br[144] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_147 
+ bl[145] br[145] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_148 
+ bl[146] br[146] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_149 
+ bl[147] br[147] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_150 
+ bl[148] br[148] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_151 
+ bl[149] br[149] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_152 
+ bl[150] br[150] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_153 
+ bl[151] br[151] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_154 
+ bl[152] br[152] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_155 
+ bl[153] br[153] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_156 
+ bl[154] br[154] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_157 
+ bl[155] br[155] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_158 
+ bl[156] br[156] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_159 
+ bl[157] br[157] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_160 
+ bl[158] br[158] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_161 
+ bl[159] br[159] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_162 
+ bl[160] br[160] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_163 
+ bl[161] br[161] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_164 
+ bl[162] br[162] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_165 
+ bl[163] br[163] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_166 
+ bl[164] br[164] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_167 
+ bl[165] br[165] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_168 
+ bl[166] br[166] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_169 
+ bl[167] br[167] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_170 
+ bl[168] br[168] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_171 
+ bl[169] br[169] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_172 
+ bl[170] br[170] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_173 
+ bl[171] br[171] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_174 
+ bl[172] br[172] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_175 
+ bl[173] br[173] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_176 
+ bl[174] br[174] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_177 
+ bl[175] br[175] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_178 
+ bl[176] br[176] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_179 
+ bl[177] br[177] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_180 
+ bl[178] br[178] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_181 
+ bl[179] br[179] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_182 
+ bl[180] br[180] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_183 
+ bl[181] br[181] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_184 
+ bl[182] br[182] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_185 
+ bl[183] br[183] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_186 
+ bl[184] br[184] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_187 
+ bl[185] br[185] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_188 
+ bl[186] br[186] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_189 
+ bl[187] br[187] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_190 
+ bl[188] br[188] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_191 
+ bl[189] br[189] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_192 
+ bl[190] br[190] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_193 
+ bl[191] br[191] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_194 
+ bl[192] br[192] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_195 
+ bl[193] br[193] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_196 
+ bl[194] br[194] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_197 
+ bl[195] br[195] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_198 
+ bl[196] br[196] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_199 
+ bl[197] br[197] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_200 
+ bl[198] br[198] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_201 
+ bl[199] br[199] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_202 
+ bl[200] br[200] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_203 
+ bl[201] br[201] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_204 
+ bl[202] br[202] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_205 
+ bl[203] br[203] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_206 
+ bl[204] br[204] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_207 
+ bl[205] br[205] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_208 
+ bl[206] br[206] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_209 
+ bl[207] br[207] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_210 
+ bl[208] br[208] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_211 
+ bl[209] br[209] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_212 
+ bl[210] br[210] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_213 
+ bl[211] br[211] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_214 
+ bl[212] br[212] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_215 
+ bl[213] br[213] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_216 
+ bl[214] br[214] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_217 
+ bl[215] br[215] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_218 
+ bl[216] br[216] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_219 
+ bl[217] br[217] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_220 
+ bl[218] br[218] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_221 
+ bl[219] br[219] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_222 
+ bl[220] br[220] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_223 
+ bl[221] br[221] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_224 
+ bl[222] br[222] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_225 
+ bl[223] br[223] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_226 
+ bl[224] br[224] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_227 
+ bl[225] br[225] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_228 
+ bl[226] br[226] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_229 
+ bl[227] br[227] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_230 
+ bl[228] br[228] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_231 
+ bl[229] br[229] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_232 
+ bl[230] br[230] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_233 
+ bl[231] br[231] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_234 
+ bl[232] br[232] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_235 
+ bl[233] br[233] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_236 
+ bl[234] br[234] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_237 
+ bl[235] br[235] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_238 
+ bl[236] br[236] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_239 
+ bl[237] br[237] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_240 
+ bl[238] br[238] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_241 
+ bl[239] br[239] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_242 
+ bl[240] br[240] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_243 
+ bl[241] br[241] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_244 
+ bl[242] br[242] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_245 
+ bl[243] br[243] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_246 
+ bl[244] br[244] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_247 
+ bl[245] br[245] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_248 
+ bl[246] br[246] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_249 
+ bl[247] br[247] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_250 
+ bl[248] br[248] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_251 
+ bl[249] br[249] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_252 
+ bl[250] br[250] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_253 
+ bl[251] br[251] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_254 
+ bl[252] br[252] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_255 
+ bl[253] br[253] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_256 
+ bl[254] br[254] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_257 
+ bl[255] br[255] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_258 
+ vdd vdd vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_259 
+ vdd vdd vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_0 
+ vdd vdd vss vdd vpb vnb wl[86] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_88_1 
+ rbl rbr vss vdd vpb vnb wl[86] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_88_2 
+ bl[0] br[0] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_3 
+ bl[1] br[1] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_4 
+ bl[2] br[2] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_5 
+ bl[3] br[3] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_6 
+ bl[4] br[4] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_7 
+ bl[5] br[5] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_8 
+ bl[6] br[6] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_9 
+ bl[7] br[7] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_10 
+ bl[8] br[8] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_11 
+ bl[9] br[9] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_12 
+ bl[10] br[10] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_13 
+ bl[11] br[11] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_14 
+ bl[12] br[12] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_15 
+ bl[13] br[13] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_16 
+ bl[14] br[14] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_17 
+ bl[15] br[15] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_18 
+ bl[16] br[16] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_19 
+ bl[17] br[17] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_20 
+ bl[18] br[18] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_21 
+ bl[19] br[19] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_22 
+ bl[20] br[20] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_23 
+ bl[21] br[21] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_24 
+ bl[22] br[22] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_25 
+ bl[23] br[23] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_26 
+ bl[24] br[24] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_27 
+ bl[25] br[25] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_28 
+ bl[26] br[26] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_29 
+ bl[27] br[27] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_30 
+ bl[28] br[28] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_31 
+ bl[29] br[29] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_32 
+ bl[30] br[30] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_33 
+ bl[31] br[31] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_34 
+ bl[32] br[32] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_35 
+ bl[33] br[33] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_36 
+ bl[34] br[34] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_37 
+ bl[35] br[35] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_38 
+ bl[36] br[36] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_39 
+ bl[37] br[37] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_40 
+ bl[38] br[38] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_41 
+ bl[39] br[39] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_42 
+ bl[40] br[40] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_43 
+ bl[41] br[41] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_44 
+ bl[42] br[42] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_45 
+ bl[43] br[43] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_46 
+ bl[44] br[44] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_47 
+ bl[45] br[45] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_48 
+ bl[46] br[46] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_49 
+ bl[47] br[47] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_50 
+ bl[48] br[48] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_51 
+ bl[49] br[49] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_52 
+ bl[50] br[50] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_53 
+ bl[51] br[51] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_54 
+ bl[52] br[52] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_55 
+ bl[53] br[53] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_56 
+ bl[54] br[54] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_57 
+ bl[55] br[55] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_58 
+ bl[56] br[56] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_59 
+ bl[57] br[57] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_60 
+ bl[58] br[58] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_61 
+ bl[59] br[59] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_62 
+ bl[60] br[60] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_63 
+ bl[61] br[61] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_64 
+ bl[62] br[62] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_65 
+ bl[63] br[63] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_66 
+ bl[64] br[64] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_67 
+ bl[65] br[65] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_68 
+ bl[66] br[66] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_69 
+ bl[67] br[67] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_70 
+ bl[68] br[68] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_71 
+ bl[69] br[69] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_72 
+ bl[70] br[70] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_73 
+ bl[71] br[71] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_74 
+ bl[72] br[72] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_75 
+ bl[73] br[73] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_76 
+ bl[74] br[74] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_77 
+ bl[75] br[75] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_78 
+ bl[76] br[76] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_79 
+ bl[77] br[77] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_80 
+ bl[78] br[78] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_81 
+ bl[79] br[79] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_82 
+ bl[80] br[80] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_83 
+ bl[81] br[81] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_84 
+ bl[82] br[82] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_85 
+ bl[83] br[83] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_86 
+ bl[84] br[84] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_87 
+ bl[85] br[85] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_88 
+ bl[86] br[86] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_89 
+ bl[87] br[87] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_90 
+ bl[88] br[88] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_91 
+ bl[89] br[89] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_92 
+ bl[90] br[90] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_93 
+ bl[91] br[91] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_94 
+ bl[92] br[92] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_95 
+ bl[93] br[93] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_96 
+ bl[94] br[94] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_97 
+ bl[95] br[95] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_98 
+ bl[96] br[96] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_99 
+ bl[97] br[97] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_100 
+ bl[98] br[98] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_101 
+ bl[99] br[99] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_102 
+ bl[100] br[100] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_103 
+ bl[101] br[101] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_104 
+ bl[102] br[102] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_105 
+ bl[103] br[103] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_106 
+ bl[104] br[104] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_107 
+ bl[105] br[105] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_108 
+ bl[106] br[106] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_109 
+ bl[107] br[107] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_110 
+ bl[108] br[108] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_111 
+ bl[109] br[109] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_112 
+ bl[110] br[110] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_113 
+ bl[111] br[111] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_114 
+ bl[112] br[112] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_115 
+ bl[113] br[113] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_116 
+ bl[114] br[114] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_117 
+ bl[115] br[115] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_118 
+ bl[116] br[116] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_119 
+ bl[117] br[117] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_120 
+ bl[118] br[118] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_121 
+ bl[119] br[119] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_122 
+ bl[120] br[120] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_123 
+ bl[121] br[121] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_124 
+ bl[122] br[122] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_125 
+ bl[123] br[123] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_126 
+ bl[124] br[124] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_127 
+ bl[125] br[125] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_128 
+ bl[126] br[126] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_129 
+ bl[127] br[127] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_130 
+ bl[128] br[128] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_131 
+ bl[129] br[129] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_132 
+ bl[130] br[130] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_133 
+ bl[131] br[131] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_134 
+ bl[132] br[132] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_135 
+ bl[133] br[133] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_136 
+ bl[134] br[134] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_137 
+ bl[135] br[135] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_138 
+ bl[136] br[136] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_139 
+ bl[137] br[137] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_140 
+ bl[138] br[138] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_141 
+ bl[139] br[139] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_142 
+ bl[140] br[140] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_143 
+ bl[141] br[141] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_144 
+ bl[142] br[142] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_145 
+ bl[143] br[143] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_146 
+ bl[144] br[144] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_147 
+ bl[145] br[145] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_148 
+ bl[146] br[146] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_149 
+ bl[147] br[147] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_150 
+ bl[148] br[148] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_151 
+ bl[149] br[149] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_152 
+ bl[150] br[150] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_153 
+ bl[151] br[151] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_154 
+ bl[152] br[152] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_155 
+ bl[153] br[153] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_156 
+ bl[154] br[154] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_157 
+ bl[155] br[155] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_158 
+ bl[156] br[156] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_159 
+ bl[157] br[157] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_160 
+ bl[158] br[158] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_161 
+ bl[159] br[159] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_162 
+ bl[160] br[160] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_163 
+ bl[161] br[161] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_164 
+ bl[162] br[162] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_165 
+ bl[163] br[163] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_166 
+ bl[164] br[164] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_167 
+ bl[165] br[165] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_168 
+ bl[166] br[166] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_169 
+ bl[167] br[167] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_170 
+ bl[168] br[168] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_171 
+ bl[169] br[169] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_172 
+ bl[170] br[170] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_173 
+ bl[171] br[171] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_174 
+ bl[172] br[172] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_175 
+ bl[173] br[173] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_176 
+ bl[174] br[174] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_177 
+ bl[175] br[175] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_178 
+ bl[176] br[176] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_179 
+ bl[177] br[177] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_180 
+ bl[178] br[178] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_181 
+ bl[179] br[179] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_182 
+ bl[180] br[180] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_183 
+ bl[181] br[181] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_184 
+ bl[182] br[182] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_185 
+ bl[183] br[183] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_186 
+ bl[184] br[184] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_187 
+ bl[185] br[185] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_188 
+ bl[186] br[186] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_189 
+ bl[187] br[187] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_190 
+ bl[188] br[188] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_191 
+ bl[189] br[189] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_192 
+ bl[190] br[190] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_193 
+ bl[191] br[191] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_194 
+ bl[192] br[192] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_195 
+ bl[193] br[193] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_196 
+ bl[194] br[194] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_197 
+ bl[195] br[195] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_198 
+ bl[196] br[196] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_199 
+ bl[197] br[197] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_200 
+ bl[198] br[198] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_201 
+ bl[199] br[199] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_202 
+ bl[200] br[200] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_203 
+ bl[201] br[201] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_204 
+ bl[202] br[202] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_205 
+ bl[203] br[203] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_206 
+ bl[204] br[204] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_207 
+ bl[205] br[205] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_208 
+ bl[206] br[206] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_209 
+ bl[207] br[207] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_210 
+ bl[208] br[208] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_211 
+ bl[209] br[209] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_212 
+ bl[210] br[210] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_213 
+ bl[211] br[211] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_214 
+ bl[212] br[212] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_215 
+ bl[213] br[213] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_216 
+ bl[214] br[214] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_217 
+ bl[215] br[215] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_218 
+ bl[216] br[216] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_219 
+ bl[217] br[217] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_220 
+ bl[218] br[218] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_221 
+ bl[219] br[219] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_222 
+ bl[220] br[220] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_223 
+ bl[221] br[221] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_224 
+ bl[222] br[222] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_225 
+ bl[223] br[223] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_226 
+ bl[224] br[224] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_227 
+ bl[225] br[225] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_228 
+ bl[226] br[226] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_229 
+ bl[227] br[227] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_230 
+ bl[228] br[228] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_231 
+ bl[229] br[229] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_232 
+ bl[230] br[230] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_233 
+ bl[231] br[231] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_234 
+ bl[232] br[232] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_235 
+ bl[233] br[233] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_236 
+ bl[234] br[234] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_237 
+ bl[235] br[235] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_238 
+ bl[236] br[236] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_239 
+ bl[237] br[237] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_240 
+ bl[238] br[238] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_241 
+ bl[239] br[239] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_242 
+ bl[240] br[240] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_243 
+ bl[241] br[241] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_244 
+ bl[242] br[242] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_245 
+ bl[243] br[243] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_246 
+ bl[244] br[244] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_247 
+ bl[245] br[245] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_248 
+ bl[246] br[246] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_249 
+ bl[247] br[247] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_250 
+ bl[248] br[248] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_251 
+ bl[249] br[249] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_252 
+ bl[250] br[250] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_253 
+ bl[251] br[251] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_254 
+ bl[252] br[252] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_255 
+ bl[253] br[253] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_256 
+ bl[254] br[254] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_257 
+ bl[255] br[255] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_258 
+ vdd vdd vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_259 
+ vdd vdd vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_0 
+ vdd vdd vss vdd vpb vnb wl[87] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_89_1 
+ rbl rbr vss vdd vpb vnb wl[87] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_89_2 
+ bl[0] br[0] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_3 
+ bl[1] br[1] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_4 
+ bl[2] br[2] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_5 
+ bl[3] br[3] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_6 
+ bl[4] br[4] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_7 
+ bl[5] br[5] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_8 
+ bl[6] br[6] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_9 
+ bl[7] br[7] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_10 
+ bl[8] br[8] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_11 
+ bl[9] br[9] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_12 
+ bl[10] br[10] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_13 
+ bl[11] br[11] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_14 
+ bl[12] br[12] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_15 
+ bl[13] br[13] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_16 
+ bl[14] br[14] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_17 
+ bl[15] br[15] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_18 
+ bl[16] br[16] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_19 
+ bl[17] br[17] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_20 
+ bl[18] br[18] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_21 
+ bl[19] br[19] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_22 
+ bl[20] br[20] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_23 
+ bl[21] br[21] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_24 
+ bl[22] br[22] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_25 
+ bl[23] br[23] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_26 
+ bl[24] br[24] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_27 
+ bl[25] br[25] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_28 
+ bl[26] br[26] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_29 
+ bl[27] br[27] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_30 
+ bl[28] br[28] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_31 
+ bl[29] br[29] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_32 
+ bl[30] br[30] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_33 
+ bl[31] br[31] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_34 
+ bl[32] br[32] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_35 
+ bl[33] br[33] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_36 
+ bl[34] br[34] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_37 
+ bl[35] br[35] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_38 
+ bl[36] br[36] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_39 
+ bl[37] br[37] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_40 
+ bl[38] br[38] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_41 
+ bl[39] br[39] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_42 
+ bl[40] br[40] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_43 
+ bl[41] br[41] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_44 
+ bl[42] br[42] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_45 
+ bl[43] br[43] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_46 
+ bl[44] br[44] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_47 
+ bl[45] br[45] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_48 
+ bl[46] br[46] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_49 
+ bl[47] br[47] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_50 
+ bl[48] br[48] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_51 
+ bl[49] br[49] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_52 
+ bl[50] br[50] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_53 
+ bl[51] br[51] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_54 
+ bl[52] br[52] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_55 
+ bl[53] br[53] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_56 
+ bl[54] br[54] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_57 
+ bl[55] br[55] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_58 
+ bl[56] br[56] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_59 
+ bl[57] br[57] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_60 
+ bl[58] br[58] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_61 
+ bl[59] br[59] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_62 
+ bl[60] br[60] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_63 
+ bl[61] br[61] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_64 
+ bl[62] br[62] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_65 
+ bl[63] br[63] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_66 
+ bl[64] br[64] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_67 
+ bl[65] br[65] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_68 
+ bl[66] br[66] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_69 
+ bl[67] br[67] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_70 
+ bl[68] br[68] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_71 
+ bl[69] br[69] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_72 
+ bl[70] br[70] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_73 
+ bl[71] br[71] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_74 
+ bl[72] br[72] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_75 
+ bl[73] br[73] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_76 
+ bl[74] br[74] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_77 
+ bl[75] br[75] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_78 
+ bl[76] br[76] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_79 
+ bl[77] br[77] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_80 
+ bl[78] br[78] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_81 
+ bl[79] br[79] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_82 
+ bl[80] br[80] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_83 
+ bl[81] br[81] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_84 
+ bl[82] br[82] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_85 
+ bl[83] br[83] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_86 
+ bl[84] br[84] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_87 
+ bl[85] br[85] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_88 
+ bl[86] br[86] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_89 
+ bl[87] br[87] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_90 
+ bl[88] br[88] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_91 
+ bl[89] br[89] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_92 
+ bl[90] br[90] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_93 
+ bl[91] br[91] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_94 
+ bl[92] br[92] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_95 
+ bl[93] br[93] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_96 
+ bl[94] br[94] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_97 
+ bl[95] br[95] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_98 
+ bl[96] br[96] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_99 
+ bl[97] br[97] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_100 
+ bl[98] br[98] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_101 
+ bl[99] br[99] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_102 
+ bl[100] br[100] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_103 
+ bl[101] br[101] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_104 
+ bl[102] br[102] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_105 
+ bl[103] br[103] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_106 
+ bl[104] br[104] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_107 
+ bl[105] br[105] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_108 
+ bl[106] br[106] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_109 
+ bl[107] br[107] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_110 
+ bl[108] br[108] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_111 
+ bl[109] br[109] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_112 
+ bl[110] br[110] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_113 
+ bl[111] br[111] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_114 
+ bl[112] br[112] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_115 
+ bl[113] br[113] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_116 
+ bl[114] br[114] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_117 
+ bl[115] br[115] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_118 
+ bl[116] br[116] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_119 
+ bl[117] br[117] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_120 
+ bl[118] br[118] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_121 
+ bl[119] br[119] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_122 
+ bl[120] br[120] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_123 
+ bl[121] br[121] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_124 
+ bl[122] br[122] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_125 
+ bl[123] br[123] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_126 
+ bl[124] br[124] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_127 
+ bl[125] br[125] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_128 
+ bl[126] br[126] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_129 
+ bl[127] br[127] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_130 
+ bl[128] br[128] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_131 
+ bl[129] br[129] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_132 
+ bl[130] br[130] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_133 
+ bl[131] br[131] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_134 
+ bl[132] br[132] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_135 
+ bl[133] br[133] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_136 
+ bl[134] br[134] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_137 
+ bl[135] br[135] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_138 
+ bl[136] br[136] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_139 
+ bl[137] br[137] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_140 
+ bl[138] br[138] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_141 
+ bl[139] br[139] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_142 
+ bl[140] br[140] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_143 
+ bl[141] br[141] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_144 
+ bl[142] br[142] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_145 
+ bl[143] br[143] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_146 
+ bl[144] br[144] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_147 
+ bl[145] br[145] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_148 
+ bl[146] br[146] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_149 
+ bl[147] br[147] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_150 
+ bl[148] br[148] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_151 
+ bl[149] br[149] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_152 
+ bl[150] br[150] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_153 
+ bl[151] br[151] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_154 
+ bl[152] br[152] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_155 
+ bl[153] br[153] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_156 
+ bl[154] br[154] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_157 
+ bl[155] br[155] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_158 
+ bl[156] br[156] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_159 
+ bl[157] br[157] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_160 
+ bl[158] br[158] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_161 
+ bl[159] br[159] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_162 
+ bl[160] br[160] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_163 
+ bl[161] br[161] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_164 
+ bl[162] br[162] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_165 
+ bl[163] br[163] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_166 
+ bl[164] br[164] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_167 
+ bl[165] br[165] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_168 
+ bl[166] br[166] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_169 
+ bl[167] br[167] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_170 
+ bl[168] br[168] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_171 
+ bl[169] br[169] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_172 
+ bl[170] br[170] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_173 
+ bl[171] br[171] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_174 
+ bl[172] br[172] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_175 
+ bl[173] br[173] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_176 
+ bl[174] br[174] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_177 
+ bl[175] br[175] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_178 
+ bl[176] br[176] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_179 
+ bl[177] br[177] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_180 
+ bl[178] br[178] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_181 
+ bl[179] br[179] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_182 
+ bl[180] br[180] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_183 
+ bl[181] br[181] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_184 
+ bl[182] br[182] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_185 
+ bl[183] br[183] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_186 
+ bl[184] br[184] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_187 
+ bl[185] br[185] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_188 
+ bl[186] br[186] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_189 
+ bl[187] br[187] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_190 
+ bl[188] br[188] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_191 
+ bl[189] br[189] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_192 
+ bl[190] br[190] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_193 
+ bl[191] br[191] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_194 
+ bl[192] br[192] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_195 
+ bl[193] br[193] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_196 
+ bl[194] br[194] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_197 
+ bl[195] br[195] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_198 
+ bl[196] br[196] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_199 
+ bl[197] br[197] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_200 
+ bl[198] br[198] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_201 
+ bl[199] br[199] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_202 
+ bl[200] br[200] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_203 
+ bl[201] br[201] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_204 
+ bl[202] br[202] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_205 
+ bl[203] br[203] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_206 
+ bl[204] br[204] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_207 
+ bl[205] br[205] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_208 
+ bl[206] br[206] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_209 
+ bl[207] br[207] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_210 
+ bl[208] br[208] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_211 
+ bl[209] br[209] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_212 
+ bl[210] br[210] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_213 
+ bl[211] br[211] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_214 
+ bl[212] br[212] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_215 
+ bl[213] br[213] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_216 
+ bl[214] br[214] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_217 
+ bl[215] br[215] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_218 
+ bl[216] br[216] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_219 
+ bl[217] br[217] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_220 
+ bl[218] br[218] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_221 
+ bl[219] br[219] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_222 
+ bl[220] br[220] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_223 
+ bl[221] br[221] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_224 
+ bl[222] br[222] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_225 
+ bl[223] br[223] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_226 
+ bl[224] br[224] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_227 
+ bl[225] br[225] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_228 
+ bl[226] br[226] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_229 
+ bl[227] br[227] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_230 
+ bl[228] br[228] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_231 
+ bl[229] br[229] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_232 
+ bl[230] br[230] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_233 
+ bl[231] br[231] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_234 
+ bl[232] br[232] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_235 
+ bl[233] br[233] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_236 
+ bl[234] br[234] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_237 
+ bl[235] br[235] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_238 
+ bl[236] br[236] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_239 
+ bl[237] br[237] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_240 
+ bl[238] br[238] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_241 
+ bl[239] br[239] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_242 
+ bl[240] br[240] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_243 
+ bl[241] br[241] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_244 
+ bl[242] br[242] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_245 
+ bl[243] br[243] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_246 
+ bl[244] br[244] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_247 
+ bl[245] br[245] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_248 
+ bl[246] br[246] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_249 
+ bl[247] br[247] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_250 
+ bl[248] br[248] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_251 
+ bl[249] br[249] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_252 
+ bl[250] br[250] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_253 
+ bl[251] br[251] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_254 
+ bl[252] br[252] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_255 
+ bl[253] br[253] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_256 
+ bl[254] br[254] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_257 
+ bl[255] br[255] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_258 
+ vdd vdd vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_259 
+ vdd vdd vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_0 
+ vdd vdd vss vdd vpb vnb wl[88] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_90_1 
+ rbl rbr vss vdd vpb vnb wl[88] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_90_2 
+ bl[0] br[0] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_3 
+ bl[1] br[1] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_4 
+ bl[2] br[2] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_5 
+ bl[3] br[3] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_6 
+ bl[4] br[4] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_7 
+ bl[5] br[5] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_8 
+ bl[6] br[6] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_9 
+ bl[7] br[7] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_10 
+ bl[8] br[8] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_11 
+ bl[9] br[9] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_12 
+ bl[10] br[10] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_13 
+ bl[11] br[11] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_14 
+ bl[12] br[12] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_15 
+ bl[13] br[13] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_16 
+ bl[14] br[14] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_17 
+ bl[15] br[15] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_18 
+ bl[16] br[16] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_19 
+ bl[17] br[17] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_20 
+ bl[18] br[18] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_21 
+ bl[19] br[19] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_22 
+ bl[20] br[20] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_23 
+ bl[21] br[21] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_24 
+ bl[22] br[22] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_25 
+ bl[23] br[23] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_26 
+ bl[24] br[24] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_27 
+ bl[25] br[25] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_28 
+ bl[26] br[26] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_29 
+ bl[27] br[27] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_30 
+ bl[28] br[28] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_31 
+ bl[29] br[29] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_32 
+ bl[30] br[30] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_33 
+ bl[31] br[31] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_34 
+ bl[32] br[32] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_35 
+ bl[33] br[33] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_36 
+ bl[34] br[34] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_37 
+ bl[35] br[35] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_38 
+ bl[36] br[36] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_39 
+ bl[37] br[37] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_40 
+ bl[38] br[38] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_41 
+ bl[39] br[39] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_42 
+ bl[40] br[40] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_43 
+ bl[41] br[41] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_44 
+ bl[42] br[42] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_45 
+ bl[43] br[43] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_46 
+ bl[44] br[44] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_47 
+ bl[45] br[45] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_48 
+ bl[46] br[46] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_49 
+ bl[47] br[47] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_50 
+ bl[48] br[48] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_51 
+ bl[49] br[49] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_52 
+ bl[50] br[50] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_53 
+ bl[51] br[51] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_54 
+ bl[52] br[52] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_55 
+ bl[53] br[53] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_56 
+ bl[54] br[54] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_57 
+ bl[55] br[55] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_58 
+ bl[56] br[56] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_59 
+ bl[57] br[57] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_60 
+ bl[58] br[58] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_61 
+ bl[59] br[59] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_62 
+ bl[60] br[60] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_63 
+ bl[61] br[61] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_64 
+ bl[62] br[62] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_65 
+ bl[63] br[63] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_66 
+ bl[64] br[64] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_67 
+ bl[65] br[65] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_68 
+ bl[66] br[66] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_69 
+ bl[67] br[67] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_70 
+ bl[68] br[68] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_71 
+ bl[69] br[69] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_72 
+ bl[70] br[70] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_73 
+ bl[71] br[71] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_74 
+ bl[72] br[72] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_75 
+ bl[73] br[73] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_76 
+ bl[74] br[74] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_77 
+ bl[75] br[75] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_78 
+ bl[76] br[76] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_79 
+ bl[77] br[77] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_80 
+ bl[78] br[78] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_81 
+ bl[79] br[79] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_82 
+ bl[80] br[80] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_83 
+ bl[81] br[81] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_84 
+ bl[82] br[82] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_85 
+ bl[83] br[83] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_86 
+ bl[84] br[84] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_87 
+ bl[85] br[85] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_88 
+ bl[86] br[86] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_89 
+ bl[87] br[87] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_90 
+ bl[88] br[88] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_91 
+ bl[89] br[89] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_92 
+ bl[90] br[90] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_93 
+ bl[91] br[91] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_94 
+ bl[92] br[92] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_95 
+ bl[93] br[93] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_96 
+ bl[94] br[94] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_97 
+ bl[95] br[95] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_98 
+ bl[96] br[96] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_99 
+ bl[97] br[97] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_100 
+ bl[98] br[98] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_101 
+ bl[99] br[99] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_102 
+ bl[100] br[100] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_103 
+ bl[101] br[101] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_104 
+ bl[102] br[102] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_105 
+ bl[103] br[103] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_106 
+ bl[104] br[104] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_107 
+ bl[105] br[105] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_108 
+ bl[106] br[106] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_109 
+ bl[107] br[107] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_110 
+ bl[108] br[108] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_111 
+ bl[109] br[109] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_112 
+ bl[110] br[110] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_113 
+ bl[111] br[111] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_114 
+ bl[112] br[112] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_115 
+ bl[113] br[113] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_116 
+ bl[114] br[114] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_117 
+ bl[115] br[115] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_118 
+ bl[116] br[116] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_119 
+ bl[117] br[117] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_120 
+ bl[118] br[118] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_121 
+ bl[119] br[119] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_122 
+ bl[120] br[120] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_123 
+ bl[121] br[121] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_124 
+ bl[122] br[122] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_125 
+ bl[123] br[123] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_126 
+ bl[124] br[124] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_127 
+ bl[125] br[125] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_128 
+ bl[126] br[126] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_129 
+ bl[127] br[127] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_130 
+ bl[128] br[128] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_131 
+ bl[129] br[129] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_132 
+ bl[130] br[130] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_133 
+ bl[131] br[131] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_134 
+ bl[132] br[132] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_135 
+ bl[133] br[133] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_136 
+ bl[134] br[134] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_137 
+ bl[135] br[135] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_138 
+ bl[136] br[136] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_139 
+ bl[137] br[137] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_140 
+ bl[138] br[138] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_141 
+ bl[139] br[139] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_142 
+ bl[140] br[140] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_143 
+ bl[141] br[141] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_144 
+ bl[142] br[142] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_145 
+ bl[143] br[143] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_146 
+ bl[144] br[144] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_147 
+ bl[145] br[145] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_148 
+ bl[146] br[146] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_149 
+ bl[147] br[147] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_150 
+ bl[148] br[148] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_151 
+ bl[149] br[149] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_152 
+ bl[150] br[150] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_153 
+ bl[151] br[151] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_154 
+ bl[152] br[152] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_155 
+ bl[153] br[153] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_156 
+ bl[154] br[154] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_157 
+ bl[155] br[155] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_158 
+ bl[156] br[156] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_159 
+ bl[157] br[157] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_160 
+ bl[158] br[158] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_161 
+ bl[159] br[159] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_162 
+ bl[160] br[160] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_163 
+ bl[161] br[161] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_164 
+ bl[162] br[162] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_165 
+ bl[163] br[163] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_166 
+ bl[164] br[164] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_167 
+ bl[165] br[165] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_168 
+ bl[166] br[166] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_169 
+ bl[167] br[167] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_170 
+ bl[168] br[168] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_171 
+ bl[169] br[169] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_172 
+ bl[170] br[170] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_173 
+ bl[171] br[171] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_174 
+ bl[172] br[172] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_175 
+ bl[173] br[173] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_176 
+ bl[174] br[174] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_177 
+ bl[175] br[175] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_178 
+ bl[176] br[176] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_179 
+ bl[177] br[177] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_180 
+ bl[178] br[178] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_181 
+ bl[179] br[179] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_182 
+ bl[180] br[180] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_183 
+ bl[181] br[181] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_184 
+ bl[182] br[182] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_185 
+ bl[183] br[183] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_186 
+ bl[184] br[184] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_187 
+ bl[185] br[185] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_188 
+ bl[186] br[186] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_189 
+ bl[187] br[187] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_190 
+ bl[188] br[188] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_191 
+ bl[189] br[189] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_192 
+ bl[190] br[190] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_193 
+ bl[191] br[191] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_194 
+ bl[192] br[192] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_195 
+ bl[193] br[193] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_196 
+ bl[194] br[194] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_197 
+ bl[195] br[195] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_198 
+ bl[196] br[196] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_199 
+ bl[197] br[197] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_200 
+ bl[198] br[198] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_201 
+ bl[199] br[199] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_202 
+ bl[200] br[200] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_203 
+ bl[201] br[201] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_204 
+ bl[202] br[202] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_205 
+ bl[203] br[203] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_206 
+ bl[204] br[204] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_207 
+ bl[205] br[205] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_208 
+ bl[206] br[206] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_209 
+ bl[207] br[207] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_210 
+ bl[208] br[208] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_211 
+ bl[209] br[209] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_212 
+ bl[210] br[210] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_213 
+ bl[211] br[211] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_214 
+ bl[212] br[212] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_215 
+ bl[213] br[213] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_216 
+ bl[214] br[214] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_217 
+ bl[215] br[215] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_218 
+ bl[216] br[216] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_219 
+ bl[217] br[217] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_220 
+ bl[218] br[218] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_221 
+ bl[219] br[219] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_222 
+ bl[220] br[220] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_223 
+ bl[221] br[221] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_224 
+ bl[222] br[222] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_225 
+ bl[223] br[223] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_226 
+ bl[224] br[224] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_227 
+ bl[225] br[225] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_228 
+ bl[226] br[226] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_229 
+ bl[227] br[227] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_230 
+ bl[228] br[228] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_231 
+ bl[229] br[229] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_232 
+ bl[230] br[230] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_233 
+ bl[231] br[231] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_234 
+ bl[232] br[232] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_235 
+ bl[233] br[233] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_236 
+ bl[234] br[234] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_237 
+ bl[235] br[235] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_238 
+ bl[236] br[236] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_239 
+ bl[237] br[237] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_240 
+ bl[238] br[238] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_241 
+ bl[239] br[239] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_242 
+ bl[240] br[240] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_243 
+ bl[241] br[241] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_244 
+ bl[242] br[242] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_245 
+ bl[243] br[243] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_246 
+ bl[244] br[244] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_247 
+ bl[245] br[245] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_248 
+ bl[246] br[246] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_249 
+ bl[247] br[247] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_250 
+ bl[248] br[248] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_251 
+ bl[249] br[249] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_252 
+ bl[250] br[250] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_253 
+ bl[251] br[251] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_254 
+ bl[252] br[252] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_255 
+ bl[253] br[253] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_256 
+ bl[254] br[254] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_257 
+ bl[255] br[255] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_258 
+ vdd vdd vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_259 
+ vdd vdd vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_0 
+ vdd vdd vss vdd vpb vnb wl[89] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_91_1 
+ rbl rbr vss vdd vpb vnb wl[89] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_91_2 
+ bl[0] br[0] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_3 
+ bl[1] br[1] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_4 
+ bl[2] br[2] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_5 
+ bl[3] br[3] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_6 
+ bl[4] br[4] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_7 
+ bl[5] br[5] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_8 
+ bl[6] br[6] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_9 
+ bl[7] br[7] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_10 
+ bl[8] br[8] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_11 
+ bl[9] br[9] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_12 
+ bl[10] br[10] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_13 
+ bl[11] br[11] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_14 
+ bl[12] br[12] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_15 
+ bl[13] br[13] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_16 
+ bl[14] br[14] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_17 
+ bl[15] br[15] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_18 
+ bl[16] br[16] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_19 
+ bl[17] br[17] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_20 
+ bl[18] br[18] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_21 
+ bl[19] br[19] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_22 
+ bl[20] br[20] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_23 
+ bl[21] br[21] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_24 
+ bl[22] br[22] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_25 
+ bl[23] br[23] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_26 
+ bl[24] br[24] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_27 
+ bl[25] br[25] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_28 
+ bl[26] br[26] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_29 
+ bl[27] br[27] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_30 
+ bl[28] br[28] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_31 
+ bl[29] br[29] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_32 
+ bl[30] br[30] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_33 
+ bl[31] br[31] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_34 
+ bl[32] br[32] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_35 
+ bl[33] br[33] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_36 
+ bl[34] br[34] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_37 
+ bl[35] br[35] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_38 
+ bl[36] br[36] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_39 
+ bl[37] br[37] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_40 
+ bl[38] br[38] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_41 
+ bl[39] br[39] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_42 
+ bl[40] br[40] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_43 
+ bl[41] br[41] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_44 
+ bl[42] br[42] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_45 
+ bl[43] br[43] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_46 
+ bl[44] br[44] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_47 
+ bl[45] br[45] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_48 
+ bl[46] br[46] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_49 
+ bl[47] br[47] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_50 
+ bl[48] br[48] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_51 
+ bl[49] br[49] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_52 
+ bl[50] br[50] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_53 
+ bl[51] br[51] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_54 
+ bl[52] br[52] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_55 
+ bl[53] br[53] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_56 
+ bl[54] br[54] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_57 
+ bl[55] br[55] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_58 
+ bl[56] br[56] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_59 
+ bl[57] br[57] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_60 
+ bl[58] br[58] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_61 
+ bl[59] br[59] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_62 
+ bl[60] br[60] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_63 
+ bl[61] br[61] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_64 
+ bl[62] br[62] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_65 
+ bl[63] br[63] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_66 
+ bl[64] br[64] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_67 
+ bl[65] br[65] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_68 
+ bl[66] br[66] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_69 
+ bl[67] br[67] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_70 
+ bl[68] br[68] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_71 
+ bl[69] br[69] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_72 
+ bl[70] br[70] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_73 
+ bl[71] br[71] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_74 
+ bl[72] br[72] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_75 
+ bl[73] br[73] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_76 
+ bl[74] br[74] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_77 
+ bl[75] br[75] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_78 
+ bl[76] br[76] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_79 
+ bl[77] br[77] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_80 
+ bl[78] br[78] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_81 
+ bl[79] br[79] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_82 
+ bl[80] br[80] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_83 
+ bl[81] br[81] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_84 
+ bl[82] br[82] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_85 
+ bl[83] br[83] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_86 
+ bl[84] br[84] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_87 
+ bl[85] br[85] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_88 
+ bl[86] br[86] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_89 
+ bl[87] br[87] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_90 
+ bl[88] br[88] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_91 
+ bl[89] br[89] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_92 
+ bl[90] br[90] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_93 
+ bl[91] br[91] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_94 
+ bl[92] br[92] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_95 
+ bl[93] br[93] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_96 
+ bl[94] br[94] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_97 
+ bl[95] br[95] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_98 
+ bl[96] br[96] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_99 
+ bl[97] br[97] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_100 
+ bl[98] br[98] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_101 
+ bl[99] br[99] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_102 
+ bl[100] br[100] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_103 
+ bl[101] br[101] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_104 
+ bl[102] br[102] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_105 
+ bl[103] br[103] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_106 
+ bl[104] br[104] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_107 
+ bl[105] br[105] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_108 
+ bl[106] br[106] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_109 
+ bl[107] br[107] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_110 
+ bl[108] br[108] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_111 
+ bl[109] br[109] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_112 
+ bl[110] br[110] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_113 
+ bl[111] br[111] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_114 
+ bl[112] br[112] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_115 
+ bl[113] br[113] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_116 
+ bl[114] br[114] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_117 
+ bl[115] br[115] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_118 
+ bl[116] br[116] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_119 
+ bl[117] br[117] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_120 
+ bl[118] br[118] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_121 
+ bl[119] br[119] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_122 
+ bl[120] br[120] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_123 
+ bl[121] br[121] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_124 
+ bl[122] br[122] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_125 
+ bl[123] br[123] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_126 
+ bl[124] br[124] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_127 
+ bl[125] br[125] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_128 
+ bl[126] br[126] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_129 
+ bl[127] br[127] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_130 
+ bl[128] br[128] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_131 
+ bl[129] br[129] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_132 
+ bl[130] br[130] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_133 
+ bl[131] br[131] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_134 
+ bl[132] br[132] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_135 
+ bl[133] br[133] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_136 
+ bl[134] br[134] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_137 
+ bl[135] br[135] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_138 
+ bl[136] br[136] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_139 
+ bl[137] br[137] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_140 
+ bl[138] br[138] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_141 
+ bl[139] br[139] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_142 
+ bl[140] br[140] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_143 
+ bl[141] br[141] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_144 
+ bl[142] br[142] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_145 
+ bl[143] br[143] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_146 
+ bl[144] br[144] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_147 
+ bl[145] br[145] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_148 
+ bl[146] br[146] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_149 
+ bl[147] br[147] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_150 
+ bl[148] br[148] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_151 
+ bl[149] br[149] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_152 
+ bl[150] br[150] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_153 
+ bl[151] br[151] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_154 
+ bl[152] br[152] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_155 
+ bl[153] br[153] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_156 
+ bl[154] br[154] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_157 
+ bl[155] br[155] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_158 
+ bl[156] br[156] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_159 
+ bl[157] br[157] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_160 
+ bl[158] br[158] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_161 
+ bl[159] br[159] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_162 
+ bl[160] br[160] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_163 
+ bl[161] br[161] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_164 
+ bl[162] br[162] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_165 
+ bl[163] br[163] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_166 
+ bl[164] br[164] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_167 
+ bl[165] br[165] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_168 
+ bl[166] br[166] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_169 
+ bl[167] br[167] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_170 
+ bl[168] br[168] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_171 
+ bl[169] br[169] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_172 
+ bl[170] br[170] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_173 
+ bl[171] br[171] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_174 
+ bl[172] br[172] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_175 
+ bl[173] br[173] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_176 
+ bl[174] br[174] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_177 
+ bl[175] br[175] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_178 
+ bl[176] br[176] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_179 
+ bl[177] br[177] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_180 
+ bl[178] br[178] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_181 
+ bl[179] br[179] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_182 
+ bl[180] br[180] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_183 
+ bl[181] br[181] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_184 
+ bl[182] br[182] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_185 
+ bl[183] br[183] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_186 
+ bl[184] br[184] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_187 
+ bl[185] br[185] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_188 
+ bl[186] br[186] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_189 
+ bl[187] br[187] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_190 
+ bl[188] br[188] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_191 
+ bl[189] br[189] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_192 
+ bl[190] br[190] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_193 
+ bl[191] br[191] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_194 
+ bl[192] br[192] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_195 
+ bl[193] br[193] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_196 
+ bl[194] br[194] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_197 
+ bl[195] br[195] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_198 
+ bl[196] br[196] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_199 
+ bl[197] br[197] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_200 
+ bl[198] br[198] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_201 
+ bl[199] br[199] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_202 
+ bl[200] br[200] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_203 
+ bl[201] br[201] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_204 
+ bl[202] br[202] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_205 
+ bl[203] br[203] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_206 
+ bl[204] br[204] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_207 
+ bl[205] br[205] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_208 
+ bl[206] br[206] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_209 
+ bl[207] br[207] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_210 
+ bl[208] br[208] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_211 
+ bl[209] br[209] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_212 
+ bl[210] br[210] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_213 
+ bl[211] br[211] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_214 
+ bl[212] br[212] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_215 
+ bl[213] br[213] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_216 
+ bl[214] br[214] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_217 
+ bl[215] br[215] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_218 
+ bl[216] br[216] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_219 
+ bl[217] br[217] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_220 
+ bl[218] br[218] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_221 
+ bl[219] br[219] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_222 
+ bl[220] br[220] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_223 
+ bl[221] br[221] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_224 
+ bl[222] br[222] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_225 
+ bl[223] br[223] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_226 
+ bl[224] br[224] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_227 
+ bl[225] br[225] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_228 
+ bl[226] br[226] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_229 
+ bl[227] br[227] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_230 
+ bl[228] br[228] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_231 
+ bl[229] br[229] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_232 
+ bl[230] br[230] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_233 
+ bl[231] br[231] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_234 
+ bl[232] br[232] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_235 
+ bl[233] br[233] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_236 
+ bl[234] br[234] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_237 
+ bl[235] br[235] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_238 
+ bl[236] br[236] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_239 
+ bl[237] br[237] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_240 
+ bl[238] br[238] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_241 
+ bl[239] br[239] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_242 
+ bl[240] br[240] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_243 
+ bl[241] br[241] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_244 
+ bl[242] br[242] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_245 
+ bl[243] br[243] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_246 
+ bl[244] br[244] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_247 
+ bl[245] br[245] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_248 
+ bl[246] br[246] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_249 
+ bl[247] br[247] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_250 
+ bl[248] br[248] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_251 
+ bl[249] br[249] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_252 
+ bl[250] br[250] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_253 
+ bl[251] br[251] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_254 
+ bl[252] br[252] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_255 
+ bl[253] br[253] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_256 
+ bl[254] br[254] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_257 
+ bl[255] br[255] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_258 
+ vdd vdd vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_259 
+ vdd vdd vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_0 
+ vdd vdd vss vdd vpb vnb wl[90] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_92_1 
+ rbl rbr vss vdd vpb vnb wl[90] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_92_2 
+ bl[0] br[0] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_3 
+ bl[1] br[1] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_4 
+ bl[2] br[2] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_5 
+ bl[3] br[3] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_6 
+ bl[4] br[4] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_7 
+ bl[5] br[5] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_8 
+ bl[6] br[6] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_9 
+ bl[7] br[7] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_10 
+ bl[8] br[8] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_11 
+ bl[9] br[9] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_12 
+ bl[10] br[10] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_13 
+ bl[11] br[11] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_14 
+ bl[12] br[12] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_15 
+ bl[13] br[13] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_16 
+ bl[14] br[14] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_17 
+ bl[15] br[15] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_18 
+ bl[16] br[16] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_19 
+ bl[17] br[17] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_20 
+ bl[18] br[18] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_21 
+ bl[19] br[19] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_22 
+ bl[20] br[20] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_23 
+ bl[21] br[21] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_24 
+ bl[22] br[22] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_25 
+ bl[23] br[23] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_26 
+ bl[24] br[24] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_27 
+ bl[25] br[25] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_28 
+ bl[26] br[26] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_29 
+ bl[27] br[27] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_30 
+ bl[28] br[28] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_31 
+ bl[29] br[29] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_32 
+ bl[30] br[30] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_33 
+ bl[31] br[31] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_34 
+ bl[32] br[32] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_35 
+ bl[33] br[33] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_36 
+ bl[34] br[34] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_37 
+ bl[35] br[35] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_38 
+ bl[36] br[36] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_39 
+ bl[37] br[37] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_40 
+ bl[38] br[38] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_41 
+ bl[39] br[39] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_42 
+ bl[40] br[40] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_43 
+ bl[41] br[41] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_44 
+ bl[42] br[42] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_45 
+ bl[43] br[43] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_46 
+ bl[44] br[44] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_47 
+ bl[45] br[45] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_48 
+ bl[46] br[46] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_49 
+ bl[47] br[47] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_50 
+ bl[48] br[48] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_51 
+ bl[49] br[49] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_52 
+ bl[50] br[50] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_53 
+ bl[51] br[51] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_54 
+ bl[52] br[52] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_55 
+ bl[53] br[53] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_56 
+ bl[54] br[54] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_57 
+ bl[55] br[55] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_58 
+ bl[56] br[56] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_59 
+ bl[57] br[57] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_60 
+ bl[58] br[58] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_61 
+ bl[59] br[59] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_62 
+ bl[60] br[60] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_63 
+ bl[61] br[61] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_64 
+ bl[62] br[62] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_65 
+ bl[63] br[63] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_66 
+ bl[64] br[64] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_67 
+ bl[65] br[65] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_68 
+ bl[66] br[66] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_69 
+ bl[67] br[67] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_70 
+ bl[68] br[68] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_71 
+ bl[69] br[69] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_72 
+ bl[70] br[70] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_73 
+ bl[71] br[71] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_74 
+ bl[72] br[72] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_75 
+ bl[73] br[73] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_76 
+ bl[74] br[74] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_77 
+ bl[75] br[75] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_78 
+ bl[76] br[76] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_79 
+ bl[77] br[77] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_80 
+ bl[78] br[78] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_81 
+ bl[79] br[79] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_82 
+ bl[80] br[80] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_83 
+ bl[81] br[81] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_84 
+ bl[82] br[82] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_85 
+ bl[83] br[83] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_86 
+ bl[84] br[84] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_87 
+ bl[85] br[85] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_88 
+ bl[86] br[86] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_89 
+ bl[87] br[87] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_90 
+ bl[88] br[88] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_91 
+ bl[89] br[89] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_92 
+ bl[90] br[90] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_93 
+ bl[91] br[91] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_94 
+ bl[92] br[92] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_95 
+ bl[93] br[93] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_96 
+ bl[94] br[94] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_97 
+ bl[95] br[95] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_98 
+ bl[96] br[96] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_99 
+ bl[97] br[97] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_100 
+ bl[98] br[98] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_101 
+ bl[99] br[99] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_102 
+ bl[100] br[100] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_103 
+ bl[101] br[101] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_104 
+ bl[102] br[102] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_105 
+ bl[103] br[103] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_106 
+ bl[104] br[104] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_107 
+ bl[105] br[105] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_108 
+ bl[106] br[106] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_109 
+ bl[107] br[107] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_110 
+ bl[108] br[108] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_111 
+ bl[109] br[109] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_112 
+ bl[110] br[110] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_113 
+ bl[111] br[111] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_114 
+ bl[112] br[112] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_115 
+ bl[113] br[113] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_116 
+ bl[114] br[114] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_117 
+ bl[115] br[115] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_118 
+ bl[116] br[116] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_119 
+ bl[117] br[117] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_120 
+ bl[118] br[118] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_121 
+ bl[119] br[119] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_122 
+ bl[120] br[120] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_123 
+ bl[121] br[121] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_124 
+ bl[122] br[122] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_125 
+ bl[123] br[123] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_126 
+ bl[124] br[124] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_127 
+ bl[125] br[125] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_128 
+ bl[126] br[126] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_129 
+ bl[127] br[127] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_130 
+ bl[128] br[128] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_131 
+ bl[129] br[129] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_132 
+ bl[130] br[130] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_133 
+ bl[131] br[131] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_134 
+ bl[132] br[132] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_135 
+ bl[133] br[133] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_136 
+ bl[134] br[134] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_137 
+ bl[135] br[135] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_138 
+ bl[136] br[136] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_139 
+ bl[137] br[137] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_140 
+ bl[138] br[138] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_141 
+ bl[139] br[139] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_142 
+ bl[140] br[140] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_143 
+ bl[141] br[141] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_144 
+ bl[142] br[142] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_145 
+ bl[143] br[143] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_146 
+ bl[144] br[144] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_147 
+ bl[145] br[145] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_148 
+ bl[146] br[146] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_149 
+ bl[147] br[147] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_150 
+ bl[148] br[148] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_151 
+ bl[149] br[149] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_152 
+ bl[150] br[150] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_153 
+ bl[151] br[151] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_154 
+ bl[152] br[152] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_155 
+ bl[153] br[153] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_156 
+ bl[154] br[154] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_157 
+ bl[155] br[155] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_158 
+ bl[156] br[156] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_159 
+ bl[157] br[157] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_160 
+ bl[158] br[158] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_161 
+ bl[159] br[159] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_162 
+ bl[160] br[160] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_163 
+ bl[161] br[161] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_164 
+ bl[162] br[162] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_165 
+ bl[163] br[163] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_166 
+ bl[164] br[164] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_167 
+ bl[165] br[165] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_168 
+ bl[166] br[166] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_169 
+ bl[167] br[167] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_170 
+ bl[168] br[168] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_171 
+ bl[169] br[169] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_172 
+ bl[170] br[170] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_173 
+ bl[171] br[171] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_174 
+ bl[172] br[172] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_175 
+ bl[173] br[173] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_176 
+ bl[174] br[174] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_177 
+ bl[175] br[175] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_178 
+ bl[176] br[176] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_179 
+ bl[177] br[177] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_180 
+ bl[178] br[178] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_181 
+ bl[179] br[179] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_182 
+ bl[180] br[180] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_183 
+ bl[181] br[181] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_184 
+ bl[182] br[182] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_185 
+ bl[183] br[183] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_186 
+ bl[184] br[184] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_187 
+ bl[185] br[185] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_188 
+ bl[186] br[186] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_189 
+ bl[187] br[187] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_190 
+ bl[188] br[188] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_191 
+ bl[189] br[189] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_192 
+ bl[190] br[190] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_193 
+ bl[191] br[191] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_194 
+ bl[192] br[192] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_195 
+ bl[193] br[193] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_196 
+ bl[194] br[194] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_197 
+ bl[195] br[195] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_198 
+ bl[196] br[196] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_199 
+ bl[197] br[197] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_200 
+ bl[198] br[198] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_201 
+ bl[199] br[199] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_202 
+ bl[200] br[200] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_203 
+ bl[201] br[201] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_204 
+ bl[202] br[202] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_205 
+ bl[203] br[203] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_206 
+ bl[204] br[204] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_207 
+ bl[205] br[205] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_208 
+ bl[206] br[206] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_209 
+ bl[207] br[207] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_210 
+ bl[208] br[208] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_211 
+ bl[209] br[209] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_212 
+ bl[210] br[210] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_213 
+ bl[211] br[211] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_214 
+ bl[212] br[212] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_215 
+ bl[213] br[213] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_216 
+ bl[214] br[214] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_217 
+ bl[215] br[215] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_218 
+ bl[216] br[216] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_219 
+ bl[217] br[217] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_220 
+ bl[218] br[218] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_221 
+ bl[219] br[219] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_222 
+ bl[220] br[220] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_223 
+ bl[221] br[221] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_224 
+ bl[222] br[222] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_225 
+ bl[223] br[223] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_226 
+ bl[224] br[224] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_227 
+ bl[225] br[225] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_228 
+ bl[226] br[226] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_229 
+ bl[227] br[227] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_230 
+ bl[228] br[228] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_231 
+ bl[229] br[229] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_232 
+ bl[230] br[230] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_233 
+ bl[231] br[231] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_234 
+ bl[232] br[232] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_235 
+ bl[233] br[233] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_236 
+ bl[234] br[234] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_237 
+ bl[235] br[235] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_238 
+ bl[236] br[236] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_239 
+ bl[237] br[237] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_240 
+ bl[238] br[238] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_241 
+ bl[239] br[239] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_242 
+ bl[240] br[240] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_243 
+ bl[241] br[241] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_244 
+ bl[242] br[242] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_245 
+ bl[243] br[243] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_246 
+ bl[244] br[244] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_247 
+ bl[245] br[245] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_248 
+ bl[246] br[246] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_249 
+ bl[247] br[247] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_250 
+ bl[248] br[248] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_251 
+ bl[249] br[249] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_252 
+ bl[250] br[250] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_253 
+ bl[251] br[251] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_254 
+ bl[252] br[252] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_255 
+ bl[253] br[253] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_256 
+ bl[254] br[254] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_257 
+ bl[255] br[255] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_258 
+ vdd vdd vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_259 
+ vdd vdd vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_0 
+ vdd vdd vss vdd vpb vnb wl[91] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_93_1 
+ rbl rbr vss vdd vpb vnb wl[91] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_93_2 
+ bl[0] br[0] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_3 
+ bl[1] br[1] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_4 
+ bl[2] br[2] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_5 
+ bl[3] br[3] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_6 
+ bl[4] br[4] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_7 
+ bl[5] br[5] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_8 
+ bl[6] br[6] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_9 
+ bl[7] br[7] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_10 
+ bl[8] br[8] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_11 
+ bl[9] br[9] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_12 
+ bl[10] br[10] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_13 
+ bl[11] br[11] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_14 
+ bl[12] br[12] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_15 
+ bl[13] br[13] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_16 
+ bl[14] br[14] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_17 
+ bl[15] br[15] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_18 
+ bl[16] br[16] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_19 
+ bl[17] br[17] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_20 
+ bl[18] br[18] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_21 
+ bl[19] br[19] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_22 
+ bl[20] br[20] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_23 
+ bl[21] br[21] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_24 
+ bl[22] br[22] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_25 
+ bl[23] br[23] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_26 
+ bl[24] br[24] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_27 
+ bl[25] br[25] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_28 
+ bl[26] br[26] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_29 
+ bl[27] br[27] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_30 
+ bl[28] br[28] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_31 
+ bl[29] br[29] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_32 
+ bl[30] br[30] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_33 
+ bl[31] br[31] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_34 
+ bl[32] br[32] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_35 
+ bl[33] br[33] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_36 
+ bl[34] br[34] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_37 
+ bl[35] br[35] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_38 
+ bl[36] br[36] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_39 
+ bl[37] br[37] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_40 
+ bl[38] br[38] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_41 
+ bl[39] br[39] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_42 
+ bl[40] br[40] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_43 
+ bl[41] br[41] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_44 
+ bl[42] br[42] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_45 
+ bl[43] br[43] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_46 
+ bl[44] br[44] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_47 
+ bl[45] br[45] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_48 
+ bl[46] br[46] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_49 
+ bl[47] br[47] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_50 
+ bl[48] br[48] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_51 
+ bl[49] br[49] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_52 
+ bl[50] br[50] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_53 
+ bl[51] br[51] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_54 
+ bl[52] br[52] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_55 
+ bl[53] br[53] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_56 
+ bl[54] br[54] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_57 
+ bl[55] br[55] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_58 
+ bl[56] br[56] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_59 
+ bl[57] br[57] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_60 
+ bl[58] br[58] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_61 
+ bl[59] br[59] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_62 
+ bl[60] br[60] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_63 
+ bl[61] br[61] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_64 
+ bl[62] br[62] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_65 
+ bl[63] br[63] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_66 
+ bl[64] br[64] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_67 
+ bl[65] br[65] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_68 
+ bl[66] br[66] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_69 
+ bl[67] br[67] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_70 
+ bl[68] br[68] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_71 
+ bl[69] br[69] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_72 
+ bl[70] br[70] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_73 
+ bl[71] br[71] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_74 
+ bl[72] br[72] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_75 
+ bl[73] br[73] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_76 
+ bl[74] br[74] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_77 
+ bl[75] br[75] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_78 
+ bl[76] br[76] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_79 
+ bl[77] br[77] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_80 
+ bl[78] br[78] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_81 
+ bl[79] br[79] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_82 
+ bl[80] br[80] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_83 
+ bl[81] br[81] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_84 
+ bl[82] br[82] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_85 
+ bl[83] br[83] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_86 
+ bl[84] br[84] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_87 
+ bl[85] br[85] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_88 
+ bl[86] br[86] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_89 
+ bl[87] br[87] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_90 
+ bl[88] br[88] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_91 
+ bl[89] br[89] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_92 
+ bl[90] br[90] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_93 
+ bl[91] br[91] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_94 
+ bl[92] br[92] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_95 
+ bl[93] br[93] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_96 
+ bl[94] br[94] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_97 
+ bl[95] br[95] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_98 
+ bl[96] br[96] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_99 
+ bl[97] br[97] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_100 
+ bl[98] br[98] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_101 
+ bl[99] br[99] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_102 
+ bl[100] br[100] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_103 
+ bl[101] br[101] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_104 
+ bl[102] br[102] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_105 
+ bl[103] br[103] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_106 
+ bl[104] br[104] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_107 
+ bl[105] br[105] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_108 
+ bl[106] br[106] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_109 
+ bl[107] br[107] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_110 
+ bl[108] br[108] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_111 
+ bl[109] br[109] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_112 
+ bl[110] br[110] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_113 
+ bl[111] br[111] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_114 
+ bl[112] br[112] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_115 
+ bl[113] br[113] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_116 
+ bl[114] br[114] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_117 
+ bl[115] br[115] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_118 
+ bl[116] br[116] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_119 
+ bl[117] br[117] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_120 
+ bl[118] br[118] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_121 
+ bl[119] br[119] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_122 
+ bl[120] br[120] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_123 
+ bl[121] br[121] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_124 
+ bl[122] br[122] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_125 
+ bl[123] br[123] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_126 
+ bl[124] br[124] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_127 
+ bl[125] br[125] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_128 
+ bl[126] br[126] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_129 
+ bl[127] br[127] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_130 
+ bl[128] br[128] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_131 
+ bl[129] br[129] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_132 
+ bl[130] br[130] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_133 
+ bl[131] br[131] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_134 
+ bl[132] br[132] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_135 
+ bl[133] br[133] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_136 
+ bl[134] br[134] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_137 
+ bl[135] br[135] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_138 
+ bl[136] br[136] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_139 
+ bl[137] br[137] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_140 
+ bl[138] br[138] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_141 
+ bl[139] br[139] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_142 
+ bl[140] br[140] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_143 
+ bl[141] br[141] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_144 
+ bl[142] br[142] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_145 
+ bl[143] br[143] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_146 
+ bl[144] br[144] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_147 
+ bl[145] br[145] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_148 
+ bl[146] br[146] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_149 
+ bl[147] br[147] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_150 
+ bl[148] br[148] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_151 
+ bl[149] br[149] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_152 
+ bl[150] br[150] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_153 
+ bl[151] br[151] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_154 
+ bl[152] br[152] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_155 
+ bl[153] br[153] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_156 
+ bl[154] br[154] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_157 
+ bl[155] br[155] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_158 
+ bl[156] br[156] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_159 
+ bl[157] br[157] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_160 
+ bl[158] br[158] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_161 
+ bl[159] br[159] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_162 
+ bl[160] br[160] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_163 
+ bl[161] br[161] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_164 
+ bl[162] br[162] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_165 
+ bl[163] br[163] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_166 
+ bl[164] br[164] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_167 
+ bl[165] br[165] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_168 
+ bl[166] br[166] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_169 
+ bl[167] br[167] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_170 
+ bl[168] br[168] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_171 
+ bl[169] br[169] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_172 
+ bl[170] br[170] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_173 
+ bl[171] br[171] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_174 
+ bl[172] br[172] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_175 
+ bl[173] br[173] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_176 
+ bl[174] br[174] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_177 
+ bl[175] br[175] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_178 
+ bl[176] br[176] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_179 
+ bl[177] br[177] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_180 
+ bl[178] br[178] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_181 
+ bl[179] br[179] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_182 
+ bl[180] br[180] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_183 
+ bl[181] br[181] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_184 
+ bl[182] br[182] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_185 
+ bl[183] br[183] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_186 
+ bl[184] br[184] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_187 
+ bl[185] br[185] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_188 
+ bl[186] br[186] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_189 
+ bl[187] br[187] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_190 
+ bl[188] br[188] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_191 
+ bl[189] br[189] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_192 
+ bl[190] br[190] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_193 
+ bl[191] br[191] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_194 
+ bl[192] br[192] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_195 
+ bl[193] br[193] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_196 
+ bl[194] br[194] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_197 
+ bl[195] br[195] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_198 
+ bl[196] br[196] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_199 
+ bl[197] br[197] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_200 
+ bl[198] br[198] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_201 
+ bl[199] br[199] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_202 
+ bl[200] br[200] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_203 
+ bl[201] br[201] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_204 
+ bl[202] br[202] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_205 
+ bl[203] br[203] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_206 
+ bl[204] br[204] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_207 
+ bl[205] br[205] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_208 
+ bl[206] br[206] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_209 
+ bl[207] br[207] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_210 
+ bl[208] br[208] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_211 
+ bl[209] br[209] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_212 
+ bl[210] br[210] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_213 
+ bl[211] br[211] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_214 
+ bl[212] br[212] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_215 
+ bl[213] br[213] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_216 
+ bl[214] br[214] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_217 
+ bl[215] br[215] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_218 
+ bl[216] br[216] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_219 
+ bl[217] br[217] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_220 
+ bl[218] br[218] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_221 
+ bl[219] br[219] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_222 
+ bl[220] br[220] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_223 
+ bl[221] br[221] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_224 
+ bl[222] br[222] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_225 
+ bl[223] br[223] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_226 
+ bl[224] br[224] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_227 
+ bl[225] br[225] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_228 
+ bl[226] br[226] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_229 
+ bl[227] br[227] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_230 
+ bl[228] br[228] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_231 
+ bl[229] br[229] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_232 
+ bl[230] br[230] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_233 
+ bl[231] br[231] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_234 
+ bl[232] br[232] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_235 
+ bl[233] br[233] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_236 
+ bl[234] br[234] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_237 
+ bl[235] br[235] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_238 
+ bl[236] br[236] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_239 
+ bl[237] br[237] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_240 
+ bl[238] br[238] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_241 
+ bl[239] br[239] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_242 
+ bl[240] br[240] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_243 
+ bl[241] br[241] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_244 
+ bl[242] br[242] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_245 
+ bl[243] br[243] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_246 
+ bl[244] br[244] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_247 
+ bl[245] br[245] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_248 
+ bl[246] br[246] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_249 
+ bl[247] br[247] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_250 
+ bl[248] br[248] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_251 
+ bl[249] br[249] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_252 
+ bl[250] br[250] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_253 
+ bl[251] br[251] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_254 
+ bl[252] br[252] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_255 
+ bl[253] br[253] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_256 
+ bl[254] br[254] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_257 
+ bl[255] br[255] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_258 
+ vdd vdd vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_259 
+ vdd vdd vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_0 
+ vdd vdd vss vdd vpb vnb wl[92] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_94_1 
+ rbl rbr vss vdd vpb vnb wl[92] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_94_2 
+ bl[0] br[0] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_3 
+ bl[1] br[1] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_4 
+ bl[2] br[2] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_5 
+ bl[3] br[3] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_6 
+ bl[4] br[4] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_7 
+ bl[5] br[5] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_8 
+ bl[6] br[6] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_9 
+ bl[7] br[7] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_10 
+ bl[8] br[8] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_11 
+ bl[9] br[9] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_12 
+ bl[10] br[10] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_13 
+ bl[11] br[11] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_14 
+ bl[12] br[12] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_15 
+ bl[13] br[13] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_16 
+ bl[14] br[14] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_17 
+ bl[15] br[15] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_18 
+ bl[16] br[16] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_19 
+ bl[17] br[17] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_20 
+ bl[18] br[18] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_21 
+ bl[19] br[19] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_22 
+ bl[20] br[20] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_23 
+ bl[21] br[21] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_24 
+ bl[22] br[22] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_25 
+ bl[23] br[23] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_26 
+ bl[24] br[24] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_27 
+ bl[25] br[25] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_28 
+ bl[26] br[26] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_29 
+ bl[27] br[27] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_30 
+ bl[28] br[28] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_31 
+ bl[29] br[29] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_32 
+ bl[30] br[30] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_33 
+ bl[31] br[31] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_34 
+ bl[32] br[32] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_35 
+ bl[33] br[33] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_36 
+ bl[34] br[34] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_37 
+ bl[35] br[35] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_38 
+ bl[36] br[36] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_39 
+ bl[37] br[37] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_40 
+ bl[38] br[38] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_41 
+ bl[39] br[39] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_42 
+ bl[40] br[40] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_43 
+ bl[41] br[41] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_44 
+ bl[42] br[42] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_45 
+ bl[43] br[43] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_46 
+ bl[44] br[44] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_47 
+ bl[45] br[45] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_48 
+ bl[46] br[46] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_49 
+ bl[47] br[47] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_50 
+ bl[48] br[48] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_51 
+ bl[49] br[49] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_52 
+ bl[50] br[50] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_53 
+ bl[51] br[51] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_54 
+ bl[52] br[52] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_55 
+ bl[53] br[53] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_56 
+ bl[54] br[54] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_57 
+ bl[55] br[55] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_58 
+ bl[56] br[56] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_59 
+ bl[57] br[57] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_60 
+ bl[58] br[58] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_61 
+ bl[59] br[59] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_62 
+ bl[60] br[60] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_63 
+ bl[61] br[61] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_64 
+ bl[62] br[62] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_65 
+ bl[63] br[63] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_66 
+ bl[64] br[64] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_67 
+ bl[65] br[65] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_68 
+ bl[66] br[66] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_69 
+ bl[67] br[67] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_70 
+ bl[68] br[68] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_71 
+ bl[69] br[69] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_72 
+ bl[70] br[70] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_73 
+ bl[71] br[71] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_74 
+ bl[72] br[72] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_75 
+ bl[73] br[73] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_76 
+ bl[74] br[74] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_77 
+ bl[75] br[75] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_78 
+ bl[76] br[76] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_79 
+ bl[77] br[77] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_80 
+ bl[78] br[78] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_81 
+ bl[79] br[79] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_82 
+ bl[80] br[80] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_83 
+ bl[81] br[81] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_84 
+ bl[82] br[82] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_85 
+ bl[83] br[83] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_86 
+ bl[84] br[84] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_87 
+ bl[85] br[85] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_88 
+ bl[86] br[86] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_89 
+ bl[87] br[87] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_90 
+ bl[88] br[88] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_91 
+ bl[89] br[89] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_92 
+ bl[90] br[90] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_93 
+ bl[91] br[91] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_94 
+ bl[92] br[92] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_95 
+ bl[93] br[93] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_96 
+ bl[94] br[94] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_97 
+ bl[95] br[95] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_98 
+ bl[96] br[96] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_99 
+ bl[97] br[97] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_100 
+ bl[98] br[98] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_101 
+ bl[99] br[99] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_102 
+ bl[100] br[100] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_103 
+ bl[101] br[101] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_104 
+ bl[102] br[102] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_105 
+ bl[103] br[103] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_106 
+ bl[104] br[104] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_107 
+ bl[105] br[105] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_108 
+ bl[106] br[106] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_109 
+ bl[107] br[107] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_110 
+ bl[108] br[108] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_111 
+ bl[109] br[109] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_112 
+ bl[110] br[110] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_113 
+ bl[111] br[111] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_114 
+ bl[112] br[112] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_115 
+ bl[113] br[113] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_116 
+ bl[114] br[114] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_117 
+ bl[115] br[115] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_118 
+ bl[116] br[116] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_119 
+ bl[117] br[117] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_120 
+ bl[118] br[118] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_121 
+ bl[119] br[119] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_122 
+ bl[120] br[120] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_123 
+ bl[121] br[121] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_124 
+ bl[122] br[122] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_125 
+ bl[123] br[123] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_126 
+ bl[124] br[124] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_127 
+ bl[125] br[125] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_128 
+ bl[126] br[126] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_129 
+ bl[127] br[127] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_130 
+ bl[128] br[128] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_131 
+ bl[129] br[129] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_132 
+ bl[130] br[130] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_133 
+ bl[131] br[131] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_134 
+ bl[132] br[132] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_135 
+ bl[133] br[133] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_136 
+ bl[134] br[134] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_137 
+ bl[135] br[135] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_138 
+ bl[136] br[136] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_139 
+ bl[137] br[137] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_140 
+ bl[138] br[138] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_141 
+ bl[139] br[139] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_142 
+ bl[140] br[140] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_143 
+ bl[141] br[141] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_144 
+ bl[142] br[142] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_145 
+ bl[143] br[143] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_146 
+ bl[144] br[144] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_147 
+ bl[145] br[145] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_148 
+ bl[146] br[146] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_149 
+ bl[147] br[147] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_150 
+ bl[148] br[148] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_151 
+ bl[149] br[149] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_152 
+ bl[150] br[150] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_153 
+ bl[151] br[151] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_154 
+ bl[152] br[152] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_155 
+ bl[153] br[153] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_156 
+ bl[154] br[154] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_157 
+ bl[155] br[155] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_158 
+ bl[156] br[156] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_159 
+ bl[157] br[157] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_160 
+ bl[158] br[158] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_161 
+ bl[159] br[159] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_162 
+ bl[160] br[160] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_163 
+ bl[161] br[161] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_164 
+ bl[162] br[162] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_165 
+ bl[163] br[163] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_166 
+ bl[164] br[164] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_167 
+ bl[165] br[165] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_168 
+ bl[166] br[166] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_169 
+ bl[167] br[167] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_170 
+ bl[168] br[168] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_171 
+ bl[169] br[169] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_172 
+ bl[170] br[170] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_173 
+ bl[171] br[171] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_174 
+ bl[172] br[172] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_175 
+ bl[173] br[173] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_176 
+ bl[174] br[174] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_177 
+ bl[175] br[175] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_178 
+ bl[176] br[176] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_179 
+ bl[177] br[177] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_180 
+ bl[178] br[178] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_181 
+ bl[179] br[179] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_182 
+ bl[180] br[180] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_183 
+ bl[181] br[181] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_184 
+ bl[182] br[182] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_185 
+ bl[183] br[183] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_186 
+ bl[184] br[184] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_187 
+ bl[185] br[185] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_188 
+ bl[186] br[186] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_189 
+ bl[187] br[187] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_190 
+ bl[188] br[188] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_191 
+ bl[189] br[189] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_192 
+ bl[190] br[190] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_193 
+ bl[191] br[191] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_194 
+ bl[192] br[192] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_195 
+ bl[193] br[193] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_196 
+ bl[194] br[194] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_197 
+ bl[195] br[195] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_198 
+ bl[196] br[196] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_199 
+ bl[197] br[197] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_200 
+ bl[198] br[198] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_201 
+ bl[199] br[199] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_202 
+ bl[200] br[200] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_203 
+ bl[201] br[201] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_204 
+ bl[202] br[202] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_205 
+ bl[203] br[203] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_206 
+ bl[204] br[204] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_207 
+ bl[205] br[205] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_208 
+ bl[206] br[206] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_209 
+ bl[207] br[207] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_210 
+ bl[208] br[208] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_211 
+ bl[209] br[209] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_212 
+ bl[210] br[210] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_213 
+ bl[211] br[211] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_214 
+ bl[212] br[212] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_215 
+ bl[213] br[213] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_216 
+ bl[214] br[214] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_217 
+ bl[215] br[215] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_218 
+ bl[216] br[216] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_219 
+ bl[217] br[217] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_220 
+ bl[218] br[218] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_221 
+ bl[219] br[219] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_222 
+ bl[220] br[220] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_223 
+ bl[221] br[221] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_224 
+ bl[222] br[222] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_225 
+ bl[223] br[223] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_226 
+ bl[224] br[224] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_227 
+ bl[225] br[225] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_228 
+ bl[226] br[226] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_229 
+ bl[227] br[227] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_230 
+ bl[228] br[228] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_231 
+ bl[229] br[229] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_232 
+ bl[230] br[230] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_233 
+ bl[231] br[231] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_234 
+ bl[232] br[232] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_235 
+ bl[233] br[233] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_236 
+ bl[234] br[234] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_237 
+ bl[235] br[235] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_238 
+ bl[236] br[236] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_239 
+ bl[237] br[237] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_240 
+ bl[238] br[238] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_241 
+ bl[239] br[239] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_242 
+ bl[240] br[240] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_243 
+ bl[241] br[241] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_244 
+ bl[242] br[242] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_245 
+ bl[243] br[243] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_246 
+ bl[244] br[244] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_247 
+ bl[245] br[245] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_248 
+ bl[246] br[246] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_249 
+ bl[247] br[247] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_250 
+ bl[248] br[248] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_251 
+ bl[249] br[249] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_252 
+ bl[250] br[250] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_253 
+ bl[251] br[251] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_254 
+ bl[252] br[252] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_255 
+ bl[253] br[253] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_256 
+ bl[254] br[254] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_257 
+ bl[255] br[255] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_258 
+ vdd vdd vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_259 
+ vdd vdd vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_0 
+ vdd vdd vss vdd vpb vnb wl[93] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_95_1 
+ rbl rbr vss vdd vpb vnb wl[93] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_95_2 
+ bl[0] br[0] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_3 
+ bl[1] br[1] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_4 
+ bl[2] br[2] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_5 
+ bl[3] br[3] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_6 
+ bl[4] br[4] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_7 
+ bl[5] br[5] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_8 
+ bl[6] br[6] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_9 
+ bl[7] br[7] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_10 
+ bl[8] br[8] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_11 
+ bl[9] br[9] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_12 
+ bl[10] br[10] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_13 
+ bl[11] br[11] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_14 
+ bl[12] br[12] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_15 
+ bl[13] br[13] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_16 
+ bl[14] br[14] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_17 
+ bl[15] br[15] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_18 
+ bl[16] br[16] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_19 
+ bl[17] br[17] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_20 
+ bl[18] br[18] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_21 
+ bl[19] br[19] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_22 
+ bl[20] br[20] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_23 
+ bl[21] br[21] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_24 
+ bl[22] br[22] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_25 
+ bl[23] br[23] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_26 
+ bl[24] br[24] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_27 
+ bl[25] br[25] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_28 
+ bl[26] br[26] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_29 
+ bl[27] br[27] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_30 
+ bl[28] br[28] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_31 
+ bl[29] br[29] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_32 
+ bl[30] br[30] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_33 
+ bl[31] br[31] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_34 
+ bl[32] br[32] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_35 
+ bl[33] br[33] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_36 
+ bl[34] br[34] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_37 
+ bl[35] br[35] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_38 
+ bl[36] br[36] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_39 
+ bl[37] br[37] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_40 
+ bl[38] br[38] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_41 
+ bl[39] br[39] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_42 
+ bl[40] br[40] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_43 
+ bl[41] br[41] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_44 
+ bl[42] br[42] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_45 
+ bl[43] br[43] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_46 
+ bl[44] br[44] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_47 
+ bl[45] br[45] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_48 
+ bl[46] br[46] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_49 
+ bl[47] br[47] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_50 
+ bl[48] br[48] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_51 
+ bl[49] br[49] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_52 
+ bl[50] br[50] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_53 
+ bl[51] br[51] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_54 
+ bl[52] br[52] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_55 
+ bl[53] br[53] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_56 
+ bl[54] br[54] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_57 
+ bl[55] br[55] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_58 
+ bl[56] br[56] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_59 
+ bl[57] br[57] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_60 
+ bl[58] br[58] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_61 
+ bl[59] br[59] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_62 
+ bl[60] br[60] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_63 
+ bl[61] br[61] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_64 
+ bl[62] br[62] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_65 
+ bl[63] br[63] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_66 
+ bl[64] br[64] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_67 
+ bl[65] br[65] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_68 
+ bl[66] br[66] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_69 
+ bl[67] br[67] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_70 
+ bl[68] br[68] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_71 
+ bl[69] br[69] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_72 
+ bl[70] br[70] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_73 
+ bl[71] br[71] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_74 
+ bl[72] br[72] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_75 
+ bl[73] br[73] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_76 
+ bl[74] br[74] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_77 
+ bl[75] br[75] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_78 
+ bl[76] br[76] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_79 
+ bl[77] br[77] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_80 
+ bl[78] br[78] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_81 
+ bl[79] br[79] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_82 
+ bl[80] br[80] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_83 
+ bl[81] br[81] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_84 
+ bl[82] br[82] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_85 
+ bl[83] br[83] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_86 
+ bl[84] br[84] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_87 
+ bl[85] br[85] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_88 
+ bl[86] br[86] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_89 
+ bl[87] br[87] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_90 
+ bl[88] br[88] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_91 
+ bl[89] br[89] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_92 
+ bl[90] br[90] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_93 
+ bl[91] br[91] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_94 
+ bl[92] br[92] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_95 
+ bl[93] br[93] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_96 
+ bl[94] br[94] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_97 
+ bl[95] br[95] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_98 
+ bl[96] br[96] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_99 
+ bl[97] br[97] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_100 
+ bl[98] br[98] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_101 
+ bl[99] br[99] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_102 
+ bl[100] br[100] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_103 
+ bl[101] br[101] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_104 
+ bl[102] br[102] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_105 
+ bl[103] br[103] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_106 
+ bl[104] br[104] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_107 
+ bl[105] br[105] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_108 
+ bl[106] br[106] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_109 
+ bl[107] br[107] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_110 
+ bl[108] br[108] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_111 
+ bl[109] br[109] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_112 
+ bl[110] br[110] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_113 
+ bl[111] br[111] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_114 
+ bl[112] br[112] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_115 
+ bl[113] br[113] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_116 
+ bl[114] br[114] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_117 
+ bl[115] br[115] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_118 
+ bl[116] br[116] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_119 
+ bl[117] br[117] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_120 
+ bl[118] br[118] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_121 
+ bl[119] br[119] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_122 
+ bl[120] br[120] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_123 
+ bl[121] br[121] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_124 
+ bl[122] br[122] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_125 
+ bl[123] br[123] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_126 
+ bl[124] br[124] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_127 
+ bl[125] br[125] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_128 
+ bl[126] br[126] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_129 
+ bl[127] br[127] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_130 
+ bl[128] br[128] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_131 
+ bl[129] br[129] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_132 
+ bl[130] br[130] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_133 
+ bl[131] br[131] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_134 
+ bl[132] br[132] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_135 
+ bl[133] br[133] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_136 
+ bl[134] br[134] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_137 
+ bl[135] br[135] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_138 
+ bl[136] br[136] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_139 
+ bl[137] br[137] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_140 
+ bl[138] br[138] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_141 
+ bl[139] br[139] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_142 
+ bl[140] br[140] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_143 
+ bl[141] br[141] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_144 
+ bl[142] br[142] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_145 
+ bl[143] br[143] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_146 
+ bl[144] br[144] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_147 
+ bl[145] br[145] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_148 
+ bl[146] br[146] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_149 
+ bl[147] br[147] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_150 
+ bl[148] br[148] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_151 
+ bl[149] br[149] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_152 
+ bl[150] br[150] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_153 
+ bl[151] br[151] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_154 
+ bl[152] br[152] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_155 
+ bl[153] br[153] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_156 
+ bl[154] br[154] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_157 
+ bl[155] br[155] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_158 
+ bl[156] br[156] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_159 
+ bl[157] br[157] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_160 
+ bl[158] br[158] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_161 
+ bl[159] br[159] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_162 
+ bl[160] br[160] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_163 
+ bl[161] br[161] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_164 
+ bl[162] br[162] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_165 
+ bl[163] br[163] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_166 
+ bl[164] br[164] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_167 
+ bl[165] br[165] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_168 
+ bl[166] br[166] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_169 
+ bl[167] br[167] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_170 
+ bl[168] br[168] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_171 
+ bl[169] br[169] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_172 
+ bl[170] br[170] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_173 
+ bl[171] br[171] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_174 
+ bl[172] br[172] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_175 
+ bl[173] br[173] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_176 
+ bl[174] br[174] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_177 
+ bl[175] br[175] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_178 
+ bl[176] br[176] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_179 
+ bl[177] br[177] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_180 
+ bl[178] br[178] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_181 
+ bl[179] br[179] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_182 
+ bl[180] br[180] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_183 
+ bl[181] br[181] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_184 
+ bl[182] br[182] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_185 
+ bl[183] br[183] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_186 
+ bl[184] br[184] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_187 
+ bl[185] br[185] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_188 
+ bl[186] br[186] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_189 
+ bl[187] br[187] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_190 
+ bl[188] br[188] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_191 
+ bl[189] br[189] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_192 
+ bl[190] br[190] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_193 
+ bl[191] br[191] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_194 
+ bl[192] br[192] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_195 
+ bl[193] br[193] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_196 
+ bl[194] br[194] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_197 
+ bl[195] br[195] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_198 
+ bl[196] br[196] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_199 
+ bl[197] br[197] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_200 
+ bl[198] br[198] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_201 
+ bl[199] br[199] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_202 
+ bl[200] br[200] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_203 
+ bl[201] br[201] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_204 
+ bl[202] br[202] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_205 
+ bl[203] br[203] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_206 
+ bl[204] br[204] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_207 
+ bl[205] br[205] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_208 
+ bl[206] br[206] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_209 
+ bl[207] br[207] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_210 
+ bl[208] br[208] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_211 
+ bl[209] br[209] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_212 
+ bl[210] br[210] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_213 
+ bl[211] br[211] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_214 
+ bl[212] br[212] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_215 
+ bl[213] br[213] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_216 
+ bl[214] br[214] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_217 
+ bl[215] br[215] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_218 
+ bl[216] br[216] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_219 
+ bl[217] br[217] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_220 
+ bl[218] br[218] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_221 
+ bl[219] br[219] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_222 
+ bl[220] br[220] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_223 
+ bl[221] br[221] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_224 
+ bl[222] br[222] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_225 
+ bl[223] br[223] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_226 
+ bl[224] br[224] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_227 
+ bl[225] br[225] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_228 
+ bl[226] br[226] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_229 
+ bl[227] br[227] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_230 
+ bl[228] br[228] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_231 
+ bl[229] br[229] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_232 
+ bl[230] br[230] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_233 
+ bl[231] br[231] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_234 
+ bl[232] br[232] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_235 
+ bl[233] br[233] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_236 
+ bl[234] br[234] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_237 
+ bl[235] br[235] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_238 
+ bl[236] br[236] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_239 
+ bl[237] br[237] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_240 
+ bl[238] br[238] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_241 
+ bl[239] br[239] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_242 
+ bl[240] br[240] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_243 
+ bl[241] br[241] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_244 
+ bl[242] br[242] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_245 
+ bl[243] br[243] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_246 
+ bl[244] br[244] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_247 
+ bl[245] br[245] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_248 
+ bl[246] br[246] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_249 
+ bl[247] br[247] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_250 
+ bl[248] br[248] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_251 
+ bl[249] br[249] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_252 
+ bl[250] br[250] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_253 
+ bl[251] br[251] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_254 
+ bl[252] br[252] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_255 
+ bl[253] br[253] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_256 
+ bl[254] br[254] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_257 
+ bl[255] br[255] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_258 
+ vdd vdd vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_259 
+ vdd vdd vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_0 
+ vdd vdd vss vdd vpb vnb wl[94] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_96_1 
+ rbl rbr vss vdd vpb vnb wl[94] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_96_2 
+ bl[0] br[0] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_3 
+ bl[1] br[1] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_4 
+ bl[2] br[2] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_5 
+ bl[3] br[3] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_6 
+ bl[4] br[4] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_7 
+ bl[5] br[5] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_8 
+ bl[6] br[6] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_9 
+ bl[7] br[7] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_10 
+ bl[8] br[8] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_11 
+ bl[9] br[9] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_12 
+ bl[10] br[10] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_13 
+ bl[11] br[11] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_14 
+ bl[12] br[12] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_15 
+ bl[13] br[13] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_16 
+ bl[14] br[14] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_17 
+ bl[15] br[15] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_18 
+ bl[16] br[16] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_19 
+ bl[17] br[17] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_20 
+ bl[18] br[18] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_21 
+ bl[19] br[19] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_22 
+ bl[20] br[20] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_23 
+ bl[21] br[21] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_24 
+ bl[22] br[22] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_25 
+ bl[23] br[23] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_26 
+ bl[24] br[24] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_27 
+ bl[25] br[25] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_28 
+ bl[26] br[26] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_29 
+ bl[27] br[27] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_30 
+ bl[28] br[28] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_31 
+ bl[29] br[29] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_32 
+ bl[30] br[30] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_33 
+ bl[31] br[31] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_34 
+ bl[32] br[32] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_35 
+ bl[33] br[33] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_36 
+ bl[34] br[34] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_37 
+ bl[35] br[35] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_38 
+ bl[36] br[36] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_39 
+ bl[37] br[37] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_40 
+ bl[38] br[38] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_41 
+ bl[39] br[39] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_42 
+ bl[40] br[40] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_43 
+ bl[41] br[41] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_44 
+ bl[42] br[42] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_45 
+ bl[43] br[43] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_46 
+ bl[44] br[44] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_47 
+ bl[45] br[45] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_48 
+ bl[46] br[46] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_49 
+ bl[47] br[47] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_50 
+ bl[48] br[48] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_51 
+ bl[49] br[49] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_52 
+ bl[50] br[50] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_53 
+ bl[51] br[51] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_54 
+ bl[52] br[52] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_55 
+ bl[53] br[53] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_56 
+ bl[54] br[54] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_57 
+ bl[55] br[55] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_58 
+ bl[56] br[56] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_59 
+ bl[57] br[57] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_60 
+ bl[58] br[58] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_61 
+ bl[59] br[59] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_62 
+ bl[60] br[60] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_63 
+ bl[61] br[61] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_64 
+ bl[62] br[62] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_65 
+ bl[63] br[63] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_66 
+ bl[64] br[64] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_67 
+ bl[65] br[65] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_68 
+ bl[66] br[66] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_69 
+ bl[67] br[67] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_70 
+ bl[68] br[68] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_71 
+ bl[69] br[69] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_72 
+ bl[70] br[70] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_73 
+ bl[71] br[71] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_74 
+ bl[72] br[72] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_75 
+ bl[73] br[73] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_76 
+ bl[74] br[74] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_77 
+ bl[75] br[75] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_78 
+ bl[76] br[76] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_79 
+ bl[77] br[77] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_80 
+ bl[78] br[78] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_81 
+ bl[79] br[79] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_82 
+ bl[80] br[80] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_83 
+ bl[81] br[81] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_84 
+ bl[82] br[82] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_85 
+ bl[83] br[83] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_86 
+ bl[84] br[84] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_87 
+ bl[85] br[85] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_88 
+ bl[86] br[86] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_89 
+ bl[87] br[87] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_90 
+ bl[88] br[88] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_91 
+ bl[89] br[89] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_92 
+ bl[90] br[90] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_93 
+ bl[91] br[91] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_94 
+ bl[92] br[92] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_95 
+ bl[93] br[93] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_96 
+ bl[94] br[94] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_97 
+ bl[95] br[95] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_98 
+ bl[96] br[96] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_99 
+ bl[97] br[97] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_100 
+ bl[98] br[98] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_101 
+ bl[99] br[99] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_102 
+ bl[100] br[100] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_103 
+ bl[101] br[101] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_104 
+ bl[102] br[102] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_105 
+ bl[103] br[103] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_106 
+ bl[104] br[104] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_107 
+ bl[105] br[105] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_108 
+ bl[106] br[106] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_109 
+ bl[107] br[107] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_110 
+ bl[108] br[108] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_111 
+ bl[109] br[109] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_112 
+ bl[110] br[110] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_113 
+ bl[111] br[111] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_114 
+ bl[112] br[112] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_115 
+ bl[113] br[113] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_116 
+ bl[114] br[114] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_117 
+ bl[115] br[115] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_118 
+ bl[116] br[116] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_119 
+ bl[117] br[117] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_120 
+ bl[118] br[118] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_121 
+ bl[119] br[119] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_122 
+ bl[120] br[120] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_123 
+ bl[121] br[121] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_124 
+ bl[122] br[122] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_125 
+ bl[123] br[123] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_126 
+ bl[124] br[124] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_127 
+ bl[125] br[125] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_128 
+ bl[126] br[126] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_129 
+ bl[127] br[127] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_130 
+ bl[128] br[128] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_131 
+ bl[129] br[129] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_132 
+ bl[130] br[130] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_133 
+ bl[131] br[131] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_134 
+ bl[132] br[132] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_135 
+ bl[133] br[133] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_136 
+ bl[134] br[134] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_137 
+ bl[135] br[135] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_138 
+ bl[136] br[136] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_139 
+ bl[137] br[137] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_140 
+ bl[138] br[138] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_141 
+ bl[139] br[139] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_142 
+ bl[140] br[140] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_143 
+ bl[141] br[141] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_144 
+ bl[142] br[142] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_145 
+ bl[143] br[143] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_146 
+ bl[144] br[144] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_147 
+ bl[145] br[145] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_148 
+ bl[146] br[146] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_149 
+ bl[147] br[147] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_150 
+ bl[148] br[148] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_151 
+ bl[149] br[149] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_152 
+ bl[150] br[150] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_153 
+ bl[151] br[151] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_154 
+ bl[152] br[152] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_155 
+ bl[153] br[153] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_156 
+ bl[154] br[154] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_157 
+ bl[155] br[155] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_158 
+ bl[156] br[156] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_159 
+ bl[157] br[157] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_160 
+ bl[158] br[158] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_161 
+ bl[159] br[159] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_162 
+ bl[160] br[160] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_163 
+ bl[161] br[161] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_164 
+ bl[162] br[162] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_165 
+ bl[163] br[163] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_166 
+ bl[164] br[164] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_167 
+ bl[165] br[165] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_168 
+ bl[166] br[166] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_169 
+ bl[167] br[167] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_170 
+ bl[168] br[168] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_171 
+ bl[169] br[169] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_172 
+ bl[170] br[170] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_173 
+ bl[171] br[171] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_174 
+ bl[172] br[172] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_175 
+ bl[173] br[173] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_176 
+ bl[174] br[174] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_177 
+ bl[175] br[175] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_178 
+ bl[176] br[176] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_179 
+ bl[177] br[177] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_180 
+ bl[178] br[178] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_181 
+ bl[179] br[179] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_182 
+ bl[180] br[180] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_183 
+ bl[181] br[181] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_184 
+ bl[182] br[182] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_185 
+ bl[183] br[183] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_186 
+ bl[184] br[184] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_187 
+ bl[185] br[185] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_188 
+ bl[186] br[186] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_189 
+ bl[187] br[187] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_190 
+ bl[188] br[188] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_191 
+ bl[189] br[189] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_192 
+ bl[190] br[190] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_193 
+ bl[191] br[191] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_194 
+ bl[192] br[192] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_195 
+ bl[193] br[193] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_196 
+ bl[194] br[194] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_197 
+ bl[195] br[195] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_198 
+ bl[196] br[196] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_199 
+ bl[197] br[197] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_200 
+ bl[198] br[198] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_201 
+ bl[199] br[199] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_202 
+ bl[200] br[200] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_203 
+ bl[201] br[201] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_204 
+ bl[202] br[202] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_205 
+ bl[203] br[203] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_206 
+ bl[204] br[204] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_207 
+ bl[205] br[205] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_208 
+ bl[206] br[206] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_209 
+ bl[207] br[207] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_210 
+ bl[208] br[208] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_211 
+ bl[209] br[209] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_212 
+ bl[210] br[210] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_213 
+ bl[211] br[211] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_214 
+ bl[212] br[212] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_215 
+ bl[213] br[213] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_216 
+ bl[214] br[214] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_217 
+ bl[215] br[215] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_218 
+ bl[216] br[216] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_219 
+ bl[217] br[217] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_220 
+ bl[218] br[218] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_221 
+ bl[219] br[219] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_222 
+ bl[220] br[220] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_223 
+ bl[221] br[221] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_224 
+ bl[222] br[222] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_225 
+ bl[223] br[223] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_226 
+ bl[224] br[224] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_227 
+ bl[225] br[225] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_228 
+ bl[226] br[226] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_229 
+ bl[227] br[227] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_230 
+ bl[228] br[228] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_231 
+ bl[229] br[229] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_232 
+ bl[230] br[230] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_233 
+ bl[231] br[231] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_234 
+ bl[232] br[232] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_235 
+ bl[233] br[233] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_236 
+ bl[234] br[234] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_237 
+ bl[235] br[235] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_238 
+ bl[236] br[236] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_239 
+ bl[237] br[237] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_240 
+ bl[238] br[238] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_241 
+ bl[239] br[239] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_242 
+ bl[240] br[240] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_243 
+ bl[241] br[241] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_244 
+ bl[242] br[242] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_245 
+ bl[243] br[243] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_246 
+ bl[244] br[244] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_247 
+ bl[245] br[245] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_248 
+ bl[246] br[246] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_249 
+ bl[247] br[247] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_250 
+ bl[248] br[248] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_251 
+ bl[249] br[249] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_252 
+ bl[250] br[250] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_253 
+ bl[251] br[251] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_254 
+ bl[252] br[252] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_255 
+ bl[253] br[253] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_256 
+ bl[254] br[254] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_257 
+ bl[255] br[255] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_258 
+ vdd vdd vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_259 
+ vdd vdd vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_0 
+ vdd vdd vss vdd vpb vnb wl[95] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_97_1 
+ rbl rbr vss vdd vpb vnb wl[95] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_97_2 
+ bl[0] br[0] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_3 
+ bl[1] br[1] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_4 
+ bl[2] br[2] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_5 
+ bl[3] br[3] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_6 
+ bl[4] br[4] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_7 
+ bl[5] br[5] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_8 
+ bl[6] br[6] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_9 
+ bl[7] br[7] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_10 
+ bl[8] br[8] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_11 
+ bl[9] br[9] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_12 
+ bl[10] br[10] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_13 
+ bl[11] br[11] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_14 
+ bl[12] br[12] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_15 
+ bl[13] br[13] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_16 
+ bl[14] br[14] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_17 
+ bl[15] br[15] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_18 
+ bl[16] br[16] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_19 
+ bl[17] br[17] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_20 
+ bl[18] br[18] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_21 
+ bl[19] br[19] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_22 
+ bl[20] br[20] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_23 
+ bl[21] br[21] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_24 
+ bl[22] br[22] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_25 
+ bl[23] br[23] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_26 
+ bl[24] br[24] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_27 
+ bl[25] br[25] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_28 
+ bl[26] br[26] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_29 
+ bl[27] br[27] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_30 
+ bl[28] br[28] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_31 
+ bl[29] br[29] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_32 
+ bl[30] br[30] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_33 
+ bl[31] br[31] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_34 
+ bl[32] br[32] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_35 
+ bl[33] br[33] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_36 
+ bl[34] br[34] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_37 
+ bl[35] br[35] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_38 
+ bl[36] br[36] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_39 
+ bl[37] br[37] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_40 
+ bl[38] br[38] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_41 
+ bl[39] br[39] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_42 
+ bl[40] br[40] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_43 
+ bl[41] br[41] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_44 
+ bl[42] br[42] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_45 
+ bl[43] br[43] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_46 
+ bl[44] br[44] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_47 
+ bl[45] br[45] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_48 
+ bl[46] br[46] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_49 
+ bl[47] br[47] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_50 
+ bl[48] br[48] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_51 
+ bl[49] br[49] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_52 
+ bl[50] br[50] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_53 
+ bl[51] br[51] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_54 
+ bl[52] br[52] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_55 
+ bl[53] br[53] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_56 
+ bl[54] br[54] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_57 
+ bl[55] br[55] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_58 
+ bl[56] br[56] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_59 
+ bl[57] br[57] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_60 
+ bl[58] br[58] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_61 
+ bl[59] br[59] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_62 
+ bl[60] br[60] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_63 
+ bl[61] br[61] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_64 
+ bl[62] br[62] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_65 
+ bl[63] br[63] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_66 
+ bl[64] br[64] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_67 
+ bl[65] br[65] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_68 
+ bl[66] br[66] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_69 
+ bl[67] br[67] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_70 
+ bl[68] br[68] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_71 
+ bl[69] br[69] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_72 
+ bl[70] br[70] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_73 
+ bl[71] br[71] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_74 
+ bl[72] br[72] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_75 
+ bl[73] br[73] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_76 
+ bl[74] br[74] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_77 
+ bl[75] br[75] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_78 
+ bl[76] br[76] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_79 
+ bl[77] br[77] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_80 
+ bl[78] br[78] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_81 
+ bl[79] br[79] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_82 
+ bl[80] br[80] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_83 
+ bl[81] br[81] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_84 
+ bl[82] br[82] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_85 
+ bl[83] br[83] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_86 
+ bl[84] br[84] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_87 
+ bl[85] br[85] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_88 
+ bl[86] br[86] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_89 
+ bl[87] br[87] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_90 
+ bl[88] br[88] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_91 
+ bl[89] br[89] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_92 
+ bl[90] br[90] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_93 
+ bl[91] br[91] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_94 
+ bl[92] br[92] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_95 
+ bl[93] br[93] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_96 
+ bl[94] br[94] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_97 
+ bl[95] br[95] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_98 
+ bl[96] br[96] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_99 
+ bl[97] br[97] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_100 
+ bl[98] br[98] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_101 
+ bl[99] br[99] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_102 
+ bl[100] br[100] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_103 
+ bl[101] br[101] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_104 
+ bl[102] br[102] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_105 
+ bl[103] br[103] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_106 
+ bl[104] br[104] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_107 
+ bl[105] br[105] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_108 
+ bl[106] br[106] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_109 
+ bl[107] br[107] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_110 
+ bl[108] br[108] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_111 
+ bl[109] br[109] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_112 
+ bl[110] br[110] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_113 
+ bl[111] br[111] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_114 
+ bl[112] br[112] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_115 
+ bl[113] br[113] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_116 
+ bl[114] br[114] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_117 
+ bl[115] br[115] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_118 
+ bl[116] br[116] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_119 
+ bl[117] br[117] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_120 
+ bl[118] br[118] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_121 
+ bl[119] br[119] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_122 
+ bl[120] br[120] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_123 
+ bl[121] br[121] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_124 
+ bl[122] br[122] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_125 
+ bl[123] br[123] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_126 
+ bl[124] br[124] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_127 
+ bl[125] br[125] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_128 
+ bl[126] br[126] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_129 
+ bl[127] br[127] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_130 
+ bl[128] br[128] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_131 
+ bl[129] br[129] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_132 
+ bl[130] br[130] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_133 
+ bl[131] br[131] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_134 
+ bl[132] br[132] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_135 
+ bl[133] br[133] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_136 
+ bl[134] br[134] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_137 
+ bl[135] br[135] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_138 
+ bl[136] br[136] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_139 
+ bl[137] br[137] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_140 
+ bl[138] br[138] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_141 
+ bl[139] br[139] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_142 
+ bl[140] br[140] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_143 
+ bl[141] br[141] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_144 
+ bl[142] br[142] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_145 
+ bl[143] br[143] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_146 
+ bl[144] br[144] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_147 
+ bl[145] br[145] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_148 
+ bl[146] br[146] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_149 
+ bl[147] br[147] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_150 
+ bl[148] br[148] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_151 
+ bl[149] br[149] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_152 
+ bl[150] br[150] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_153 
+ bl[151] br[151] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_154 
+ bl[152] br[152] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_155 
+ bl[153] br[153] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_156 
+ bl[154] br[154] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_157 
+ bl[155] br[155] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_158 
+ bl[156] br[156] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_159 
+ bl[157] br[157] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_160 
+ bl[158] br[158] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_161 
+ bl[159] br[159] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_162 
+ bl[160] br[160] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_163 
+ bl[161] br[161] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_164 
+ bl[162] br[162] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_165 
+ bl[163] br[163] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_166 
+ bl[164] br[164] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_167 
+ bl[165] br[165] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_168 
+ bl[166] br[166] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_169 
+ bl[167] br[167] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_170 
+ bl[168] br[168] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_171 
+ bl[169] br[169] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_172 
+ bl[170] br[170] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_173 
+ bl[171] br[171] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_174 
+ bl[172] br[172] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_175 
+ bl[173] br[173] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_176 
+ bl[174] br[174] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_177 
+ bl[175] br[175] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_178 
+ bl[176] br[176] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_179 
+ bl[177] br[177] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_180 
+ bl[178] br[178] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_181 
+ bl[179] br[179] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_182 
+ bl[180] br[180] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_183 
+ bl[181] br[181] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_184 
+ bl[182] br[182] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_185 
+ bl[183] br[183] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_186 
+ bl[184] br[184] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_187 
+ bl[185] br[185] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_188 
+ bl[186] br[186] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_189 
+ bl[187] br[187] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_190 
+ bl[188] br[188] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_191 
+ bl[189] br[189] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_192 
+ bl[190] br[190] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_193 
+ bl[191] br[191] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_194 
+ bl[192] br[192] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_195 
+ bl[193] br[193] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_196 
+ bl[194] br[194] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_197 
+ bl[195] br[195] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_198 
+ bl[196] br[196] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_199 
+ bl[197] br[197] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_200 
+ bl[198] br[198] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_201 
+ bl[199] br[199] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_202 
+ bl[200] br[200] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_203 
+ bl[201] br[201] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_204 
+ bl[202] br[202] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_205 
+ bl[203] br[203] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_206 
+ bl[204] br[204] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_207 
+ bl[205] br[205] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_208 
+ bl[206] br[206] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_209 
+ bl[207] br[207] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_210 
+ bl[208] br[208] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_211 
+ bl[209] br[209] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_212 
+ bl[210] br[210] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_213 
+ bl[211] br[211] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_214 
+ bl[212] br[212] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_215 
+ bl[213] br[213] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_216 
+ bl[214] br[214] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_217 
+ bl[215] br[215] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_218 
+ bl[216] br[216] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_219 
+ bl[217] br[217] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_220 
+ bl[218] br[218] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_221 
+ bl[219] br[219] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_222 
+ bl[220] br[220] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_223 
+ bl[221] br[221] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_224 
+ bl[222] br[222] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_225 
+ bl[223] br[223] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_226 
+ bl[224] br[224] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_227 
+ bl[225] br[225] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_228 
+ bl[226] br[226] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_229 
+ bl[227] br[227] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_230 
+ bl[228] br[228] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_231 
+ bl[229] br[229] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_232 
+ bl[230] br[230] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_233 
+ bl[231] br[231] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_234 
+ bl[232] br[232] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_235 
+ bl[233] br[233] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_236 
+ bl[234] br[234] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_237 
+ bl[235] br[235] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_238 
+ bl[236] br[236] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_239 
+ bl[237] br[237] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_240 
+ bl[238] br[238] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_241 
+ bl[239] br[239] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_242 
+ bl[240] br[240] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_243 
+ bl[241] br[241] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_244 
+ bl[242] br[242] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_245 
+ bl[243] br[243] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_246 
+ bl[244] br[244] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_247 
+ bl[245] br[245] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_248 
+ bl[246] br[246] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_249 
+ bl[247] br[247] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_250 
+ bl[248] br[248] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_251 
+ bl[249] br[249] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_252 
+ bl[250] br[250] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_253 
+ bl[251] br[251] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_254 
+ bl[252] br[252] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_255 
+ bl[253] br[253] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_256 
+ bl[254] br[254] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_257 
+ bl[255] br[255] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_258 
+ vdd vdd vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_259 
+ vdd vdd vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_0 
+ vdd vdd vss vdd vpb vnb wl[96] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_98_1 
+ rbl rbr vss vdd vpb vnb wl[96] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_98_2 
+ bl[0] br[0] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_3 
+ bl[1] br[1] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_4 
+ bl[2] br[2] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_5 
+ bl[3] br[3] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_6 
+ bl[4] br[4] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_7 
+ bl[5] br[5] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_8 
+ bl[6] br[6] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_9 
+ bl[7] br[7] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_10 
+ bl[8] br[8] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_11 
+ bl[9] br[9] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_12 
+ bl[10] br[10] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_13 
+ bl[11] br[11] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_14 
+ bl[12] br[12] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_15 
+ bl[13] br[13] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_16 
+ bl[14] br[14] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_17 
+ bl[15] br[15] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_18 
+ bl[16] br[16] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_19 
+ bl[17] br[17] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_20 
+ bl[18] br[18] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_21 
+ bl[19] br[19] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_22 
+ bl[20] br[20] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_23 
+ bl[21] br[21] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_24 
+ bl[22] br[22] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_25 
+ bl[23] br[23] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_26 
+ bl[24] br[24] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_27 
+ bl[25] br[25] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_28 
+ bl[26] br[26] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_29 
+ bl[27] br[27] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_30 
+ bl[28] br[28] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_31 
+ bl[29] br[29] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_32 
+ bl[30] br[30] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_33 
+ bl[31] br[31] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_34 
+ bl[32] br[32] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_35 
+ bl[33] br[33] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_36 
+ bl[34] br[34] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_37 
+ bl[35] br[35] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_38 
+ bl[36] br[36] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_39 
+ bl[37] br[37] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_40 
+ bl[38] br[38] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_41 
+ bl[39] br[39] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_42 
+ bl[40] br[40] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_43 
+ bl[41] br[41] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_44 
+ bl[42] br[42] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_45 
+ bl[43] br[43] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_46 
+ bl[44] br[44] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_47 
+ bl[45] br[45] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_48 
+ bl[46] br[46] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_49 
+ bl[47] br[47] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_50 
+ bl[48] br[48] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_51 
+ bl[49] br[49] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_52 
+ bl[50] br[50] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_53 
+ bl[51] br[51] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_54 
+ bl[52] br[52] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_55 
+ bl[53] br[53] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_56 
+ bl[54] br[54] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_57 
+ bl[55] br[55] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_58 
+ bl[56] br[56] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_59 
+ bl[57] br[57] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_60 
+ bl[58] br[58] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_61 
+ bl[59] br[59] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_62 
+ bl[60] br[60] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_63 
+ bl[61] br[61] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_64 
+ bl[62] br[62] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_65 
+ bl[63] br[63] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_66 
+ bl[64] br[64] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_67 
+ bl[65] br[65] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_68 
+ bl[66] br[66] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_69 
+ bl[67] br[67] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_70 
+ bl[68] br[68] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_71 
+ bl[69] br[69] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_72 
+ bl[70] br[70] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_73 
+ bl[71] br[71] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_74 
+ bl[72] br[72] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_75 
+ bl[73] br[73] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_76 
+ bl[74] br[74] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_77 
+ bl[75] br[75] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_78 
+ bl[76] br[76] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_79 
+ bl[77] br[77] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_80 
+ bl[78] br[78] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_81 
+ bl[79] br[79] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_82 
+ bl[80] br[80] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_83 
+ bl[81] br[81] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_84 
+ bl[82] br[82] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_85 
+ bl[83] br[83] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_86 
+ bl[84] br[84] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_87 
+ bl[85] br[85] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_88 
+ bl[86] br[86] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_89 
+ bl[87] br[87] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_90 
+ bl[88] br[88] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_91 
+ bl[89] br[89] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_92 
+ bl[90] br[90] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_93 
+ bl[91] br[91] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_94 
+ bl[92] br[92] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_95 
+ bl[93] br[93] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_96 
+ bl[94] br[94] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_97 
+ bl[95] br[95] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_98 
+ bl[96] br[96] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_99 
+ bl[97] br[97] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_100 
+ bl[98] br[98] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_101 
+ bl[99] br[99] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_102 
+ bl[100] br[100] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_103 
+ bl[101] br[101] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_104 
+ bl[102] br[102] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_105 
+ bl[103] br[103] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_106 
+ bl[104] br[104] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_107 
+ bl[105] br[105] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_108 
+ bl[106] br[106] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_109 
+ bl[107] br[107] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_110 
+ bl[108] br[108] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_111 
+ bl[109] br[109] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_112 
+ bl[110] br[110] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_113 
+ bl[111] br[111] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_114 
+ bl[112] br[112] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_115 
+ bl[113] br[113] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_116 
+ bl[114] br[114] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_117 
+ bl[115] br[115] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_118 
+ bl[116] br[116] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_119 
+ bl[117] br[117] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_120 
+ bl[118] br[118] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_121 
+ bl[119] br[119] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_122 
+ bl[120] br[120] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_123 
+ bl[121] br[121] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_124 
+ bl[122] br[122] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_125 
+ bl[123] br[123] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_126 
+ bl[124] br[124] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_127 
+ bl[125] br[125] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_128 
+ bl[126] br[126] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_129 
+ bl[127] br[127] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_130 
+ bl[128] br[128] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_131 
+ bl[129] br[129] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_132 
+ bl[130] br[130] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_133 
+ bl[131] br[131] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_134 
+ bl[132] br[132] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_135 
+ bl[133] br[133] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_136 
+ bl[134] br[134] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_137 
+ bl[135] br[135] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_138 
+ bl[136] br[136] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_139 
+ bl[137] br[137] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_140 
+ bl[138] br[138] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_141 
+ bl[139] br[139] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_142 
+ bl[140] br[140] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_143 
+ bl[141] br[141] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_144 
+ bl[142] br[142] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_145 
+ bl[143] br[143] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_146 
+ bl[144] br[144] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_147 
+ bl[145] br[145] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_148 
+ bl[146] br[146] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_149 
+ bl[147] br[147] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_150 
+ bl[148] br[148] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_151 
+ bl[149] br[149] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_152 
+ bl[150] br[150] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_153 
+ bl[151] br[151] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_154 
+ bl[152] br[152] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_155 
+ bl[153] br[153] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_156 
+ bl[154] br[154] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_157 
+ bl[155] br[155] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_158 
+ bl[156] br[156] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_159 
+ bl[157] br[157] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_160 
+ bl[158] br[158] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_161 
+ bl[159] br[159] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_162 
+ bl[160] br[160] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_163 
+ bl[161] br[161] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_164 
+ bl[162] br[162] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_165 
+ bl[163] br[163] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_166 
+ bl[164] br[164] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_167 
+ bl[165] br[165] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_168 
+ bl[166] br[166] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_169 
+ bl[167] br[167] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_170 
+ bl[168] br[168] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_171 
+ bl[169] br[169] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_172 
+ bl[170] br[170] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_173 
+ bl[171] br[171] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_174 
+ bl[172] br[172] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_175 
+ bl[173] br[173] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_176 
+ bl[174] br[174] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_177 
+ bl[175] br[175] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_178 
+ bl[176] br[176] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_179 
+ bl[177] br[177] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_180 
+ bl[178] br[178] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_181 
+ bl[179] br[179] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_182 
+ bl[180] br[180] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_183 
+ bl[181] br[181] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_184 
+ bl[182] br[182] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_185 
+ bl[183] br[183] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_186 
+ bl[184] br[184] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_187 
+ bl[185] br[185] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_188 
+ bl[186] br[186] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_189 
+ bl[187] br[187] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_190 
+ bl[188] br[188] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_191 
+ bl[189] br[189] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_192 
+ bl[190] br[190] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_193 
+ bl[191] br[191] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_194 
+ bl[192] br[192] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_195 
+ bl[193] br[193] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_196 
+ bl[194] br[194] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_197 
+ bl[195] br[195] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_198 
+ bl[196] br[196] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_199 
+ bl[197] br[197] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_200 
+ bl[198] br[198] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_201 
+ bl[199] br[199] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_202 
+ bl[200] br[200] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_203 
+ bl[201] br[201] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_204 
+ bl[202] br[202] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_205 
+ bl[203] br[203] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_206 
+ bl[204] br[204] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_207 
+ bl[205] br[205] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_208 
+ bl[206] br[206] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_209 
+ bl[207] br[207] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_210 
+ bl[208] br[208] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_211 
+ bl[209] br[209] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_212 
+ bl[210] br[210] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_213 
+ bl[211] br[211] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_214 
+ bl[212] br[212] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_215 
+ bl[213] br[213] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_216 
+ bl[214] br[214] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_217 
+ bl[215] br[215] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_218 
+ bl[216] br[216] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_219 
+ bl[217] br[217] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_220 
+ bl[218] br[218] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_221 
+ bl[219] br[219] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_222 
+ bl[220] br[220] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_223 
+ bl[221] br[221] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_224 
+ bl[222] br[222] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_225 
+ bl[223] br[223] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_226 
+ bl[224] br[224] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_227 
+ bl[225] br[225] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_228 
+ bl[226] br[226] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_229 
+ bl[227] br[227] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_230 
+ bl[228] br[228] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_231 
+ bl[229] br[229] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_232 
+ bl[230] br[230] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_233 
+ bl[231] br[231] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_234 
+ bl[232] br[232] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_235 
+ bl[233] br[233] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_236 
+ bl[234] br[234] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_237 
+ bl[235] br[235] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_238 
+ bl[236] br[236] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_239 
+ bl[237] br[237] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_240 
+ bl[238] br[238] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_241 
+ bl[239] br[239] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_242 
+ bl[240] br[240] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_243 
+ bl[241] br[241] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_244 
+ bl[242] br[242] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_245 
+ bl[243] br[243] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_246 
+ bl[244] br[244] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_247 
+ bl[245] br[245] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_248 
+ bl[246] br[246] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_249 
+ bl[247] br[247] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_250 
+ bl[248] br[248] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_251 
+ bl[249] br[249] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_252 
+ bl[250] br[250] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_253 
+ bl[251] br[251] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_254 
+ bl[252] br[252] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_255 
+ bl[253] br[253] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_256 
+ bl[254] br[254] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_257 
+ bl[255] br[255] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_258 
+ vdd vdd vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_259 
+ vdd vdd vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_0 
+ vdd vdd vss vdd vpb vnb wl[97] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_99_1 
+ rbl rbr vss vdd vpb vnb wl[97] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_99_2 
+ bl[0] br[0] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_3 
+ bl[1] br[1] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_4 
+ bl[2] br[2] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_5 
+ bl[3] br[3] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_6 
+ bl[4] br[4] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_7 
+ bl[5] br[5] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_8 
+ bl[6] br[6] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_9 
+ bl[7] br[7] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_10 
+ bl[8] br[8] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_11 
+ bl[9] br[9] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_12 
+ bl[10] br[10] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_13 
+ bl[11] br[11] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_14 
+ bl[12] br[12] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_15 
+ bl[13] br[13] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_16 
+ bl[14] br[14] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_17 
+ bl[15] br[15] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_18 
+ bl[16] br[16] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_19 
+ bl[17] br[17] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_20 
+ bl[18] br[18] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_21 
+ bl[19] br[19] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_22 
+ bl[20] br[20] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_23 
+ bl[21] br[21] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_24 
+ bl[22] br[22] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_25 
+ bl[23] br[23] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_26 
+ bl[24] br[24] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_27 
+ bl[25] br[25] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_28 
+ bl[26] br[26] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_29 
+ bl[27] br[27] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_30 
+ bl[28] br[28] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_31 
+ bl[29] br[29] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_32 
+ bl[30] br[30] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_33 
+ bl[31] br[31] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_34 
+ bl[32] br[32] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_35 
+ bl[33] br[33] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_36 
+ bl[34] br[34] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_37 
+ bl[35] br[35] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_38 
+ bl[36] br[36] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_39 
+ bl[37] br[37] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_40 
+ bl[38] br[38] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_41 
+ bl[39] br[39] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_42 
+ bl[40] br[40] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_43 
+ bl[41] br[41] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_44 
+ bl[42] br[42] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_45 
+ bl[43] br[43] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_46 
+ bl[44] br[44] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_47 
+ bl[45] br[45] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_48 
+ bl[46] br[46] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_49 
+ bl[47] br[47] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_50 
+ bl[48] br[48] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_51 
+ bl[49] br[49] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_52 
+ bl[50] br[50] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_53 
+ bl[51] br[51] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_54 
+ bl[52] br[52] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_55 
+ bl[53] br[53] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_56 
+ bl[54] br[54] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_57 
+ bl[55] br[55] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_58 
+ bl[56] br[56] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_59 
+ bl[57] br[57] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_60 
+ bl[58] br[58] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_61 
+ bl[59] br[59] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_62 
+ bl[60] br[60] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_63 
+ bl[61] br[61] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_64 
+ bl[62] br[62] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_65 
+ bl[63] br[63] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_66 
+ bl[64] br[64] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_67 
+ bl[65] br[65] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_68 
+ bl[66] br[66] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_69 
+ bl[67] br[67] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_70 
+ bl[68] br[68] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_71 
+ bl[69] br[69] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_72 
+ bl[70] br[70] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_73 
+ bl[71] br[71] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_74 
+ bl[72] br[72] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_75 
+ bl[73] br[73] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_76 
+ bl[74] br[74] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_77 
+ bl[75] br[75] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_78 
+ bl[76] br[76] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_79 
+ bl[77] br[77] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_80 
+ bl[78] br[78] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_81 
+ bl[79] br[79] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_82 
+ bl[80] br[80] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_83 
+ bl[81] br[81] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_84 
+ bl[82] br[82] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_85 
+ bl[83] br[83] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_86 
+ bl[84] br[84] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_87 
+ bl[85] br[85] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_88 
+ bl[86] br[86] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_89 
+ bl[87] br[87] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_90 
+ bl[88] br[88] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_91 
+ bl[89] br[89] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_92 
+ bl[90] br[90] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_93 
+ bl[91] br[91] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_94 
+ bl[92] br[92] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_95 
+ bl[93] br[93] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_96 
+ bl[94] br[94] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_97 
+ bl[95] br[95] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_98 
+ bl[96] br[96] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_99 
+ bl[97] br[97] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_100 
+ bl[98] br[98] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_101 
+ bl[99] br[99] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_102 
+ bl[100] br[100] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_103 
+ bl[101] br[101] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_104 
+ bl[102] br[102] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_105 
+ bl[103] br[103] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_106 
+ bl[104] br[104] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_107 
+ bl[105] br[105] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_108 
+ bl[106] br[106] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_109 
+ bl[107] br[107] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_110 
+ bl[108] br[108] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_111 
+ bl[109] br[109] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_112 
+ bl[110] br[110] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_113 
+ bl[111] br[111] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_114 
+ bl[112] br[112] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_115 
+ bl[113] br[113] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_116 
+ bl[114] br[114] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_117 
+ bl[115] br[115] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_118 
+ bl[116] br[116] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_119 
+ bl[117] br[117] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_120 
+ bl[118] br[118] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_121 
+ bl[119] br[119] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_122 
+ bl[120] br[120] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_123 
+ bl[121] br[121] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_124 
+ bl[122] br[122] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_125 
+ bl[123] br[123] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_126 
+ bl[124] br[124] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_127 
+ bl[125] br[125] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_128 
+ bl[126] br[126] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_129 
+ bl[127] br[127] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_130 
+ bl[128] br[128] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_131 
+ bl[129] br[129] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_132 
+ bl[130] br[130] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_133 
+ bl[131] br[131] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_134 
+ bl[132] br[132] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_135 
+ bl[133] br[133] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_136 
+ bl[134] br[134] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_137 
+ bl[135] br[135] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_138 
+ bl[136] br[136] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_139 
+ bl[137] br[137] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_140 
+ bl[138] br[138] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_141 
+ bl[139] br[139] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_142 
+ bl[140] br[140] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_143 
+ bl[141] br[141] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_144 
+ bl[142] br[142] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_145 
+ bl[143] br[143] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_146 
+ bl[144] br[144] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_147 
+ bl[145] br[145] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_148 
+ bl[146] br[146] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_149 
+ bl[147] br[147] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_150 
+ bl[148] br[148] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_151 
+ bl[149] br[149] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_152 
+ bl[150] br[150] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_153 
+ bl[151] br[151] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_154 
+ bl[152] br[152] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_155 
+ bl[153] br[153] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_156 
+ bl[154] br[154] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_157 
+ bl[155] br[155] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_158 
+ bl[156] br[156] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_159 
+ bl[157] br[157] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_160 
+ bl[158] br[158] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_161 
+ bl[159] br[159] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_162 
+ bl[160] br[160] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_163 
+ bl[161] br[161] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_164 
+ bl[162] br[162] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_165 
+ bl[163] br[163] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_166 
+ bl[164] br[164] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_167 
+ bl[165] br[165] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_168 
+ bl[166] br[166] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_169 
+ bl[167] br[167] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_170 
+ bl[168] br[168] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_171 
+ bl[169] br[169] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_172 
+ bl[170] br[170] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_173 
+ bl[171] br[171] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_174 
+ bl[172] br[172] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_175 
+ bl[173] br[173] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_176 
+ bl[174] br[174] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_177 
+ bl[175] br[175] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_178 
+ bl[176] br[176] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_179 
+ bl[177] br[177] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_180 
+ bl[178] br[178] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_181 
+ bl[179] br[179] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_182 
+ bl[180] br[180] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_183 
+ bl[181] br[181] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_184 
+ bl[182] br[182] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_185 
+ bl[183] br[183] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_186 
+ bl[184] br[184] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_187 
+ bl[185] br[185] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_188 
+ bl[186] br[186] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_189 
+ bl[187] br[187] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_190 
+ bl[188] br[188] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_191 
+ bl[189] br[189] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_192 
+ bl[190] br[190] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_193 
+ bl[191] br[191] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_194 
+ bl[192] br[192] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_195 
+ bl[193] br[193] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_196 
+ bl[194] br[194] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_197 
+ bl[195] br[195] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_198 
+ bl[196] br[196] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_199 
+ bl[197] br[197] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_200 
+ bl[198] br[198] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_201 
+ bl[199] br[199] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_202 
+ bl[200] br[200] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_203 
+ bl[201] br[201] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_204 
+ bl[202] br[202] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_205 
+ bl[203] br[203] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_206 
+ bl[204] br[204] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_207 
+ bl[205] br[205] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_208 
+ bl[206] br[206] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_209 
+ bl[207] br[207] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_210 
+ bl[208] br[208] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_211 
+ bl[209] br[209] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_212 
+ bl[210] br[210] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_213 
+ bl[211] br[211] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_214 
+ bl[212] br[212] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_215 
+ bl[213] br[213] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_216 
+ bl[214] br[214] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_217 
+ bl[215] br[215] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_218 
+ bl[216] br[216] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_219 
+ bl[217] br[217] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_220 
+ bl[218] br[218] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_221 
+ bl[219] br[219] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_222 
+ bl[220] br[220] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_223 
+ bl[221] br[221] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_224 
+ bl[222] br[222] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_225 
+ bl[223] br[223] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_226 
+ bl[224] br[224] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_227 
+ bl[225] br[225] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_228 
+ bl[226] br[226] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_229 
+ bl[227] br[227] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_230 
+ bl[228] br[228] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_231 
+ bl[229] br[229] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_232 
+ bl[230] br[230] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_233 
+ bl[231] br[231] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_234 
+ bl[232] br[232] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_235 
+ bl[233] br[233] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_236 
+ bl[234] br[234] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_237 
+ bl[235] br[235] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_238 
+ bl[236] br[236] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_239 
+ bl[237] br[237] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_240 
+ bl[238] br[238] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_241 
+ bl[239] br[239] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_242 
+ bl[240] br[240] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_243 
+ bl[241] br[241] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_244 
+ bl[242] br[242] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_245 
+ bl[243] br[243] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_246 
+ bl[244] br[244] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_247 
+ bl[245] br[245] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_248 
+ bl[246] br[246] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_249 
+ bl[247] br[247] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_250 
+ bl[248] br[248] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_251 
+ bl[249] br[249] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_252 
+ bl[250] br[250] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_253 
+ bl[251] br[251] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_254 
+ bl[252] br[252] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_255 
+ bl[253] br[253] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_256 
+ bl[254] br[254] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_257 
+ bl[255] br[255] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_258 
+ vdd vdd vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_259 
+ vdd vdd vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_0 
+ vdd vdd vss vdd vpb vnb wl[98] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_100_1 
+ rbl rbr vss vdd vpb vnb wl[98] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_100_2 
+ bl[0] br[0] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_3 
+ bl[1] br[1] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_4 
+ bl[2] br[2] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_5 
+ bl[3] br[3] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_6 
+ bl[4] br[4] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_7 
+ bl[5] br[5] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_8 
+ bl[6] br[6] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_9 
+ bl[7] br[7] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_10 
+ bl[8] br[8] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_11 
+ bl[9] br[9] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_12 
+ bl[10] br[10] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_13 
+ bl[11] br[11] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_14 
+ bl[12] br[12] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_15 
+ bl[13] br[13] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_16 
+ bl[14] br[14] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_17 
+ bl[15] br[15] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_18 
+ bl[16] br[16] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_19 
+ bl[17] br[17] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_20 
+ bl[18] br[18] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_21 
+ bl[19] br[19] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_22 
+ bl[20] br[20] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_23 
+ bl[21] br[21] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_24 
+ bl[22] br[22] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_25 
+ bl[23] br[23] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_26 
+ bl[24] br[24] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_27 
+ bl[25] br[25] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_28 
+ bl[26] br[26] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_29 
+ bl[27] br[27] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_30 
+ bl[28] br[28] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_31 
+ bl[29] br[29] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_32 
+ bl[30] br[30] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_33 
+ bl[31] br[31] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_34 
+ bl[32] br[32] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_35 
+ bl[33] br[33] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_36 
+ bl[34] br[34] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_37 
+ bl[35] br[35] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_38 
+ bl[36] br[36] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_39 
+ bl[37] br[37] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_40 
+ bl[38] br[38] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_41 
+ bl[39] br[39] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_42 
+ bl[40] br[40] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_43 
+ bl[41] br[41] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_44 
+ bl[42] br[42] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_45 
+ bl[43] br[43] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_46 
+ bl[44] br[44] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_47 
+ bl[45] br[45] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_48 
+ bl[46] br[46] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_49 
+ bl[47] br[47] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_50 
+ bl[48] br[48] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_51 
+ bl[49] br[49] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_52 
+ bl[50] br[50] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_53 
+ bl[51] br[51] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_54 
+ bl[52] br[52] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_55 
+ bl[53] br[53] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_56 
+ bl[54] br[54] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_57 
+ bl[55] br[55] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_58 
+ bl[56] br[56] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_59 
+ bl[57] br[57] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_60 
+ bl[58] br[58] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_61 
+ bl[59] br[59] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_62 
+ bl[60] br[60] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_63 
+ bl[61] br[61] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_64 
+ bl[62] br[62] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_65 
+ bl[63] br[63] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_66 
+ bl[64] br[64] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_67 
+ bl[65] br[65] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_68 
+ bl[66] br[66] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_69 
+ bl[67] br[67] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_70 
+ bl[68] br[68] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_71 
+ bl[69] br[69] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_72 
+ bl[70] br[70] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_73 
+ bl[71] br[71] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_74 
+ bl[72] br[72] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_75 
+ bl[73] br[73] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_76 
+ bl[74] br[74] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_77 
+ bl[75] br[75] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_78 
+ bl[76] br[76] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_79 
+ bl[77] br[77] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_80 
+ bl[78] br[78] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_81 
+ bl[79] br[79] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_82 
+ bl[80] br[80] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_83 
+ bl[81] br[81] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_84 
+ bl[82] br[82] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_85 
+ bl[83] br[83] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_86 
+ bl[84] br[84] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_87 
+ bl[85] br[85] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_88 
+ bl[86] br[86] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_89 
+ bl[87] br[87] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_90 
+ bl[88] br[88] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_91 
+ bl[89] br[89] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_92 
+ bl[90] br[90] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_93 
+ bl[91] br[91] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_94 
+ bl[92] br[92] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_95 
+ bl[93] br[93] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_96 
+ bl[94] br[94] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_97 
+ bl[95] br[95] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_98 
+ bl[96] br[96] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_99 
+ bl[97] br[97] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_100 
+ bl[98] br[98] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_101 
+ bl[99] br[99] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_102 
+ bl[100] br[100] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_103 
+ bl[101] br[101] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_104 
+ bl[102] br[102] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_105 
+ bl[103] br[103] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_106 
+ bl[104] br[104] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_107 
+ bl[105] br[105] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_108 
+ bl[106] br[106] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_109 
+ bl[107] br[107] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_110 
+ bl[108] br[108] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_111 
+ bl[109] br[109] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_112 
+ bl[110] br[110] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_113 
+ bl[111] br[111] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_114 
+ bl[112] br[112] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_115 
+ bl[113] br[113] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_116 
+ bl[114] br[114] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_117 
+ bl[115] br[115] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_118 
+ bl[116] br[116] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_119 
+ bl[117] br[117] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_120 
+ bl[118] br[118] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_121 
+ bl[119] br[119] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_122 
+ bl[120] br[120] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_123 
+ bl[121] br[121] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_124 
+ bl[122] br[122] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_125 
+ bl[123] br[123] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_126 
+ bl[124] br[124] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_127 
+ bl[125] br[125] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_128 
+ bl[126] br[126] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_129 
+ bl[127] br[127] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_130 
+ bl[128] br[128] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_131 
+ bl[129] br[129] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_132 
+ bl[130] br[130] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_133 
+ bl[131] br[131] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_134 
+ bl[132] br[132] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_135 
+ bl[133] br[133] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_136 
+ bl[134] br[134] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_137 
+ bl[135] br[135] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_138 
+ bl[136] br[136] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_139 
+ bl[137] br[137] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_140 
+ bl[138] br[138] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_141 
+ bl[139] br[139] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_142 
+ bl[140] br[140] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_143 
+ bl[141] br[141] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_144 
+ bl[142] br[142] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_145 
+ bl[143] br[143] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_146 
+ bl[144] br[144] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_147 
+ bl[145] br[145] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_148 
+ bl[146] br[146] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_149 
+ bl[147] br[147] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_150 
+ bl[148] br[148] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_151 
+ bl[149] br[149] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_152 
+ bl[150] br[150] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_153 
+ bl[151] br[151] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_154 
+ bl[152] br[152] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_155 
+ bl[153] br[153] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_156 
+ bl[154] br[154] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_157 
+ bl[155] br[155] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_158 
+ bl[156] br[156] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_159 
+ bl[157] br[157] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_160 
+ bl[158] br[158] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_161 
+ bl[159] br[159] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_162 
+ bl[160] br[160] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_163 
+ bl[161] br[161] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_164 
+ bl[162] br[162] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_165 
+ bl[163] br[163] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_166 
+ bl[164] br[164] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_167 
+ bl[165] br[165] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_168 
+ bl[166] br[166] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_169 
+ bl[167] br[167] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_170 
+ bl[168] br[168] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_171 
+ bl[169] br[169] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_172 
+ bl[170] br[170] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_173 
+ bl[171] br[171] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_174 
+ bl[172] br[172] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_175 
+ bl[173] br[173] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_176 
+ bl[174] br[174] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_177 
+ bl[175] br[175] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_178 
+ bl[176] br[176] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_179 
+ bl[177] br[177] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_180 
+ bl[178] br[178] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_181 
+ bl[179] br[179] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_182 
+ bl[180] br[180] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_183 
+ bl[181] br[181] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_184 
+ bl[182] br[182] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_185 
+ bl[183] br[183] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_186 
+ bl[184] br[184] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_187 
+ bl[185] br[185] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_188 
+ bl[186] br[186] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_189 
+ bl[187] br[187] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_190 
+ bl[188] br[188] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_191 
+ bl[189] br[189] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_192 
+ bl[190] br[190] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_193 
+ bl[191] br[191] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_194 
+ bl[192] br[192] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_195 
+ bl[193] br[193] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_196 
+ bl[194] br[194] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_197 
+ bl[195] br[195] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_198 
+ bl[196] br[196] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_199 
+ bl[197] br[197] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_200 
+ bl[198] br[198] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_201 
+ bl[199] br[199] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_202 
+ bl[200] br[200] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_203 
+ bl[201] br[201] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_204 
+ bl[202] br[202] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_205 
+ bl[203] br[203] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_206 
+ bl[204] br[204] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_207 
+ bl[205] br[205] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_208 
+ bl[206] br[206] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_209 
+ bl[207] br[207] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_210 
+ bl[208] br[208] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_211 
+ bl[209] br[209] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_212 
+ bl[210] br[210] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_213 
+ bl[211] br[211] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_214 
+ bl[212] br[212] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_215 
+ bl[213] br[213] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_216 
+ bl[214] br[214] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_217 
+ bl[215] br[215] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_218 
+ bl[216] br[216] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_219 
+ bl[217] br[217] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_220 
+ bl[218] br[218] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_221 
+ bl[219] br[219] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_222 
+ bl[220] br[220] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_223 
+ bl[221] br[221] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_224 
+ bl[222] br[222] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_225 
+ bl[223] br[223] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_226 
+ bl[224] br[224] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_227 
+ bl[225] br[225] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_228 
+ bl[226] br[226] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_229 
+ bl[227] br[227] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_230 
+ bl[228] br[228] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_231 
+ bl[229] br[229] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_232 
+ bl[230] br[230] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_233 
+ bl[231] br[231] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_234 
+ bl[232] br[232] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_235 
+ bl[233] br[233] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_236 
+ bl[234] br[234] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_237 
+ bl[235] br[235] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_238 
+ bl[236] br[236] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_239 
+ bl[237] br[237] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_240 
+ bl[238] br[238] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_241 
+ bl[239] br[239] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_242 
+ bl[240] br[240] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_243 
+ bl[241] br[241] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_244 
+ bl[242] br[242] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_245 
+ bl[243] br[243] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_246 
+ bl[244] br[244] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_247 
+ bl[245] br[245] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_248 
+ bl[246] br[246] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_249 
+ bl[247] br[247] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_250 
+ bl[248] br[248] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_251 
+ bl[249] br[249] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_252 
+ bl[250] br[250] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_253 
+ bl[251] br[251] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_254 
+ bl[252] br[252] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_255 
+ bl[253] br[253] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_256 
+ bl[254] br[254] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_257 
+ bl[255] br[255] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_258 
+ vdd vdd vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_259 
+ vdd vdd vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_0 
+ vdd vdd vss vdd vpb vnb wl[99] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_101_1 
+ rbl rbr vss vdd vpb vnb wl[99] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_101_2 
+ bl[0] br[0] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_3 
+ bl[1] br[1] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_4 
+ bl[2] br[2] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_5 
+ bl[3] br[3] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_6 
+ bl[4] br[4] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_7 
+ bl[5] br[5] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_8 
+ bl[6] br[6] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_9 
+ bl[7] br[7] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_10 
+ bl[8] br[8] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_11 
+ bl[9] br[9] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_12 
+ bl[10] br[10] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_13 
+ bl[11] br[11] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_14 
+ bl[12] br[12] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_15 
+ bl[13] br[13] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_16 
+ bl[14] br[14] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_17 
+ bl[15] br[15] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_18 
+ bl[16] br[16] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_19 
+ bl[17] br[17] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_20 
+ bl[18] br[18] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_21 
+ bl[19] br[19] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_22 
+ bl[20] br[20] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_23 
+ bl[21] br[21] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_24 
+ bl[22] br[22] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_25 
+ bl[23] br[23] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_26 
+ bl[24] br[24] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_27 
+ bl[25] br[25] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_28 
+ bl[26] br[26] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_29 
+ bl[27] br[27] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_30 
+ bl[28] br[28] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_31 
+ bl[29] br[29] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_32 
+ bl[30] br[30] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_33 
+ bl[31] br[31] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_34 
+ bl[32] br[32] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_35 
+ bl[33] br[33] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_36 
+ bl[34] br[34] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_37 
+ bl[35] br[35] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_38 
+ bl[36] br[36] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_39 
+ bl[37] br[37] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_40 
+ bl[38] br[38] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_41 
+ bl[39] br[39] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_42 
+ bl[40] br[40] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_43 
+ bl[41] br[41] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_44 
+ bl[42] br[42] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_45 
+ bl[43] br[43] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_46 
+ bl[44] br[44] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_47 
+ bl[45] br[45] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_48 
+ bl[46] br[46] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_49 
+ bl[47] br[47] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_50 
+ bl[48] br[48] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_51 
+ bl[49] br[49] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_52 
+ bl[50] br[50] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_53 
+ bl[51] br[51] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_54 
+ bl[52] br[52] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_55 
+ bl[53] br[53] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_56 
+ bl[54] br[54] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_57 
+ bl[55] br[55] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_58 
+ bl[56] br[56] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_59 
+ bl[57] br[57] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_60 
+ bl[58] br[58] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_61 
+ bl[59] br[59] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_62 
+ bl[60] br[60] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_63 
+ bl[61] br[61] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_64 
+ bl[62] br[62] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_65 
+ bl[63] br[63] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_66 
+ bl[64] br[64] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_67 
+ bl[65] br[65] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_68 
+ bl[66] br[66] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_69 
+ bl[67] br[67] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_70 
+ bl[68] br[68] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_71 
+ bl[69] br[69] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_72 
+ bl[70] br[70] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_73 
+ bl[71] br[71] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_74 
+ bl[72] br[72] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_75 
+ bl[73] br[73] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_76 
+ bl[74] br[74] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_77 
+ bl[75] br[75] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_78 
+ bl[76] br[76] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_79 
+ bl[77] br[77] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_80 
+ bl[78] br[78] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_81 
+ bl[79] br[79] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_82 
+ bl[80] br[80] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_83 
+ bl[81] br[81] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_84 
+ bl[82] br[82] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_85 
+ bl[83] br[83] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_86 
+ bl[84] br[84] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_87 
+ bl[85] br[85] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_88 
+ bl[86] br[86] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_89 
+ bl[87] br[87] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_90 
+ bl[88] br[88] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_91 
+ bl[89] br[89] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_92 
+ bl[90] br[90] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_93 
+ bl[91] br[91] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_94 
+ bl[92] br[92] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_95 
+ bl[93] br[93] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_96 
+ bl[94] br[94] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_97 
+ bl[95] br[95] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_98 
+ bl[96] br[96] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_99 
+ bl[97] br[97] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_100 
+ bl[98] br[98] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_101 
+ bl[99] br[99] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_102 
+ bl[100] br[100] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_103 
+ bl[101] br[101] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_104 
+ bl[102] br[102] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_105 
+ bl[103] br[103] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_106 
+ bl[104] br[104] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_107 
+ bl[105] br[105] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_108 
+ bl[106] br[106] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_109 
+ bl[107] br[107] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_110 
+ bl[108] br[108] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_111 
+ bl[109] br[109] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_112 
+ bl[110] br[110] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_113 
+ bl[111] br[111] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_114 
+ bl[112] br[112] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_115 
+ bl[113] br[113] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_116 
+ bl[114] br[114] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_117 
+ bl[115] br[115] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_118 
+ bl[116] br[116] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_119 
+ bl[117] br[117] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_120 
+ bl[118] br[118] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_121 
+ bl[119] br[119] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_122 
+ bl[120] br[120] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_123 
+ bl[121] br[121] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_124 
+ bl[122] br[122] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_125 
+ bl[123] br[123] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_126 
+ bl[124] br[124] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_127 
+ bl[125] br[125] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_128 
+ bl[126] br[126] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_129 
+ bl[127] br[127] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_130 
+ bl[128] br[128] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_131 
+ bl[129] br[129] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_132 
+ bl[130] br[130] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_133 
+ bl[131] br[131] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_134 
+ bl[132] br[132] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_135 
+ bl[133] br[133] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_136 
+ bl[134] br[134] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_137 
+ bl[135] br[135] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_138 
+ bl[136] br[136] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_139 
+ bl[137] br[137] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_140 
+ bl[138] br[138] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_141 
+ bl[139] br[139] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_142 
+ bl[140] br[140] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_143 
+ bl[141] br[141] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_144 
+ bl[142] br[142] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_145 
+ bl[143] br[143] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_146 
+ bl[144] br[144] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_147 
+ bl[145] br[145] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_148 
+ bl[146] br[146] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_149 
+ bl[147] br[147] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_150 
+ bl[148] br[148] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_151 
+ bl[149] br[149] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_152 
+ bl[150] br[150] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_153 
+ bl[151] br[151] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_154 
+ bl[152] br[152] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_155 
+ bl[153] br[153] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_156 
+ bl[154] br[154] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_157 
+ bl[155] br[155] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_158 
+ bl[156] br[156] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_159 
+ bl[157] br[157] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_160 
+ bl[158] br[158] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_161 
+ bl[159] br[159] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_162 
+ bl[160] br[160] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_163 
+ bl[161] br[161] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_164 
+ bl[162] br[162] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_165 
+ bl[163] br[163] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_166 
+ bl[164] br[164] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_167 
+ bl[165] br[165] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_168 
+ bl[166] br[166] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_169 
+ bl[167] br[167] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_170 
+ bl[168] br[168] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_171 
+ bl[169] br[169] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_172 
+ bl[170] br[170] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_173 
+ bl[171] br[171] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_174 
+ bl[172] br[172] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_175 
+ bl[173] br[173] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_176 
+ bl[174] br[174] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_177 
+ bl[175] br[175] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_178 
+ bl[176] br[176] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_179 
+ bl[177] br[177] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_180 
+ bl[178] br[178] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_181 
+ bl[179] br[179] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_182 
+ bl[180] br[180] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_183 
+ bl[181] br[181] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_184 
+ bl[182] br[182] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_185 
+ bl[183] br[183] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_186 
+ bl[184] br[184] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_187 
+ bl[185] br[185] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_188 
+ bl[186] br[186] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_189 
+ bl[187] br[187] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_190 
+ bl[188] br[188] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_191 
+ bl[189] br[189] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_192 
+ bl[190] br[190] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_193 
+ bl[191] br[191] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_194 
+ bl[192] br[192] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_195 
+ bl[193] br[193] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_196 
+ bl[194] br[194] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_197 
+ bl[195] br[195] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_198 
+ bl[196] br[196] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_199 
+ bl[197] br[197] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_200 
+ bl[198] br[198] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_201 
+ bl[199] br[199] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_202 
+ bl[200] br[200] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_203 
+ bl[201] br[201] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_204 
+ bl[202] br[202] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_205 
+ bl[203] br[203] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_206 
+ bl[204] br[204] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_207 
+ bl[205] br[205] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_208 
+ bl[206] br[206] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_209 
+ bl[207] br[207] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_210 
+ bl[208] br[208] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_211 
+ bl[209] br[209] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_212 
+ bl[210] br[210] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_213 
+ bl[211] br[211] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_214 
+ bl[212] br[212] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_215 
+ bl[213] br[213] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_216 
+ bl[214] br[214] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_217 
+ bl[215] br[215] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_218 
+ bl[216] br[216] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_219 
+ bl[217] br[217] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_220 
+ bl[218] br[218] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_221 
+ bl[219] br[219] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_222 
+ bl[220] br[220] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_223 
+ bl[221] br[221] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_224 
+ bl[222] br[222] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_225 
+ bl[223] br[223] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_226 
+ bl[224] br[224] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_227 
+ bl[225] br[225] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_228 
+ bl[226] br[226] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_229 
+ bl[227] br[227] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_230 
+ bl[228] br[228] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_231 
+ bl[229] br[229] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_232 
+ bl[230] br[230] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_233 
+ bl[231] br[231] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_234 
+ bl[232] br[232] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_235 
+ bl[233] br[233] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_236 
+ bl[234] br[234] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_237 
+ bl[235] br[235] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_238 
+ bl[236] br[236] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_239 
+ bl[237] br[237] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_240 
+ bl[238] br[238] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_241 
+ bl[239] br[239] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_242 
+ bl[240] br[240] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_243 
+ bl[241] br[241] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_244 
+ bl[242] br[242] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_245 
+ bl[243] br[243] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_246 
+ bl[244] br[244] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_247 
+ bl[245] br[245] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_248 
+ bl[246] br[246] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_249 
+ bl[247] br[247] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_250 
+ bl[248] br[248] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_251 
+ bl[249] br[249] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_252 
+ bl[250] br[250] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_253 
+ bl[251] br[251] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_254 
+ bl[252] br[252] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_255 
+ bl[253] br[253] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_256 
+ bl[254] br[254] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_257 
+ bl[255] br[255] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_258 
+ vdd vdd vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_259 
+ vdd vdd vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_0 
+ vdd vdd vss vdd vpb vnb wl[100] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_102_1 
+ rbl rbr vss vdd vpb vnb wl[100] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_102_2 
+ bl[0] br[0] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_3 
+ bl[1] br[1] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_4 
+ bl[2] br[2] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_5 
+ bl[3] br[3] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_6 
+ bl[4] br[4] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_7 
+ bl[5] br[5] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_8 
+ bl[6] br[6] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_9 
+ bl[7] br[7] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_10 
+ bl[8] br[8] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_11 
+ bl[9] br[9] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_12 
+ bl[10] br[10] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_13 
+ bl[11] br[11] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_14 
+ bl[12] br[12] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_15 
+ bl[13] br[13] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_16 
+ bl[14] br[14] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_17 
+ bl[15] br[15] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_18 
+ bl[16] br[16] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_19 
+ bl[17] br[17] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_20 
+ bl[18] br[18] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_21 
+ bl[19] br[19] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_22 
+ bl[20] br[20] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_23 
+ bl[21] br[21] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_24 
+ bl[22] br[22] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_25 
+ bl[23] br[23] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_26 
+ bl[24] br[24] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_27 
+ bl[25] br[25] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_28 
+ bl[26] br[26] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_29 
+ bl[27] br[27] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_30 
+ bl[28] br[28] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_31 
+ bl[29] br[29] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_32 
+ bl[30] br[30] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_33 
+ bl[31] br[31] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_34 
+ bl[32] br[32] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_35 
+ bl[33] br[33] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_36 
+ bl[34] br[34] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_37 
+ bl[35] br[35] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_38 
+ bl[36] br[36] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_39 
+ bl[37] br[37] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_40 
+ bl[38] br[38] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_41 
+ bl[39] br[39] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_42 
+ bl[40] br[40] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_43 
+ bl[41] br[41] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_44 
+ bl[42] br[42] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_45 
+ bl[43] br[43] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_46 
+ bl[44] br[44] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_47 
+ bl[45] br[45] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_48 
+ bl[46] br[46] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_49 
+ bl[47] br[47] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_50 
+ bl[48] br[48] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_51 
+ bl[49] br[49] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_52 
+ bl[50] br[50] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_53 
+ bl[51] br[51] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_54 
+ bl[52] br[52] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_55 
+ bl[53] br[53] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_56 
+ bl[54] br[54] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_57 
+ bl[55] br[55] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_58 
+ bl[56] br[56] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_59 
+ bl[57] br[57] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_60 
+ bl[58] br[58] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_61 
+ bl[59] br[59] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_62 
+ bl[60] br[60] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_63 
+ bl[61] br[61] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_64 
+ bl[62] br[62] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_65 
+ bl[63] br[63] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_66 
+ bl[64] br[64] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_67 
+ bl[65] br[65] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_68 
+ bl[66] br[66] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_69 
+ bl[67] br[67] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_70 
+ bl[68] br[68] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_71 
+ bl[69] br[69] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_72 
+ bl[70] br[70] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_73 
+ bl[71] br[71] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_74 
+ bl[72] br[72] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_75 
+ bl[73] br[73] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_76 
+ bl[74] br[74] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_77 
+ bl[75] br[75] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_78 
+ bl[76] br[76] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_79 
+ bl[77] br[77] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_80 
+ bl[78] br[78] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_81 
+ bl[79] br[79] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_82 
+ bl[80] br[80] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_83 
+ bl[81] br[81] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_84 
+ bl[82] br[82] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_85 
+ bl[83] br[83] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_86 
+ bl[84] br[84] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_87 
+ bl[85] br[85] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_88 
+ bl[86] br[86] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_89 
+ bl[87] br[87] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_90 
+ bl[88] br[88] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_91 
+ bl[89] br[89] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_92 
+ bl[90] br[90] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_93 
+ bl[91] br[91] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_94 
+ bl[92] br[92] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_95 
+ bl[93] br[93] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_96 
+ bl[94] br[94] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_97 
+ bl[95] br[95] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_98 
+ bl[96] br[96] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_99 
+ bl[97] br[97] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_100 
+ bl[98] br[98] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_101 
+ bl[99] br[99] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_102 
+ bl[100] br[100] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_103 
+ bl[101] br[101] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_104 
+ bl[102] br[102] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_105 
+ bl[103] br[103] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_106 
+ bl[104] br[104] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_107 
+ bl[105] br[105] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_108 
+ bl[106] br[106] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_109 
+ bl[107] br[107] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_110 
+ bl[108] br[108] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_111 
+ bl[109] br[109] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_112 
+ bl[110] br[110] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_113 
+ bl[111] br[111] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_114 
+ bl[112] br[112] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_115 
+ bl[113] br[113] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_116 
+ bl[114] br[114] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_117 
+ bl[115] br[115] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_118 
+ bl[116] br[116] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_119 
+ bl[117] br[117] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_120 
+ bl[118] br[118] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_121 
+ bl[119] br[119] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_122 
+ bl[120] br[120] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_123 
+ bl[121] br[121] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_124 
+ bl[122] br[122] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_125 
+ bl[123] br[123] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_126 
+ bl[124] br[124] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_127 
+ bl[125] br[125] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_128 
+ bl[126] br[126] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_129 
+ bl[127] br[127] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_130 
+ bl[128] br[128] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_131 
+ bl[129] br[129] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_132 
+ bl[130] br[130] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_133 
+ bl[131] br[131] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_134 
+ bl[132] br[132] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_135 
+ bl[133] br[133] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_136 
+ bl[134] br[134] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_137 
+ bl[135] br[135] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_138 
+ bl[136] br[136] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_139 
+ bl[137] br[137] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_140 
+ bl[138] br[138] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_141 
+ bl[139] br[139] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_142 
+ bl[140] br[140] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_143 
+ bl[141] br[141] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_144 
+ bl[142] br[142] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_145 
+ bl[143] br[143] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_146 
+ bl[144] br[144] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_147 
+ bl[145] br[145] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_148 
+ bl[146] br[146] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_149 
+ bl[147] br[147] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_150 
+ bl[148] br[148] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_151 
+ bl[149] br[149] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_152 
+ bl[150] br[150] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_153 
+ bl[151] br[151] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_154 
+ bl[152] br[152] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_155 
+ bl[153] br[153] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_156 
+ bl[154] br[154] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_157 
+ bl[155] br[155] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_158 
+ bl[156] br[156] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_159 
+ bl[157] br[157] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_160 
+ bl[158] br[158] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_161 
+ bl[159] br[159] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_162 
+ bl[160] br[160] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_163 
+ bl[161] br[161] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_164 
+ bl[162] br[162] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_165 
+ bl[163] br[163] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_166 
+ bl[164] br[164] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_167 
+ bl[165] br[165] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_168 
+ bl[166] br[166] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_169 
+ bl[167] br[167] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_170 
+ bl[168] br[168] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_171 
+ bl[169] br[169] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_172 
+ bl[170] br[170] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_173 
+ bl[171] br[171] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_174 
+ bl[172] br[172] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_175 
+ bl[173] br[173] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_176 
+ bl[174] br[174] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_177 
+ bl[175] br[175] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_178 
+ bl[176] br[176] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_179 
+ bl[177] br[177] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_180 
+ bl[178] br[178] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_181 
+ bl[179] br[179] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_182 
+ bl[180] br[180] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_183 
+ bl[181] br[181] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_184 
+ bl[182] br[182] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_185 
+ bl[183] br[183] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_186 
+ bl[184] br[184] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_187 
+ bl[185] br[185] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_188 
+ bl[186] br[186] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_189 
+ bl[187] br[187] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_190 
+ bl[188] br[188] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_191 
+ bl[189] br[189] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_192 
+ bl[190] br[190] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_193 
+ bl[191] br[191] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_194 
+ bl[192] br[192] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_195 
+ bl[193] br[193] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_196 
+ bl[194] br[194] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_197 
+ bl[195] br[195] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_198 
+ bl[196] br[196] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_199 
+ bl[197] br[197] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_200 
+ bl[198] br[198] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_201 
+ bl[199] br[199] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_202 
+ bl[200] br[200] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_203 
+ bl[201] br[201] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_204 
+ bl[202] br[202] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_205 
+ bl[203] br[203] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_206 
+ bl[204] br[204] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_207 
+ bl[205] br[205] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_208 
+ bl[206] br[206] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_209 
+ bl[207] br[207] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_210 
+ bl[208] br[208] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_211 
+ bl[209] br[209] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_212 
+ bl[210] br[210] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_213 
+ bl[211] br[211] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_214 
+ bl[212] br[212] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_215 
+ bl[213] br[213] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_216 
+ bl[214] br[214] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_217 
+ bl[215] br[215] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_218 
+ bl[216] br[216] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_219 
+ bl[217] br[217] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_220 
+ bl[218] br[218] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_221 
+ bl[219] br[219] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_222 
+ bl[220] br[220] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_223 
+ bl[221] br[221] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_224 
+ bl[222] br[222] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_225 
+ bl[223] br[223] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_226 
+ bl[224] br[224] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_227 
+ bl[225] br[225] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_228 
+ bl[226] br[226] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_229 
+ bl[227] br[227] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_230 
+ bl[228] br[228] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_231 
+ bl[229] br[229] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_232 
+ bl[230] br[230] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_233 
+ bl[231] br[231] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_234 
+ bl[232] br[232] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_235 
+ bl[233] br[233] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_236 
+ bl[234] br[234] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_237 
+ bl[235] br[235] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_238 
+ bl[236] br[236] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_239 
+ bl[237] br[237] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_240 
+ bl[238] br[238] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_241 
+ bl[239] br[239] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_242 
+ bl[240] br[240] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_243 
+ bl[241] br[241] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_244 
+ bl[242] br[242] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_245 
+ bl[243] br[243] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_246 
+ bl[244] br[244] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_247 
+ bl[245] br[245] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_248 
+ bl[246] br[246] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_249 
+ bl[247] br[247] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_250 
+ bl[248] br[248] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_251 
+ bl[249] br[249] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_252 
+ bl[250] br[250] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_253 
+ bl[251] br[251] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_254 
+ bl[252] br[252] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_255 
+ bl[253] br[253] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_256 
+ bl[254] br[254] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_257 
+ bl[255] br[255] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_258 
+ vdd vdd vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_259 
+ vdd vdd vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_0 
+ vdd vdd vss vdd vpb vnb wl[101] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_103_1 
+ rbl rbr vss vdd vpb vnb wl[101] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_103_2 
+ bl[0] br[0] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_3 
+ bl[1] br[1] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_4 
+ bl[2] br[2] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_5 
+ bl[3] br[3] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_6 
+ bl[4] br[4] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_7 
+ bl[5] br[5] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_8 
+ bl[6] br[6] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_9 
+ bl[7] br[7] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_10 
+ bl[8] br[8] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_11 
+ bl[9] br[9] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_12 
+ bl[10] br[10] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_13 
+ bl[11] br[11] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_14 
+ bl[12] br[12] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_15 
+ bl[13] br[13] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_16 
+ bl[14] br[14] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_17 
+ bl[15] br[15] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_18 
+ bl[16] br[16] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_19 
+ bl[17] br[17] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_20 
+ bl[18] br[18] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_21 
+ bl[19] br[19] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_22 
+ bl[20] br[20] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_23 
+ bl[21] br[21] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_24 
+ bl[22] br[22] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_25 
+ bl[23] br[23] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_26 
+ bl[24] br[24] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_27 
+ bl[25] br[25] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_28 
+ bl[26] br[26] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_29 
+ bl[27] br[27] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_30 
+ bl[28] br[28] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_31 
+ bl[29] br[29] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_32 
+ bl[30] br[30] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_33 
+ bl[31] br[31] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_34 
+ bl[32] br[32] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_35 
+ bl[33] br[33] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_36 
+ bl[34] br[34] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_37 
+ bl[35] br[35] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_38 
+ bl[36] br[36] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_39 
+ bl[37] br[37] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_40 
+ bl[38] br[38] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_41 
+ bl[39] br[39] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_42 
+ bl[40] br[40] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_43 
+ bl[41] br[41] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_44 
+ bl[42] br[42] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_45 
+ bl[43] br[43] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_46 
+ bl[44] br[44] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_47 
+ bl[45] br[45] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_48 
+ bl[46] br[46] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_49 
+ bl[47] br[47] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_50 
+ bl[48] br[48] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_51 
+ bl[49] br[49] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_52 
+ bl[50] br[50] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_53 
+ bl[51] br[51] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_54 
+ bl[52] br[52] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_55 
+ bl[53] br[53] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_56 
+ bl[54] br[54] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_57 
+ bl[55] br[55] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_58 
+ bl[56] br[56] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_59 
+ bl[57] br[57] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_60 
+ bl[58] br[58] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_61 
+ bl[59] br[59] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_62 
+ bl[60] br[60] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_63 
+ bl[61] br[61] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_64 
+ bl[62] br[62] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_65 
+ bl[63] br[63] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_66 
+ bl[64] br[64] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_67 
+ bl[65] br[65] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_68 
+ bl[66] br[66] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_69 
+ bl[67] br[67] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_70 
+ bl[68] br[68] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_71 
+ bl[69] br[69] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_72 
+ bl[70] br[70] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_73 
+ bl[71] br[71] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_74 
+ bl[72] br[72] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_75 
+ bl[73] br[73] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_76 
+ bl[74] br[74] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_77 
+ bl[75] br[75] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_78 
+ bl[76] br[76] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_79 
+ bl[77] br[77] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_80 
+ bl[78] br[78] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_81 
+ bl[79] br[79] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_82 
+ bl[80] br[80] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_83 
+ bl[81] br[81] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_84 
+ bl[82] br[82] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_85 
+ bl[83] br[83] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_86 
+ bl[84] br[84] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_87 
+ bl[85] br[85] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_88 
+ bl[86] br[86] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_89 
+ bl[87] br[87] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_90 
+ bl[88] br[88] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_91 
+ bl[89] br[89] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_92 
+ bl[90] br[90] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_93 
+ bl[91] br[91] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_94 
+ bl[92] br[92] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_95 
+ bl[93] br[93] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_96 
+ bl[94] br[94] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_97 
+ bl[95] br[95] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_98 
+ bl[96] br[96] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_99 
+ bl[97] br[97] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_100 
+ bl[98] br[98] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_101 
+ bl[99] br[99] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_102 
+ bl[100] br[100] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_103 
+ bl[101] br[101] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_104 
+ bl[102] br[102] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_105 
+ bl[103] br[103] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_106 
+ bl[104] br[104] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_107 
+ bl[105] br[105] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_108 
+ bl[106] br[106] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_109 
+ bl[107] br[107] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_110 
+ bl[108] br[108] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_111 
+ bl[109] br[109] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_112 
+ bl[110] br[110] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_113 
+ bl[111] br[111] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_114 
+ bl[112] br[112] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_115 
+ bl[113] br[113] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_116 
+ bl[114] br[114] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_117 
+ bl[115] br[115] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_118 
+ bl[116] br[116] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_119 
+ bl[117] br[117] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_120 
+ bl[118] br[118] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_121 
+ bl[119] br[119] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_122 
+ bl[120] br[120] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_123 
+ bl[121] br[121] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_124 
+ bl[122] br[122] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_125 
+ bl[123] br[123] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_126 
+ bl[124] br[124] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_127 
+ bl[125] br[125] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_128 
+ bl[126] br[126] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_129 
+ bl[127] br[127] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_130 
+ bl[128] br[128] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_131 
+ bl[129] br[129] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_132 
+ bl[130] br[130] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_133 
+ bl[131] br[131] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_134 
+ bl[132] br[132] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_135 
+ bl[133] br[133] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_136 
+ bl[134] br[134] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_137 
+ bl[135] br[135] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_138 
+ bl[136] br[136] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_139 
+ bl[137] br[137] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_140 
+ bl[138] br[138] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_141 
+ bl[139] br[139] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_142 
+ bl[140] br[140] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_143 
+ bl[141] br[141] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_144 
+ bl[142] br[142] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_145 
+ bl[143] br[143] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_146 
+ bl[144] br[144] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_147 
+ bl[145] br[145] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_148 
+ bl[146] br[146] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_149 
+ bl[147] br[147] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_150 
+ bl[148] br[148] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_151 
+ bl[149] br[149] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_152 
+ bl[150] br[150] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_153 
+ bl[151] br[151] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_154 
+ bl[152] br[152] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_155 
+ bl[153] br[153] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_156 
+ bl[154] br[154] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_157 
+ bl[155] br[155] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_158 
+ bl[156] br[156] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_159 
+ bl[157] br[157] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_160 
+ bl[158] br[158] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_161 
+ bl[159] br[159] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_162 
+ bl[160] br[160] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_163 
+ bl[161] br[161] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_164 
+ bl[162] br[162] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_165 
+ bl[163] br[163] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_166 
+ bl[164] br[164] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_167 
+ bl[165] br[165] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_168 
+ bl[166] br[166] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_169 
+ bl[167] br[167] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_170 
+ bl[168] br[168] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_171 
+ bl[169] br[169] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_172 
+ bl[170] br[170] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_173 
+ bl[171] br[171] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_174 
+ bl[172] br[172] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_175 
+ bl[173] br[173] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_176 
+ bl[174] br[174] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_177 
+ bl[175] br[175] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_178 
+ bl[176] br[176] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_179 
+ bl[177] br[177] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_180 
+ bl[178] br[178] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_181 
+ bl[179] br[179] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_182 
+ bl[180] br[180] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_183 
+ bl[181] br[181] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_184 
+ bl[182] br[182] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_185 
+ bl[183] br[183] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_186 
+ bl[184] br[184] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_187 
+ bl[185] br[185] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_188 
+ bl[186] br[186] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_189 
+ bl[187] br[187] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_190 
+ bl[188] br[188] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_191 
+ bl[189] br[189] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_192 
+ bl[190] br[190] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_193 
+ bl[191] br[191] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_194 
+ bl[192] br[192] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_195 
+ bl[193] br[193] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_196 
+ bl[194] br[194] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_197 
+ bl[195] br[195] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_198 
+ bl[196] br[196] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_199 
+ bl[197] br[197] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_200 
+ bl[198] br[198] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_201 
+ bl[199] br[199] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_202 
+ bl[200] br[200] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_203 
+ bl[201] br[201] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_204 
+ bl[202] br[202] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_205 
+ bl[203] br[203] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_206 
+ bl[204] br[204] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_207 
+ bl[205] br[205] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_208 
+ bl[206] br[206] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_209 
+ bl[207] br[207] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_210 
+ bl[208] br[208] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_211 
+ bl[209] br[209] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_212 
+ bl[210] br[210] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_213 
+ bl[211] br[211] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_214 
+ bl[212] br[212] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_215 
+ bl[213] br[213] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_216 
+ bl[214] br[214] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_217 
+ bl[215] br[215] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_218 
+ bl[216] br[216] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_219 
+ bl[217] br[217] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_220 
+ bl[218] br[218] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_221 
+ bl[219] br[219] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_222 
+ bl[220] br[220] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_223 
+ bl[221] br[221] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_224 
+ bl[222] br[222] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_225 
+ bl[223] br[223] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_226 
+ bl[224] br[224] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_227 
+ bl[225] br[225] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_228 
+ bl[226] br[226] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_229 
+ bl[227] br[227] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_230 
+ bl[228] br[228] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_231 
+ bl[229] br[229] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_232 
+ bl[230] br[230] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_233 
+ bl[231] br[231] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_234 
+ bl[232] br[232] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_235 
+ bl[233] br[233] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_236 
+ bl[234] br[234] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_237 
+ bl[235] br[235] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_238 
+ bl[236] br[236] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_239 
+ bl[237] br[237] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_240 
+ bl[238] br[238] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_241 
+ bl[239] br[239] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_242 
+ bl[240] br[240] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_243 
+ bl[241] br[241] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_244 
+ bl[242] br[242] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_245 
+ bl[243] br[243] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_246 
+ bl[244] br[244] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_247 
+ bl[245] br[245] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_248 
+ bl[246] br[246] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_249 
+ bl[247] br[247] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_250 
+ bl[248] br[248] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_251 
+ bl[249] br[249] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_252 
+ bl[250] br[250] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_253 
+ bl[251] br[251] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_254 
+ bl[252] br[252] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_255 
+ bl[253] br[253] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_256 
+ bl[254] br[254] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_257 
+ bl[255] br[255] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_258 
+ vdd vdd vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_259 
+ vdd vdd vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_0 
+ vdd vdd vss vdd vpb vnb wl[102] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_104_1 
+ rbl rbr vss vdd vpb vnb wl[102] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_104_2 
+ bl[0] br[0] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_3 
+ bl[1] br[1] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_4 
+ bl[2] br[2] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_5 
+ bl[3] br[3] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_6 
+ bl[4] br[4] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_7 
+ bl[5] br[5] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_8 
+ bl[6] br[6] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_9 
+ bl[7] br[7] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_10 
+ bl[8] br[8] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_11 
+ bl[9] br[9] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_12 
+ bl[10] br[10] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_13 
+ bl[11] br[11] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_14 
+ bl[12] br[12] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_15 
+ bl[13] br[13] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_16 
+ bl[14] br[14] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_17 
+ bl[15] br[15] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_18 
+ bl[16] br[16] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_19 
+ bl[17] br[17] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_20 
+ bl[18] br[18] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_21 
+ bl[19] br[19] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_22 
+ bl[20] br[20] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_23 
+ bl[21] br[21] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_24 
+ bl[22] br[22] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_25 
+ bl[23] br[23] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_26 
+ bl[24] br[24] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_27 
+ bl[25] br[25] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_28 
+ bl[26] br[26] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_29 
+ bl[27] br[27] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_30 
+ bl[28] br[28] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_31 
+ bl[29] br[29] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_32 
+ bl[30] br[30] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_33 
+ bl[31] br[31] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_34 
+ bl[32] br[32] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_35 
+ bl[33] br[33] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_36 
+ bl[34] br[34] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_37 
+ bl[35] br[35] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_38 
+ bl[36] br[36] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_39 
+ bl[37] br[37] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_40 
+ bl[38] br[38] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_41 
+ bl[39] br[39] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_42 
+ bl[40] br[40] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_43 
+ bl[41] br[41] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_44 
+ bl[42] br[42] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_45 
+ bl[43] br[43] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_46 
+ bl[44] br[44] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_47 
+ bl[45] br[45] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_48 
+ bl[46] br[46] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_49 
+ bl[47] br[47] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_50 
+ bl[48] br[48] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_51 
+ bl[49] br[49] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_52 
+ bl[50] br[50] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_53 
+ bl[51] br[51] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_54 
+ bl[52] br[52] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_55 
+ bl[53] br[53] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_56 
+ bl[54] br[54] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_57 
+ bl[55] br[55] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_58 
+ bl[56] br[56] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_59 
+ bl[57] br[57] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_60 
+ bl[58] br[58] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_61 
+ bl[59] br[59] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_62 
+ bl[60] br[60] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_63 
+ bl[61] br[61] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_64 
+ bl[62] br[62] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_65 
+ bl[63] br[63] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_66 
+ bl[64] br[64] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_67 
+ bl[65] br[65] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_68 
+ bl[66] br[66] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_69 
+ bl[67] br[67] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_70 
+ bl[68] br[68] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_71 
+ bl[69] br[69] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_72 
+ bl[70] br[70] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_73 
+ bl[71] br[71] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_74 
+ bl[72] br[72] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_75 
+ bl[73] br[73] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_76 
+ bl[74] br[74] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_77 
+ bl[75] br[75] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_78 
+ bl[76] br[76] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_79 
+ bl[77] br[77] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_80 
+ bl[78] br[78] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_81 
+ bl[79] br[79] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_82 
+ bl[80] br[80] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_83 
+ bl[81] br[81] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_84 
+ bl[82] br[82] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_85 
+ bl[83] br[83] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_86 
+ bl[84] br[84] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_87 
+ bl[85] br[85] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_88 
+ bl[86] br[86] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_89 
+ bl[87] br[87] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_90 
+ bl[88] br[88] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_91 
+ bl[89] br[89] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_92 
+ bl[90] br[90] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_93 
+ bl[91] br[91] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_94 
+ bl[92] br[92] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_95 
+ bl[93] br[93] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_96 
+ bl[94] br[94] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_97 
+ bl[95] br[95] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_98 
+ bl[96] br[96] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_99 
+ bl[97] br[97] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_100 
+ bl[98] br[98] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_101 
+ bl[99] br[99] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_102 
+ bl[100] br[100] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_103 
+ bl[101] br[101] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_104 
+ bl[102] br[102] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_105 
+ bl[103] br[103] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_106 
+ bl[104] br[104] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_107 
+ bl[105] br[105] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_108 
+ bl[106] br[106] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_109 
+ bl[107] br[107] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_110 
+ bl[108] br[108] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_111 
+ bl[109] br[109] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_112 
+ bl[110] br[110] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_113 
+ bl[111] br[111] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_114 
+ bl[112] br[112] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_115 
+ bl[113] br[113] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_116 
+ bl[114] br[114] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_117 
+ bl[115] br[115] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_118 
+ bl[116] br[116] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_119 
+ bl[117] br[117] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_120 
+ bl[118] br[118] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_121 
+ bl[119] br[119] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_122 
+ bl[120] br[120] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_123 
+ bl[121] br[121] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_124 
+ bl[122] br[122] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_125 
+ bl[123] br[123] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_126 
+ bl[124] br[124] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_127 
+ bl[125] br[125] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_128 
+ bl[126] br[126] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_129 
+ bl[127] br[127] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_130 
+ bl[128] br[128] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_131 
+ bl[129] br[129] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_132 
+ bl[130] br[130] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_133 
+ bl[131] br[131] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_134 
+ bl[132] br[132] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_135 
+ bl[133] br[133] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_136 
+ bl[134] br[134] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_137 
+ bl[135] br[135] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_138 
+ bl[136] br[136] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_139 
+ bl[137] br[137] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_140 
+ bl[138] br[138] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_141 
+ bl[139] br[139] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_142 
+ bl[140] br[140] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_143 
+ bl[141] br[141] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_144 
+ bl[142] br[142] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_145 
+ bl[143] br[143] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_146 
+ bl[144] br[144] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_147 
+ bl[145] br[145] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_148 
+ bl[146] br[146] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_149 
+ bl[147] br[147] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_150 
+ bl[148] br[148] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_151 
+ bl[149] br[149] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_152 
+ bl[150] br[150] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_153 
+ bl[151] br[151] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_154 
+ bl[152] br[152] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_155 
+ bl[153] br[153] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_156 
+ bl[154] br[154] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_157 
+ bl[155] br[155] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_158 
+ bl[156] br[156] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_159 
+ bl[157] br[157] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_160 
+ bl[158] br[158] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_161 
+ bl[159] br[159] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_162 
+ bl[160] br[160] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_163 
+ bl[161] br[161] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_164 
+ bl[162] br[162] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_165 
+ bl[163] br[163] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_166 
+ bl[164] br[164] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_167 
+ bl[165] br[165] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_168 
+ bl[166] br[166] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_169 
+ bl[167] br[167] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_170 
+ bl[168] br[168] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_171 
+ bl[169] br[169] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_172 
+ bl[170] br[170] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_173 
+ bl[171] br[171] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_174 
+ bl[172] br[172] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_175 
+ bl[173] br[173] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_176 
+ bl[174] br[174] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_177 
+ bl[175] br[175] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_178 
+ bl[176] br[176] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_179 
+ bl[177] br[177] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_180 
+ bl[178] br[178] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_181 
+ bl[179] br[179] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_182 
+ bl[180] br[180] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_183 
+ bl[181] br[181] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_184 
+ bl[182] br[182] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_185 
+ bl[183] br[183] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_186 
+ bl[184] br[184] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_187 
+ bl[185] br[185] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_188 
+ bl[186] br[186] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_189 
+ bl[187] br[187] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_190 
+ bl[188] br[188] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_191 
+ bl[189] br[189] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_192 
+ bl[190] br[190] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_193 
+ bl[191] br[191] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_194 
+ bl[192] br[192] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_195 
+ bl[193] br[193] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_196 
+ bl[194] br[194] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_197 
+ bl[195] br[195] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_198 
+ bl[196] br[196] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_199 
+ bl[197] br[197] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_200 
+ bl[198] br[198] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_201 
+ bl[199] br[199] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_202 
+ bl[200] br[200] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_203 
+ bl[201] br[201] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_204 
+ bl[202] br[202] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_205 
+ bl[203] br[203] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_206 
+ bl[204] br[204] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_207 
+ bl[205] br[205] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_208 
+ bl[206] br[206] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_209 
+ bl[207] br[207] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_210 
+ bl[208] br[208] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_211 
+ bl[209] br[209] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_212 
+ bl[210] br[210] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_213 
+ bl[211] br[211] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_214 
+ bl[212] br[212] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_215 
+ bl[213] br[213] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_216 
+ bl[214] br[214] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_217 
+ bl[215] br[215] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_218 
+ bl[216] br[216] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_219 
+ bl[217] br[217] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_220 
+ bl[218] br[218] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_221 
+ bl[219] br[219] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_222 
+ bl[220] br[220] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_223 
+ bl[221] br[221] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_224 
+ bl[222] br[222] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_225 
+ bl[223] br[223] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_226 
+ bl[224] br[224] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_227 
+ bl[225] br[225] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_228 
+ bl[226] br[226] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_229 
+ bl[227] br[227] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_230 
+ bl[228] br[228] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_231 
+ bl[229] br[229] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_232 
+ bl[230] br[230] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_233 
+ bl[231] br[231] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_234 
+ bl[232] br[232] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_235 
+ bl[233] br[233] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_236 
+ bl[234] br[234] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_237 
+ bl[235] br[235] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_238 
+ bl[236] br[236] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_239 
+ bl[237] br[237] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_240 
+ bl[238] br[238] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_241 
+ bl[239] br[239] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_242 
+ bl[240] br[240] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_243 
+ bl[241] br[241] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_244 
+ bl[242] br[242] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_245 
+ bl[243] br[243] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_246 
+ bl[244] br[244] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_247 
+ bl[245] br[245] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_248 
+ bl[246] br[246] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_249 
+ bl[247] br[247] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_250 
+ bl[248] br[248] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_251 
+ bl[249] br[249] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_252 
+ bl[250] br[250] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_253 
+ bl[251] br[251] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_254 
+ bl[252] br[252] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_255 
+ bl[253] br[253] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_256 
+ bl[254] br[254] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_257 
+ bl[255] br[255] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_258 
+ vdd vdd vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_259 
+ vdd vdd vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_0 
+ vdd vdd vss vdd vpb vnb wl[103] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_105_1 
+ rbl rbr vss vdd vpb vnb wl[103] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_105_2 
+ bl[0] br[0] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_3 
+ bl[1] br[1] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_4 
+ bl[2] br[2] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_5 
+ bl[3] br[3] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_6 
+ bl[4] br[4] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_7 
+ bl[5] br[5] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_8 
+ bl[6] br[6] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_9 
+ bl[7] br[7] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_10 
+ bl[8] br[8] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_11 
+ bl[9] br[9] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_12 
+ bl[10] br[10] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_13 
+ bl[11] br[11] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_14 
+ bl[12] br[12] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_15 
+ bl[13] br[13] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_16 
+ bl[14] br[14] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_17 
+ bl[15] br[15] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_18 
+ bl[16] br[16] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_19 
+ bl[17] br[17] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_20 
+ bl[18] br[18] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_21 
+ bl[19] br[19] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_22 
+ bl[20] br[20] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_23 
+ bl[21] br[21] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_24 
+ bl[22] br[22] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_25 
+ bl[23] br[23] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_26 
+ bl[24] br[24] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_27 
+ bl[25] br[25] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_28 
+ bl[26] br[26] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_29 
+ bl[27] br[27] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_30 
+ bl[28] br[28] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_31 
+ bl[29] br[29] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_32 
+ bl[30] br[30] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_33 
+ bl[31] br[31] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_34 
+ bl[32] br[32] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_35 
+ bl[33] br[33] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_36 
+ bl[34] br[34] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_37 
+ bl[35] br[35] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_38 
+ bl[36] br[36] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_39 
+ bl[37] br[37] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_40 
+ bl[38] br[38] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_41 
+ bl[39] br[39] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_42 
+ bl[40] br[40] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_43 
+ bl[41] br[41] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_44 
+ bl[42] br[42] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_45 
+ bl[43] br[43] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_46 
+ bl[44] br[44] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_47 
+ bl[45] br[45] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_48 
+ bl[46] br[46] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_49 
+ bl[47] br[47] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_50 
+ bl[48] br[48] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_51 
+ bl[49] br[49] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_52 
+ bl[50] br[50] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_53 
+ bl[51] br[51] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_54 
+ bl[52] br[52] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_55 
+ bl[53] br[53] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_56 
+ bl[54] br[54] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_57 
+ bl[55] br[55] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_58 
+ bl[56] br[56] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_59 
+ bl[57] br[57] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_60 
+ bl[58] br[58] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_61 
+ bl[59] br[59] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_62 
+ bl[60] br[60] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_63 
+ bl[61] br[61] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_64 
+ bl[62] br[62] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_65 
+ bl[63] br[63] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_66 
+ bl[64] br[64] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_67 
+ bl[65] br[65] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_68 
+ bl[66] br[66] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_69 
+ bl[67] br[67] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_70 
+ bl[68] br[68] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_71 
+ bl[69] br[69] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_72 
+ bl[70] br[70] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_73 
+ bl[71] br[71] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_74 
+ bl[72] br[72] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_75 
+ bl[73] br[73] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_76 
+ bl[74] br[74] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_77 
+ bl[75] br[75] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_78 
+ bl[76] br[76] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_79 
+ bl[77] br[77] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_80 
+ bl[78] br[78] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_81 
+ bl[79] br[79] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_82 
+ bl[80] br[80] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_83 
+ bl[81] br[81] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_84 
+ bl[82] br[82] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_85 
+ bl[83] br[83] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_86 
+ bl[84] br[84] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_87 
+ bl[85] br[85] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_88 
+ bl[86] br[86] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_89 
+ bl[87] br[87] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_90 
+ bl[88] br[88] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_91 
+ bl[89] br[89] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_92 
+ bl[90] br[90] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_93 
+ bl[91] br[91] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_94 
+ bl[92] br[92] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_95 
+ bl[93] br[93] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_96 
+ bl[94] br[94] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_97 
+ bl[95] br[95] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_98 
+ bl[96] br[96] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_99 
+ bl[97] br[97] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_100 
+ bl[98] br[98] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_101 
+ bl[99] br[99] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_102 
+ bl[100] br[100] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_103 
+ bl[101] br[101] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_104 
+ bl[102] br[102] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_105 
+ bl[103] br[103] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_106 
+ bl[104] br[104] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_107 
+ bl[105] br[105] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_108 
+ bl[106] br[106] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_109 
+ bl[107] br[107] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_110 
+ bl[108] br[108] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_111 
+ bl[109] br[109] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_112 
+ bl[110] br[110] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_113 
+ bl[111] br[111] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_114 
+ bl[112] br[112] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_115 
+ bl[113] br[113] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_116 
+ bl[114] br[114] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_117 
+ bl[115] br[115] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_118 
+ bl[116] br[116] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_119 
+ bl[117] br[117] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_120 
+ bl[118] br[118] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_121 
+ bl[119] br[119] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_122 
+ bl[120] br[120] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_123 
+ bl[121] br[121] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_124 
+ bl[122] br[122] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_125 
+ bl[123] br[123] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_126 
+ bl[124] br[124] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_127 
+ bl[125] br[125] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_128 
+ bl[126] br[126] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_129 
+ bl[127] br[127] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_130 
+ bl[128] br[128] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_131 
+ bl[129] br[129] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_132 
+ bl[130] br[130] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_133 
+ bl[131] br[131] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_134 
+ bl[132] br[132] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_135 
+ bl[133] br[133] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_136 
+ bl[134] br[134] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_137 
+ bl[135] br[135] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_138 
+ bl[136] br[136] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_139 
+ bl[137] br[137] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_140 
+ bl[138] br[138] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_141 
+ bl[139] br[139] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_142 
+ bl[140] br[140] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_143 
+ bl[141] br[141] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_144 
+ bl[142] br[142] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_145 
+ bl[143] br[143] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_146 
+ bl[144] br[144] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_147 
+ bl[145] br[145] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_148 
+ bl[146] br[146] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_149 
+ bl[147] br[147] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_150 
+ bl[148] br[148] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_151 
+ bl[149] br[149] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_152 
+ bl[150] br[150] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_153 
+ bl[151] br[151] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_154 
+ bl[152] br[152] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_155 
+ bl[153] br[153] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_156 
+ bl[154] br[154] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_157 
+ bl[155] br[155] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_158 
+ bl[156] br[156] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_159 
+ bl[157] br[157] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_160 
+ bl[158] br[158] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_161 
+ bl[159] br[159] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_162 
+ bl[160] br[160] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_163 
+ bl[161] br[161] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_164 
+ bl[162] br[162] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_165 
+ bl[163] br[163] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_166 
+ bl[164] br[164] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_167 
+ bl[165] br[165] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_168 
+ bl[166] br[166] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_169 
+ bl[167] br[167] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_170 
+ bl[168] br[168] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_171 
+ bl[169] br[169] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_172 
+ bl[170] br[170] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_173 
+ bl[171] br[171] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_174 
+ bl[172] br[172] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_175 
+ bl[173] br[173] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_176 
+ bl[174] br[174] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_177 
+ bl[175] br[175] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_178 
+ bl[176] br[176] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_179 
+ bl[177] br[177] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_180 
+ bl[178] br[178] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_181 
+ bl[179] br[179] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_182 
+ bl[180] br[180] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_183 
+ bl[181] br[181] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_184 
+ bl[182] br[182] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_185 
+ bl[183] br[183] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_186 
+ bl[184] br[184] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_187 
+ bl[185] br[185] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_188 
+ bl[186] br[186] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_189 
+ bl[187] br[187] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_190 
+ bl[188] br[188] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_191 
+ bl[189] br[189] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_192 
+ bl[190] br[190] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_193 
+ bl[191] br[191] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_194 
+ bl[192] br[192] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_195 
+ bl[193] br[193] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_196 
+ bl[194] br[194] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_197 
+ bl[195] br[195] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_198 
+ bl[196] br[196] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_199 
+ bl[197] br[197] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_200 
+ bl[198] br[198] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_201 
+ bl[199] br[199] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_202 
+ bl[200] br[200] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_203 
+ bl[201] br[201] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_204 
+ bl[202] br[202] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_205 
+ bl[203] br[203] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_206 
+ bl[204] br[204] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_207 
+ bl[205] br[205] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_208 
+ bl[206] br[206] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_209 
+ bl[207] br[207] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_210 
+ bl[208] br[208] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_211 
+ bl[209] br[209] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_212 
+ bl[210] br[210] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_213 
+ bl[211] br[211] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_214 
+ bl[212] br[212] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_215 
+ bl[213] br[213] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_216 
+ bl[214] br[214] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_217 
+ bl[215] br[215] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_218 
+ bl[216] br[216] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_219 
+ bl[217] br[217] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_220 
+ bl[218] br[218] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_221 
+ bl[219] br[219] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_222 
+ bl[220] br[220] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_223 
+ bl[221] br[221] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_224 
+ bl[222] br[222] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_225 
+ bl[223] br[223] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_226 
+ bl[224] br[224] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_227 
+ bl[225] br[225] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_228 
+ bl[226] br[226] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_229 
+ bl[227] br[227] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_230 
+ bl[228] br[228] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_231 
+ bl[229] br[229] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_232 
+ bl[230] br[230] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_233 
+ bl[231] br[231] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_234 
+ bl[232] br[232] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_235 
+ bl[233] br[233] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_236 
+ bl[234] br[234] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_237 
+ bl[235] br[235] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_238 
+ bl[236] br[236] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_239 
+ bl[237] br[237] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_240 
+ bl[238] br[238] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_241 
+ bl[239] br[239] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_242 
+ bl[240] br[240] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_243 
+ bl[241] br[241] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_244 
+ bl[242] br[242] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_245 
+ bl[243] br[243] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_246 
+ bl[244] br[244] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_247 
+ bl[245] br[245] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_248 
+ bl[246] br[246] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_249 
+ bl[247] br[247] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_250 
+ bl[248] br[248] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_251 
+ bl[249] br[249] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_252 
+ bl[250] br[250] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_253 
+ bl[251] br[251] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_254 
+ bl[252] br[252] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_255 
+ bl[253] br[253] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_256 
+ bl[254] br[254] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_257 
+ bl[255] br[255] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_258 
+ vdd vdd vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_259 
+ vdd vdd vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_0 
+ vdd vdd vss vdd vpb vnb wl[104] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_106_1 
+ rbl rbr vss vdd vpb vnb wl[104] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_106_2 
+ bl[0] br[0] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_3 
+ bl[1] br[1] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_4 
+ bl[2] br[2] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_5 
+ bl[3] br[3] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_6 
+ bl[4] br[4] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_7 
+ bl[5] br[5] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_8 
+ bl[6] br[6] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_9 
+ bl[7] br[7] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_10 
+ bl[8] br[8] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_11 
+ bl[9] br[9] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_12 
+ bl[10] br[10] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_13 
+ bl[11] br[11] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_14 
+ bl[12] br[12] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_15 
+ bl[13] br[13] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_16 
+ bl[14] br[14] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_17 
+ bl[15] br[15] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_18 
+ bl[16] br[16] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_19 
+ bl[17] br[17] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_20 
+ bl[18] br[18] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_21 
+ bl[19] br[19] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_22 
+ bl[20] br[20] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_23 
+ bl[21] br[21] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_24 
+ bl[22] br[22] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_25 
+ bl[23] br[23] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_26 
+ bl[24] br[24] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_27 
+ bl[25] br[25] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_28 
+ bl[26] br[26] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_29 
+ bl[27] br[27] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_30 
+ bl[28] br[28] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_31 
+ bl[29] br[29] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_32 
+ bl[30] br[30] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_33 
+ bl[31] br[31] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_34 
+ bl[32] br[32] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_35 
+ bl[33] br[33] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_36 
+ bl[34] br[34] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_37 
+ bl[35] br[35] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_38 
+ bl[36] br[36] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_39 
+ bl[37] br[37] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_40 
+ bl[38] br[38] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_41 
+ bl[39] br[39] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_42 
+ bl[40] br[40] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_43 
+ bl[41] br[41] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_44 
+ bl[42] br[42] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_45 
+ bl[43] br[43] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_46 
+ bl[44] br[44] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_47 
+ bl[45] br[45] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_48 
+ bl[46] br[46] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_49 
+ bl[47] br[47] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_50 
+ bl[48] br[48] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_51 
+ bl[49] br[49] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_52 
+ bl[50] br[50] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_53 
+ bl[51] br[51] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_54 
+ bl[52] br[52] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_55 
+ bl[53] br[53] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_56 
+ bl[54] br[54] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_57 
+ bl[55] br[55] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_58 
+ bl[56] br[56] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_59 
+ bl[57] br[57] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_60 
+ bl[58] br[58] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_61 
+ bl[59] br[59] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_62 
+ bl[60] br[60] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_63 
+ bl[61] br[61] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_64 
+ bl[62] br[62] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_65 
+ bl[63] br[63] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_66 
+ bl[64] br[64] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_67 
+ bl[65] br[65] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_68 
+ bl[66] br[66] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_69 
+ bl[67] br[67] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_70 
+ bl[68] br[68] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_71 
+ bl[69] br[69] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_72 
+ bl[70] br[70] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_73 
+ bl[71] br[71] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_74 
+ bl[72] br[72] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_75 
+ bl[73] br[73] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_76 
+ bl[74] br[74] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_77 
+ bl[75] br[75] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_78 
+ bl[76] br[76] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_79 
+ bl[77] br[77] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_80 
+ bl[78] br[78] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_81 
+ bl[79] br[79] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_82 
+ bl[80] br[80] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_83 
+ bl[81] br[81] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_84 
+ bl[82] br[82] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_85 
+ bl[83] br[83] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_86 
+ bl[84] br[84] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_87 
+ bl[85] br[85] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_88 
+ bl[86] br[86] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_89 
+ bl[87] br[87] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_90 
+ bl[88] br[88] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_91 
+ bl[89] br[89] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_92 
+ bl[90] br[90] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_93 
+ bl[91] br[91] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_94 
+ bl[92] br[92] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_95 
+ bl[93] br[93] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_96 
+ bl[94] br[94] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_97 
+ bl[95] br[95] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_98 
+ bl[96] br[96] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_99 
+ bl[97] br[97] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_100 
+ bl[98] br[98] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_101 
+ bl[99] br[99] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_102 
+ bl[100] br[100] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_103 
+ bl[101] br[101] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_104 
+ bl[102] br[102] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_105 
+ bl[103] br[103] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_106 
+ bl[104] br[104] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_107 
+ bl[105] br[105] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_108 
+ bl[106] br[106] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_109 
+ bl[107] br[107] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_110 
+ bl[108] br[108] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_111 
+ bl[109] br[109] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_112 
+ bl[110] br[110] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_113 
+ bl[111] br[111] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_114 
+ bl[112] br[112] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_115 
+ bl[113] br[113] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_116 
+ bl[114] br[114] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_117 
+ bl[115] br[115] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_118 
+ bl[116] br[116] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_119 
+ bl[117] br[117] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_120 
+ bl[118] br[118] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_121 
+ bl[119] br[119] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_122 
+ bl[120] br[120] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_123 
+ bl[121] br[121] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_124 
+ bl[122] br[122] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_125 
+ bl[123] br[123] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_126 
+ bl[124] br[124] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_127 
+ bl[125] br[125] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_128 
+ bl[126] br[126] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_129 
+ bl[127] br[127] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_130 
+ bl[128] br[128] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_131 
+ bl[129] br[129] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_132 
+ bl[130] br[130] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_133 
+ bl[131] br[131] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_134 
+ bl[132] br[132] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_135 
+ bl[133] br[133] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_136 
+ bl[134] br[134] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_137 
+ bl[135] br[135] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_138 
+ bl[136] br[136] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_139 
+ bl[137] br[137] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_140 
+ bl[138] br[138] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_141 
+ bl[139] br[139] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_142 
+ bl[140] br[140] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_143 
+ bl[141] br[141] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_144 
+ bl[142] br[142] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_145 
+ bl[143] br[143] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_146 
+ bl[144] br[144] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_147 
+ bl[145] br[145] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_148 
+ bl[146] br[146] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_149 
+ bl[147] br[147] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_150 
+ bl[148] br[148] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_151 
+ bl[149] br[149] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_152 
+ bl[150] br[150] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_153 
+ bl[151] br[151] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_154 
+ bl[152] br[152] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_155 
+ bl[153] br[153] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_156 
+ bl[154] br[154] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_157 
+ bl[155] br[155] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_158 
+ bl[156] br[156] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_159 
+ bl[157] br[157] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_160 
+ bl[158] br[158] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_161 
+ bl[159] br[159] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_162 
+ bl[160] br[160] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_163 
+ bl[161] br[161] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_164 
+ bl[162] br[162] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_165 
+ bl[163] br[163] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_166 
+ bl[164] br[164] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_167 
+ bl[165] br[165] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_168 
+ bl[166] br[166] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_169 
+ bl[167] br[167] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_170 
+ bl[168] br[168] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_171 
+ bl[169] br[169] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_172 
+ bl[170] br[170] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_173 
+ bl[171] br[171] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_174 
+ bl[172] br[172] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_175 
+ bl[173] br[173] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_176 
+ bl[174] br[174] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_177 
+ bl[175] br[175] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_178 
+ bl[176] br[176] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_179 
+ bl[177] br[177] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_180 
+ bl[178] br[178] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_181 
+ bl[179] br[179] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_182 
+ bl[180] br[180] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_183 
+ bl[181] br[181] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_184 
+ bl[182] br[182] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_185 
+ bl[183] br[183] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_186 
+ bl[184] br[184] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_187 
+ bl[185] br[185] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_188 
+ bl[186] br[186] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_189 
+ bl[187] br[187] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_190 
+ bl[188] br[188] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_191 
+ bl[189] br[189] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_192 
+ bl[190] br[190] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_193 
+ bl[191] br[191] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_194 
+ bl[192] br[192] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_195 
+ bl[193] br[193] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_196 
+ bl[194] br[194] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_197 
+ bl[195] br[195] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_198 
+ bl[196] br[196] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_199 
+ bl[197] br[197] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_200 
+ bl[198] br[198] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_201 
+ bl[199] br[199] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_202 
+ bl[200] br[200] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_203 
+ bl[201] br[201] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_204 
+ bl[202] br[202] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_205 
+ bl[203] br[203] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_206 
+ bl[204] br[204] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_207 
+ bl[205] br[205] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_208 
+ bl[206] br[206] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_209 
+ bl[207] br[207] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_210 
+ bl[208] br[208] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_211 
+ bl[209] br[209] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_212 
+ bl[210] br[210] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_213 
+ bl[211] br[211] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_214 
+ bl[212] br[212] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_215 
+ bl[213] br[213] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_216 
+ bl[214] br[214] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_217 
+ bl[215] br[215] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_218 
+ bl[216] br[216] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_219 
+ bl[217] br[217] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_220 
+ bl[218] br[218] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_221 
+ bl[219] br[219] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_222 
+ bl[220] br[220] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_223 
+ bl[221] br[221] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_224 
+ bl[222] br[222] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_225 
+ bl[223] br[223] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_226 
+ bl[224] br[224] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_227 
+ bl[225] br[225] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_228 
+ bl[226] br[226] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_229 
+ bl[227] br[227] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_230 
+ bl[228] br[228] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_231 
+ bl[229] br[229] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_232 
+ bl[230] br[230] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_233 
+ bl[231] br[231] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_234 
+ bl[232] br[232] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_235 
+ bl[233] br[233] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_236 
+ bl[234] br[234] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_237 
+ bl[235] br[235] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_238 
+ bl[236] br[236] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_239 
+ bl[237] br[237] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_240 
+ bl[238] br[238] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_241 
+ bl[239] br[239] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_242 
+ bl[240] br[240] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_243 
+ bl[241] br[241] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_244 
+ bl[242] br[242] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_245 
+ bl[243] br[243] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_246 
+ bl[244] br[244] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_247 
+ bl[245] br[245] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_248 
+ bl[246] br[246] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_249 
+ bl[247] br[247] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_250 
+ bl[248] br[248] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_251 
+ bl[249] br[249] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_252 
+ bl[250] br[250] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_253 
+ bl[251] br[251] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_254 
+ bl[252] br[252] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_255 
+ bl[253] br[253] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_256 
+ bl[254] br[254] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_257 
+ bl[255] br[255] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_258 
+ vdd vdd vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_259 
+ vdd vdd vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_0 
+ vdd vdd vss vdd vpb vnb wl[105] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_107_1 
+ rbl rbr vss vdd vpb vnb wl[105] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_107_2 
+ bl[0] br[0] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_3 
+ bl[1] br[1] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_4 
+ bl[2] br[2] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_5 
+ bl[3] br[3] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_6 
+ bl[4] br[4] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_7 
+ bl[5] br[5] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_8 
+ bl[6] br[6] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_9 
+ bl[7] br[7] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_10 
+ bl[8] br[8] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_11 
+ bl[9] br[9] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_12 
+ bl[10] br[10] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_13 
+ bl[11] br[11] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_14 
+ bl[12] br[12] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_15 
+ bl[13] br[13] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_16 
+ bl[14] br[14] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_17 
+ bl[15] br[15] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_18 
+ bl[16] br[16] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_19 
+ bl[17] br[17] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_20 
+ bl[18] br[18] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_21 
+ bl[19] br[19] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_22 
+ bl[20] br[20] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_23 
+ bl[21] br[21] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_24 
+ bl[22] br[22] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_25 
+ bl[23] br[23] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_26 
+ bl[24] br[24] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_27 
+ bl[25] br[25] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_28 
+ bl[26] br[26] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_29 
+ bl[27] br[27] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_30 
+ bl[28] br[28] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_31 
+ bl[29] br[29] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_32 
+ bl[30] br[30] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_33 
+ bl[31] br[31] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_34 
+ bl[32] br[32] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_35 
+ bl[33] br[33] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_36 
+ bl[34] br[34] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_37 
+ bl[35] br[35] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_38 
+ bl[36] br[36] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_39 
+ bl[37] br[37] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_40 
+ bl[38] br[38] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_41 
+ bl[39] br[39] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_42 
+ bl[40] br[40] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_43 
+ bl[41] br[41] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_44 
+ bl[42] br[42] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_45 
+ bl[43] br[43] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_46 
+ bl[44] br[44] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_47 
+ bl[45] br[45] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_48 
+ bl[46] br[46] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_49 
+ bl[47] br[47] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_50 
+ bl[48] br[48] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_51 
+ bl[49] br[49] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_52 
+ bl[50] br[50] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_53 
+ bl[51] br[51] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_54 
+ bl[52] br[52] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_55 
+ bl[53] br[53] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_56 
+ bl[54] br[54] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_57 
+ bl[55] br[55] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_58 
+ bl[56] br[56] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_59 
+ bl[57] br[57] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_60 
+ bl[58] br[58] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_61 
+ bl[59] br[59] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_62 
+ bl[60] br[60] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_63 
+ bl[61] br[61] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_64 
+ bl[62] br[62] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_65 
+ bl[63] br[63] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_66 
+ bl[64] br[64] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_67 
+ bl[65] br[65] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_68 
+ bl[66] br[66] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_69 
+ bl[67] br[67] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_70 
+ bl[68] br[68] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_71 
+ bl[69] br[69] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_72 
+ bl[70] br[70] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_73 
+ bl[71] br[71] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_74 
+ bl[72] br[72] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_75 
+ bl[73] br[73] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_76 
+ bl[74] br[74] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_77 
+ bl[75] br[75] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_78 
+ bl[76] br[76] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_79 
+ bl[77] br[77] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_80 
+ bl[78] br[78] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_81 
+ bl[79] br[79] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_82 
+ bl[80] br[80] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_83 
+ bl[81] br[81] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_84 
+ bl[82] br[82] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_85 
+ bl[83] br[83] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_86 
+ bl[84] br[84] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_87 
+ bl[85] br[85] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_88 
+ bl[86] br[86] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_89 
+ bl[87] br[87] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_90 
+ bl[88] br[88] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_91 
+ bl[89] br[89] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_92 
+ bl[90] br[90] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_93 
+ bl[91] br[91] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_94 
+ bl[92] br[92] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_95 
+ bl[93] br[93] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_96 
+ bl[94] br[94] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_97 
+ bl[95] br[95] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_98 
+ bl[96] br[96] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_99 
+ bl[97] br[97] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_100 
+ bl[98] br[98] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_101 
+ bl[99] br[99] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_102 
+ bl[100] br[100] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_103 
+ bl[101] br[101] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_104 
+ bl[102] br[102] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_105 
+ bl[103] br[103] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_106 
+ bl[104] br[104] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_107 
+ bl[105] br[105] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_108 
+ bl[106] br[106] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_109 
+ bl[107] br[107] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_110 
+ bl[108] br[108] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_111 
+ bl[109] br[109] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_112 
+ bl[110] br[110] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_113 
+ bl[111] br[111] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_114 
+ bl[112] br[112] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_115 
+ bl[113] br[113] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_116 
+ bl[114] br[114] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_117 
+ bl[115] br[115] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_118 
+ bl[116] br[116] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_119 
+ bl[117] br[117] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_120 
+ bl[118] br[118] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_121 
+ bl[119] br[119] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_122 
+ bl[120] br[120] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_123 
+ bl[121] br[121] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_124 
+ bl[122] br[122] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_125 
+ bl[123] br[123] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_126 
+ bl[124] br[124] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_127 
+ bl[125] br[125] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_128 
+ bl[126] br[126] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_129 
+ bl[127] br[127] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_130 
+ bl[128] br[128] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_131 
+ bl[129] br[129] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_132 
+ bl[130] br[130] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_133 
+ bl[131] br[131] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_134 
+ bl[132] br[132] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_135 
+ bl[133] br[133] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_136 
+ bl[134] br[134] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_137 
+ bl[135] br[135] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_138 
+ bl[136] br[136] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_139 
+ bl[137] br[137] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_140 
+ bl[138] br[138] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_141 
+ bl[139] br[139] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_142 
+ bl[140] br[140] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_143 
+ bl[141] br[141] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_144 
+ bl[142] br[142] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_145 
+ bl[143] br[143] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_146 
+ bl[144] br[144] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_147 
+ bl[145] br[145] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_148 
+ bl[146] br[146] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_149 
+ bl[147] br[147] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_150 
+ bl[148] br[148] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_151 
+ bl[149] br[149] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_152 
+ bl[150] br[150] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_153 
+ bl[151] br[151] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_154 
+ bl[152] br[152] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_155 
+ bl[153] br[153] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_156 
+ bl[154] br[154] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_157 
+ bl[155] br[155] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_158 
+ bl[156] br[156] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_159 
+ bl[157] br[157] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_160 
+ bl[158] br[158] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_161 
+ bl[159] br[159] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_162 
+ bl[160] br[160] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_163 
+ bl[161] br[161] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_164 
+ bl[162] br[162] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_165 
+ bl[163] br[163] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_166 
+ bl[164] br[164] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_167 
+ bl[165] br[165] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_168 
+ bl[166] br[166] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_169 
+ bl[167] br[167] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_170 
+ bl[168] br[168] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_171 
+ bl[169] br[169] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_172 
+ bl[170] br[170] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_173 
+ bl[171] br[171] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_174 
+ bl[172] br[172] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_175 
+ bl[173] br[173] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_176 
+ bl[174] br[174] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_177 
+ bl[175] br[175] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_178 
+ bl[176] br[176] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_179 
+ bl[177] br[177] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_180 
+ bl[178] br[178] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_181 
+ bl[179] br[179] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_182 
+ bl[180] br[180] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_183 
+ bl[181] br[181] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_184 
+ bl[182] br[182] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_185 
+ bl[183] br[183] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_186 
+ bl[184] br[184] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_187 
+ bl[185] br[185] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_188 
+ bl[186] br[186] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_189 
+ bl[187] br[187] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_190 
+ bl[188] br[188] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_191 
+ bl[189] br[189] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_192 
+ bl[190] br[190] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_193 
+ bl[191] br[191] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_194 
+ bl[192] br[192] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_195 
+ bl[193] br[193] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_196 
+ bl[194] br[194] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_197 
+ bl[195] br[195] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_198 
+ bl[196] br[196] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_199 
+ bl[197] br[197] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_200 
+ bl[198] br[198] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_201 
+ bl[199] br[199] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_202 
+ bl[200] br[200] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_203 
+ bl[201] br[201] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_204 
+ bl[202] br[202] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_205 
+ bl[203] br[203] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_206 
+ bl[204] br[204] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_207 
+ bl[205] br[205] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_208 
+ bl[206] br[206] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_209 
+ bl[207] br[207] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_210 
+ bl[208] br[208] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_211 
+ bl[209] br[209] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_212 
+ bl[210] br[210] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_213 
+ bl[211] br[211] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_214 
+ bl[212] br[212] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_215 
+ bl[213] br[213] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_216 
+ bl[214] br[214] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_217 
+ bl[215] br[215] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_218 
+ bl[216] br[216] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_219 
+ bl[217] br[217] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_220 
+ bl[218] br[218] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_221 
+ bl[219] br[219] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_222 
+ bl[220] br[220] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_223 
+ bl[221] br[221] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_224 
+ bl[222] br[222] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_225 
+ bl[223] br[223] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_226 
+ bl[224] br[224] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_227 
+ bl[225] br[225] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_228 
+ bl[226] br[226] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_229 
+ bl[227] br[227] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_230 
+ bl[228] br[228] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_231 
+ bl[229] br[229] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_232 
+ bl[230] br[230] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_233 
+ bl[231] br[231] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_234 
+ bl[232] br[232] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_235 
+ bl[233] br[233] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_236 
+ bl[234] br[234] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_237 
+ bl[235] br[235] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_238 
+ bl[236] br[236] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_239 
+ bl[237] br[237] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_240 
+ bl[238] br[238] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_241 
+ bl[239] br[239] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_242 
+ bl[240] br[240] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_243 
+ bl[241] br[241] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_244 
+ bl[242] br[242] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_245 
+ bl[243] br[243] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_246 
+ bl[244] br[244] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_247 
+ bl[245] br[245] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_248 
+ bl[246] br[246] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_249 
+ bl[247] br[247] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_250 
+ bl[248] br[248] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_251 
+ bl[249] br[249] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_252 
+ bl[250] br[250] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_253 
+ bl[251] br[251] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_254 
+ bl[252] br[252] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_255 
+ bl[253] br[253] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_256 
+ bl[254] br[254] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_257 
+ bl[255] br[255] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_258 
+ vdd vdd vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_259 
+ vdd vdd vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_0 
+ vdd vdd vss vdd vpb vnb wl[106] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_108_1 
+ rbl rbr vss vdd vpb vnb wl[106] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_108_2 
+ bl[0] br[0] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_3 
+ bl[1] br[1] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_4 
+ bl[2] br[2] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_5 
+ bl[3] br[3] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_6 
+ bl[4] br[4] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_7 
+ bl[5] br[5] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_8 
+ bl[6] br[6] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_9 
+ bl[7] br[7] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_10 
+ bl[8] br[8] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_11 
+ bl[9] br[9] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_12 
+ bl[10] br[10] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_13 
+ bl[11] br[11] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_14 
+ bl[12] br[12] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_15 
+ bl[13] br[13] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_16 
+ bl[14] br[14] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_17 
+ bl[15] br[15] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_18 
+ bl[16] br[16] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_19 
+ bl[17] br[17] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_20 
+ bl[18] br[18] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_21 
+ bl[19] br[19] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_22 
+ bl[20] br[20] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_23 
+ bl[21] br[21] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_24 
+ bl[22] br[22] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_25 
+ bl[23] br[23] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_26 
+ bl[24] br[24] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_27 
+ bl[25] br[25] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_28 
+ bl[26] br[26] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_29 
+ bl[27] br[27] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_30 
+ bl[28] br[28] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_31 
+ bl[29] br[29] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_32 
+ bl[30] br[30] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_33 
+ bl[31] br[31] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_34 
+ bl[32] br[32] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_35 
+ bl[33] br[33] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_36 
+ bl[34] br[34] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_37 
+ bl[35] br[35] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_38 
+ bl[36] br[36] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_39 
+ bl[37] br[37] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_40 
+ bl[38] br[38] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_41 
+ bl[39] br[39] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_42 
+ bl[40] br[40] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_43 
+ bl[41] br[41] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_44 
+ bl[42] br[42] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_45 
+ bl[43] br[43] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_46 
+ bl[44] br[44] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_47 
+ bl[45] br[45] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_48 
+ bl[46] br[46] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_49 
+ bl[47] br[47] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_50 
+ bl[48] br[48] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_51 
+ bl[49] br[49] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_52 
+ bl[50] br[50] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_53 
+ bl[51] br[51] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_54 
+ bl[52] br[52] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_55 
+ bl[53] br[53] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_56 
+ bl[54] br[54] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_57 
+ bl[55] br[55] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_58 
+ bl[56] br[56] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_59 
+ bl[57] br[57] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_60 
+ bl[58] br[58] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_61 
+ bl[59] br[59] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_62 
+ bl[60] br[60] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_63 
+ bl[61] br[61] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_64 
+ bl[62] br[62] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_65 
+ bl[63] br[63] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_66 
+ bl[64] br[64] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_67 
+ bl[65] br[65] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_68 
+ bl[66] br[66] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_69 
+ bl[67] br[67] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_70 
+ bl[68] br[68] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_71 
+ bl[69] br[69] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_72 
+ bl[70] br[70] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_73 
+ bl[71] br[71] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_74 
+ bl[72] br[72] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_75 
+ bl[73] br[73] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_76 
+ bl[74] br[74] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_77 
+ bl[75] br[75] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_78 
+ bl[76] br[76] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_79 
+ bl[77] br[77] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_80 
+ bl[78] br[78] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_81 
+ bl[79] br[79] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_82 
+ bl[80] br[80] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_83 
+ bl[81] br[81] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_84 
+ bl[82] br[82] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_85 
+ bl[83] br[83] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_86 
+ bl[84] br[84] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_87 
+ bl[85] br[85] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_88 
+ bl[86] br[86] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_89 
+ bl[87] br[87] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_90 
+ bl[88] br[88] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_91 
+ bl[89] br[89] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_92 
+ bl[90] br[90] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_93 
+ bl[91] br[91] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_94 
+ bl[92] br[92] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_95 
+ bl[93] br[93] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_96 
+ bl[94] br[94] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_97 
+ bl[95] br[95] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_98 
+ bl[96] br[96] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_99 
+ bl[97] br[97] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_100 
+ bl[98] br[98] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_101 
+ bl[99] br[99] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_102 
+ bl[100] br[100] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_103 
+ bl[101] br[101] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_104 
+ bl[102] br[102] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_105 
+ bl[103] br[103] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_106 
+ bl[104] br[104] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_107 
+ bl[105] br[105] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_108 
+ bl[106] br[106] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_109 
+ bl[107] br[107] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_110 
+ bl[108] br[108] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_111 
+ bl[109] br[109] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_112 
+ bl[110] br[110] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_113 
+ bl[111] br[111] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_114 
+ bl[112] br[112] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_115 
+ bl[113] br[113] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_116 
+ bl[114] br[114] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_117 
+ bl[115] br[115] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_118 
+ bl[116] br[116] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_119 
+ bl[117] br[117] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_120 
+ bl[118] br[118] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_121 
+ bl[119] br[119] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_122 
+ bl[120] br[120] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_123 
+ bl[121] br[121] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_124 
+ bl[122] br[122] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_125 
+ bl[123] br[123] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_126 
+ bl[124] br[124] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_127 
+ bl[125] br[125] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_128 
+ bl[126] br[126] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_129 
+ bl[127] br[127] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_130 
+ bl[128] br[128] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_131 
+ bl[129] br[129] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_132 
+ bl[130] br[130] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_133 
+ bl[131] br[131] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_134 
+ bl[132] br[132] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_135 
+ bl[133] br[133] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_136 
+ bl[134] br[134] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_137 
+ bl[135] br[135] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_138 
+ bl[136] br[136] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_139 
+ bl[137] br[137] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_140 
+ bl[138] br[138] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_141 
+ bl[139] br[139] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_142 
+ bl[140] br[140] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_143 
+ bl[141] br[141] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_144 
+ bl[142] br[142] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_145 
+ bl[143] br[143] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_146 
+ bl[144] br[144] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_147 
+ bl[145] br[145] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_148 
+ bl[146] br[146] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_149 
+ bl[147] br[147] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_150 
+ bl[148] br[148] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_151 
+ bl[149] br[149] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_152 
+ bl[150] br[150] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_153 
+ bl[151] br[151] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_154 
+ bl[152] br[152] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_155 
+ bl[153] br[153] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_156 
+ bl[154] br[154] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_157 
+ bl[155] br[155] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_158 
+ bl[156] br[156] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_159 
+ bl[157] br[157] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_160 
+ bl[158] br[158] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_161 
+ bl[159] br[159] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_162 
+ bl[160] br[160] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_163 
+ bl[161] br[161] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_164 
+ bl[162] br[162] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_165 
+ bl[163] br[163] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_166 
+ bl[164] br[164] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_167 
+ bl[165] br[165] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_168 
+ bl[166] br[166] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_169 
+ bl[167] br[167] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_170 
+ bl[168] br[168] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_171 
+ bl[169] br[169] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_172 
+ bl[170] br[170] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_173 
+ bl[171] br[171] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_174 
+ bl[172] br[172] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_175 
+ bl[173] br[173] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_176 
+ bl[174] br[174] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_177 
+ bl[175] br[175] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_178 
+ bl[176] br[176] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_179 
+ bl[177] br[177] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_180 
+ bl[178] br[178] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_181 
+ bl[179] br[179] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_182 
+ bl[180] br[180] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_183 
+ bl[181] br[181] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_184 
+ bl[182] br[182] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_185 
+ bl[183] br[183] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_186 
+ bl[184] br[184] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_187 
+ bl[185] br[185] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_188 
+ bl[186] br[186] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_189 
+ bl[187] br[187] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_190 
+ bl[188] br[188] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_191 
+ bl[189] br[189] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_192 
+ bl[190] br[190] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_193 
+ bl[191] br[191] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_194 
+ bl[192] br[192] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_195 
+ bl[193] br[193] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_196 
+ bl[194] br[194] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_197 
+ bl[195] br[195] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_198 
+ bl[196] br[196] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_199 
+ bl[197] br[197] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_200 
+ bl[198] br[198] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_201 
+ bl[199] br[199] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_202 
+ bl[200] br[200] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_203 
+ bl[201] br[201] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_204 
+ bl[202] br[202] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_205 
+ bl[203] br[203] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_206 
+ bl[204] br[204] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_207 
+ bl[205] br[205] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_208 
+ bl[206] br[206] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_209 
+ bl[207] br[207] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_210 
+ bl[208] br[208] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_211 
+ bl[209] br[209] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_212 
+ bl[210] br[210] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_213 
+ bl[211] br[211] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_214 
+ bl[212] br[212] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_215 
+ bl[213] br[213] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_216 
+ bl[214] br[214] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_217 
+ bl[215] br[215] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_218 
+ bl[216] br[216] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_219 
+ bl[217] br[217] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_220 
+ bl[218] br[218] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_221 
+ bl[219] br[219] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_222 
+ bl[220] br[220] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_223 
+ bl[221] br[221] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_224 
+ bl[222] br[222] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_225 
+ bl[223] br[223] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_226 
+ bl[224] br[224] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_227 
+ bl[225] br[225] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_228 
+ bl[226] br[226] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_229 
+ bl[227] br[227] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_230 
+ bl[228] br[228] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_231 
+ bl[229] br[229] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_232 
+ bl[230] br[230] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_233 
+ bl[231] br[231] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_234 
+ bl[232] br[232] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_235 
+ bl[233] br[233] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_236 
+ bl[234] br[234] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_237 
+ bl[235] br[235] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_238 
+ bl[236] br[236] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_239 
+ bl[237] br[237] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_240 
+ bl[238] br[238] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_241 
+ bl[239] br[239] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_242 
+ bl[240] br[240] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_243 
+ bl[241] br[241] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_244 
+ bl[242] br[242] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_245 
+ bl[243] br[243] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_246 
+ bl[244] br[244] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_247 
+ bl[245] br[245] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_248 
+ bl[246] br[246] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_249 
+ bl[247] br[247] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_250 
+ bl[248] br[248] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_251 
+ bl[249] br[249] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_252 
+ bl[250] br[250] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_253 
+ bl[251] br[251] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_254 
+ bl[252] br[252] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_255 
+ bl[253] br[253] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_256 
+ bl[254] br[254] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_257 
+ bl[255] br[255] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_258 
+ vdd vdd vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_259 
+ vdd vdd vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_0 
+ vdd vdd vss vdd vpb vnb wl[107] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_109_1 
+ rbl rbr vss vdd vpb vnb wl[107] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_109_2 
+ bl[0] br[0] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_3 
+ bl[1] br[1] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_4 
+ bl[2] br[2] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_5 
+ bl[3] br[3] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_6 
+ bl[4] br[4] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_7 
+ bl[5] br[5] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_8 
+ bl[6] br[6] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_9 
+ bl[7] br[7] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_10 
+ bl[8] br[8] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_11 
+ bl[9] br[9] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_12 
+ bl[10] br[10] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_13 
+ bl[11] br[11] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_14 
+ bl[12] br[12] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_15 
+ bl[13] br[13] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_16 
+ bl[14] br[14] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_17 
+ bl[15] br[15] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_18 
+ bl[16] br[16] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_19 
+ bl[17] br[17] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_20 
+ bl[18] br[18] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_21 
+ bl[19] br[19] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_22 
+ bl[20] br[20] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_23 
+ bl[21] br[21] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_24 
+ bl[22] br[22] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_25 
+ bl[23] br[23] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_26 
+ bl[24] br[24] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_27 
+ bl[25] br[25] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_28 
+ bl[26] br[26] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_29 
+ bl[27] br[27] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_30 
+ bl[28] br[28] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_31 
+ bl[29] br[29] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_32 
+ bl[30] br[30] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_33 
+ bl[31] br[31] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_34 
+ bl[32] br[32] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_35 
+ bl[33] br[33] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_36 
+ bl[34] br[34] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_37 
+ bl[35] br[35] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_38 
+ bl[36] br[36] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_39 
+ bl[37] br[37] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_40 
+ bl[38] br[38] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_41 
+ bl[39] br[39] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_42 
+ bl[40] br[40] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_43 
+ bl[41] br[41] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_44 
+ bl[42] br[42] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_45 
+ bl[43] br[43] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_46 
+ bl[44] br[44] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_47 
+ bl[45] br[45] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_48 
+ bl[46] br[46] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_49 
+ bl[47] br[47] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_50 
+ bl[48] br[48] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_51 
+ bl[49] br[49] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_52 
+ bl[50] br[50] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_53 
+ bl[51] br[51] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_54 
+ bl[52] br[52] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_55 
+ bl[53] br[53] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_56 
+ bl[54] br[54] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_57 
+ bl[55] br[55] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_58 
+ bl[56] br[56] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_59 
+ bl[57] br[57] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_60 
+ bl[58] br[58] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_61 
+ bl[59] br[59] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_62 
+ bl[60] br[60] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_63 
+ bl[61] br[61] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_64 
+ bl[62] br[62] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_65 
+ bl[63] br[63] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_66 
+ bl[64] br[64] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_67 
+ bl[65] br[65] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_68 
+ bl[66] br[66] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_69 
+ bl[67] br[67] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_70 
+ bl[68] br[68] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_71 
+ bl[69] br[69] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_72 
+ bl[70] br[70] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_73 
+ bl[71] br[71] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_74 
+ bl[72] br[72] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_75 
+ bl[73] br[73] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_76 
+ bl[74] br[74] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_77 
+ bl[75] br[75] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_78 
+ bl[76] br[76] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_79 
+ bl[77] br[77] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_80 
+ bl[78] br[78] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_81 
+ bl[79] br[79] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_82 
+ bl[80] br[80] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_83 
+ bl[81] br[81] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_84 
+ bl[82] br[82] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_85 
+ bl[83] br[83] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_86 
+ bl[84] br[84] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_87 
+ bl[85] br[85] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_88 
+ bl[86] br[86] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_89 
+ bl[87] br[87] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_90 
+ bl[88] br[88] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_91 
+ bl[89] br[89] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_92 
+ bl[90] br[90] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_93 
+ bl[91] br[91] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_94 
+ bl[92] br[92] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_95 
+ bl[93] br[93] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_96 
+ bl[94] br[94] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_97 
+ bl[95] br[95] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_98 
+ bl[96] br[96] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_99 
+ bl[97] br[97] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_100 
+ bl[98] br[98] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_101 
+ bl[99] br[99] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_102 
+ bl[100] br[100] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_103 
+ bl[101] br[101] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_104 
+ bl[102] br[102] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_105 
+ bl[103] br[103] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_106 
+ bl[104] br[104] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_107 
+ bl[105] br[105] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_108 
+ bl[106] br[106] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_109 
+ bl[107] br[107] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_110 
+ bl[108] br[108] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_111 
+ bl[109] br[109] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_112 
+ bl[110] br[110] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_113 
+ bl[111] br[111] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_114 
+ bl[112] br[112] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_115 
+ bl[113] br[113] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_116 
+ bl[114] br[114] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_117 
+ bl[115] br[115] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_118 
+ bl[116] br[116] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_119 
+ bl[117] br[117] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_120 
+ bl[118] br[118] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_121 
+ bl[119] br[119] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_122 
+ bl[120] br[120] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_123 
+ bl[121] br[121] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_124 
+ bl[122] br[122] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_125 
+ bl[123] br[123] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_126 
+ bl[124] br[124] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_127 
+ bl[125] br[125] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_128 
+ bl[126] br[126] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_129 
+ bl[127] br[127] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_130 
+ bl[128] br[128] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_131 
+ bl[129] br[129] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_132 
+ bl[130] br[130] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_133 
+ bl[131] br[131] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_134 
+ bl[132] br[132] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_135 
+ bl[133] br[133] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_136 
+ bl[134] br[134] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_137 
+ bl[135] br[135] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_138 
+ bl[136] br[136] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_139 
+ bl[137] br[137] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_140 
+ bl[138] br[138] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_141 
+ bl[139] br[139] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_142 
+ bl[140] br[140] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_143 
+ bl[141] br[141] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_144 
+ bl[142] br[142] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_145 
+ bl[143] br[143] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_146 
+ bl[144] br[144] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_147 
+ bl[145] br[145] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_148 
+ bl[146] br[146] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_149 
+ bl[147] br[147] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_150 
+ bl[148] br[148] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_151 
+ bl[149] br[149] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_152 
+ bl[150] br[150] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_153 
+ bl[151] br[151] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_154 
+ bl[152] br[152] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_155 
+ bl[153] br[153] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_156 
+ bl[154] br[154] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_157 
+ bl[155] br[155] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_158 
+ bl[156] br[156] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_159 
+ bl[157] br[157] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_160 
+ bl[158] br[158] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_161 
+ bl[159] br[159] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_162 
+ bl[160] br[160] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_163 
+ bl[161] br[161] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_164 
+ bl[162] br[162] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_165 
+ bl[163] br[163] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_166 
+ bl[164] br[164] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_167 
+ bl[165] br[165] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_168 
+ bl[166] br[166] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_169 
+ bl[167] br[167] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_170 
+ bl[168] br[168] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_171 
+ bl[169] br[169] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_172 
+ bl[170] br[170] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_173 
+ bl[171] br[171] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_174 
+ bl[172] br[172] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_175 
+ bl[173] br[173] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_176 
+ bl[174] br[174] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_177 
+ bl[175] br[175] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_178 
+ bl[176] br[176] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_179 
+ bl[177] br[177] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_180 
+ bl[178] br[178] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_181 
+ bl[179] br[179] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_182 
+ bl[180] br[180] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_183 
+ bl[181] br[181] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_184 
+ bl[182] br[182] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_185 
+ bl[183] br[183] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_186 
+ bl[184] br[184] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_187 
+ bl[185] br[185] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_188 
+ bl[186] br[186] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_189 
+ bl[187] br[187] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_190 
+ bl[188] br[188] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_191 
+ bl[189] br[189] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_192 
+ bl[190] br[190] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_193 
+ bl[191] br[191] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_194 
+ bl[192] br[192] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_195 
+ bl[193] br[193] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_196 
+ bl[194] br[194] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_197 
+ bl[195] br[195] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_198 
+ bl[196] br[196] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_199 
+ bl[197] br[197] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_200 
+ bl[198] br[198] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_201 
+ bl[199] br[199] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_202 
+ bl[200] br[200] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_203 
+ bl[201] br[201] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_204 
+ bl[202] br[202] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_205 
+ bl[203] br[203] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_206 
+ bl[204] br[204] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_207 
+ bl[205] br[205] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_208 
+ bl[206] br[206] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_209 
+ bl[207] br[207] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_210 
+ bl[208] br[208] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_211 
+ bl[209] br[209] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_212 
+ bl[210] br[210] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_213 
+ bl[211] br[211] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_214 
+ bl[212] br[212] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_215 
+ bl[213] br[213] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_216 
+ bl[214] br[214] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_217 
+ bl[215] br[215] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_218 
+ bl[216] br[216] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_219 
+ bl[217] br[217] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_220 
+ bl[218] br[218] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_221 
+ bl[219] br[219] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_222 
+ bl[220] br[220] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_223 
+ bl[221] br[221] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_224 
+ bl[222] br[222] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_225 
+ bl[223] br[223] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_226 
+ bl[224] br[224] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_227 
+ bl[225] br[225] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_228 
+ bl[226] br[226] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_229 
+ bl[227] br[227] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_230 
+ bl[228] br[228] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_231 
+ bl[229] br[229] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_232 
+ bl[230] br[230] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_233 
+ bl[231] br[231] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_234 
+ bl[232] br[232] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_235 
+ bl[233] br[233] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_236 
+ bl[234] br[234] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_237 
+ bl[235] br[235] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_238 
+ bl[236] br[236] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_239 
+ bl[237] br[237] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_240 
+ bl[238] br[238] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_241 
+ bl[239] br[239] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_242 
+ bl[240] br[240] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_243 
+ bl[241] br[241] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_244 
+ bl[242] br[242] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_245 
+ bl[243] br[243] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_246 
+ bl[244] br[244] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_247 
+ bl[245] br[245] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_248 
+ bl[246] br[246] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_249 
+ bl[247] br[247] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_250 
+ bl[248] br[248] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_251 
+ bl[249] br[249] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_252 
+ bl[250] br[250] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_253 
+ bl[251] br[251] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_254 
+ bl[252] br[252] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_255 
+ bl[253] br[253] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_256 
+ bl[254] br[254] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_257 
+ bl[255] br[255] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_258 
+ vdd vdd vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_259 
+ vdd vdd vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_0 
+ vdd vdd vss vdd vpb vnb wl[108] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_110_1 
+ rbl rbr vss vdd vpb vnb wl[108] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_110_2 
+ bl[0] br[0] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_3 
+ bl[1] br[1] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_4 
+ bl[2] br[2] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_5 
+ bl[3] br[3] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_6 
+ bl[4] br[4] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_7 
+ bl[5] br[5] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_8 
+ bl[6] br[6] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_9 
+ bl[7] br[7] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_10 
+ bl[8] br[8] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_11 
+ bl[9] br[9] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_12 
+ bl[10] br[10] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_13 
+ bl[11] br[11] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_14 
+ bl[12] br[12] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_15 
+ bl[13] br[13] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_16 
+ bl[14] br[14] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_17 
+ bl[15] br[15] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_18 
+ bl[16] br[16] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_19 
+ bl[17] br[17] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_20 
+ bl[18] br[18] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_21 
+ bl[19] br[19] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_22 
+ bl[20] br[20] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_23 
+ bl[21] br[21] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_24 
+ bl[22] br[22] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_25 
+ bl[23] br[23] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_26 
+ bl[24] br[24] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_27 
+ bl[25] br[25] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_28 
+ bl[26] br[26] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_29 
+ bl[27] br[27] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_30 
+ bl[28] br[28] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_31 
+ bl[29] br[29] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_32 
+ bl[30] br[30] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_33 
+ bl[31] br[31] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_34 
+ bl[32] br[32] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_35 
+ bl[33] br[33] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_36 
+ bl[34] br[34] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_37 
+ bl[35] br[35] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_38 
+ bl[36] br[36] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_39 
+ bl[37] br[37] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_40 
+ bl[38] br[38] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_41 
+ bl[39] br[39] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_42 
+ bl[40] br[40] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_43 
+ bl[41] br[41] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_44 
+ bl[42] br[42] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_45 
+ bl[43] br[43] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_46 
+ bl[44] br[44] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_47 
+ bl[45] br[45] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_48 
+ bl[46] br[46] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_49 
+ bl[47] br[47] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_50 
+ bl[48] br[48] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_51 
+ bl[49] br[49] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_52 
+ bl[50] br[50] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_53 
+ bl[51] br[51] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_54 
+ bl[52] br[52] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_55 
+ bl[53] br[53] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_56 
+ bl[54] br[54] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_57 
+ bl[55] br[55] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_58 
+ bl[56] br[56] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_59 
+ bl[57] br[57] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_60 
+ bl[58] br[58] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_61 
+ bl[59] br[59] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_62 
+ bl[60] br[60] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_63 
+ bl[61] br[61] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_64 
+ bl[62] br[62] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_65 
+ bl[63] br[63] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_66 
+ bl[64] br[64] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_67 
+ bl[65] br[65] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_68 
+ bl[66] br[66] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_69 
+ bl[67] br[67] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_70 
+ bl[68] br[68] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_71 
+ bl[69] br[69] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_72 
+ bl[70] br[70] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_73 
+ bl[71] br[71] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_74 
+ bl[72] br[72] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_75 
+ bl[73] br[73] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_76 
+ bl[74] br[74] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_77 
+ bl[75] br[75] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_78 
+ bl[76] br[76] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_79 
+ bl[77] br[77] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_80 
+ bl[78] br[78] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_81 
+ bl[79] br[79] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_82 
+ bl[80] br[80] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_83 
+ bl[81] br[81] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_84 
+ bl[82] br[82] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_85 
+ bl[83] br[83] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_86 
+ bl[84] br[84] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_87 
+ bl[85] br[85] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_88 
+ bl[86] br[86] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_89 
+ bl[87] br[87] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_90 
+ bl[88] br[88] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_91 
+ bl[89] br[89] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_92 
+ bl[90] br[90] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_93 
+ bl[91] br[91] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_94 
+ bl[92] br[92] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_95 
+ bl[93] br[93] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_96 
+ bl[94] br[94] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_97 
+ bl[95] br[95] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_98 
+ bl[96] br[96] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_99 
+ bl[97] br[97] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_100 
+ bl[98] br[98] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_101 
+ bl[99] br[99] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_102 
+ bl[100] br[100] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_103 
+ bl[101] br[101] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_104 
+ bl[102] br[102] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_105 
+ bl[103] br[103] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_106 
+ bl[104] br[104] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_107 
+ bl[105] br[105] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_108 
+ bl[106] br[106] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_109 
+ bl[107] br[107] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_110 
+ bl[108] br[108] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_111 
+ bl[109] br[109] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_112 
+ bl[110] br[110] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_113 
+ bl[111] br[111] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_114 
+ bl[112] br[112] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_115 
+ bl[113] br[113] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_116 
+ bl[114] br[114] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_117 
+ bl[115] br[115] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_118 
+ bl[116] br[116] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_119 
+ bl[117] br[117] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_120 
+ bl[118] br[118] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_121 
+ bl[119] br[119] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_122 
+ bl[120] br[120] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_123 
+ bl[121] br[121] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_124 
+ bl[122] br[122] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_125 
+ bl[123] br[123] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_126 
+ bl[124] br[124] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_127 
+ bl[125] br[125] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_128 
+ bl[126] br[126] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_129 
+ bl[127] br[127] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_130 
+ bl[128] br[128] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_131 
+ bl[129] br[129] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_132 
+ bl[130] br[130] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_133 
+ bl[131] br[131] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_134 
+ bl[132] br[132] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_135 
+ bl[133] br[133] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_136 
+ bl[134] br[134] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_137 
+ bl[135] br[135] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_138 
+ bl[136] br[136] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_139 
+ bl[137] br[137] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_140 
+ bl[138] br[138] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_141 
+ bl[139] br[139] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_142 
+ bl[140] br[140] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_143 
+ bl[141] br[141] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_144 
+ bl[142] br[142] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_145 
+ bl[143] br[143] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_146 
+ bl[144] br[144] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_147 
+ bl[145] br[145] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_148 
+ bl[146] br[146] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_149 
+ bl[147] br[147] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_150 
+ bl[148] br[148] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_151 
+ bl[149] br[149] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_152 
+ bl[150] br[150] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_153 
+ bl[151] br[151] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_154 
+ bl[152] br[152] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_155 
+ bl[153] br[153] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_156 
+ bl[154] br[154] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_157 
+ bl[155] br[155] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_158 
+ bl[156] br[156] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_159 
+ bl[157] br[157] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_160 
+ bl[158] br[158] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_161 
+ bl[159] br[159] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_162 
+ bl[160] br[160] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_163 
+ bl[161] br[161] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_164 
+ bl[162] br[162] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_165 
+ bl[163] br[163] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_166 
+ bl[164] br[164] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_167 
+ bl[165] br[165] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_168 
+ bl[166] br[166] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_169 
+ bl[167] br[167] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_170 
+ bl[168] br[168] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_171 
+ bl[169] br[169] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_172 
+ bl[170] br[170] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_173 
+ bl[171] br[171] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_174 
+ bl[172] br[172] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_175 
+ bl[173] br[173] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_176 
+ bl[174] br[174] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_177 
+ bl[175] br[175] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_178 
+ bl[176] br[176] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_179 
+ bl[177] br[177] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_180 
+ bl[178] br[178] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_181 
+ bl[179] br[179] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_182 
+ bl[180] br[180] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_183 
+ bl[181] br[181] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_184 
+ bl[182] br[182] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_185 
+ bl[183] br[183] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_186 
+ bl[184] br[184] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_187 
+ bl[185] br[185] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_188 
+ bl[186] br[186] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_189 
+ bl[187] br[187] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_190 
+ bl[188] br[188] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_191 
+ bl[189] br[189] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_192 
+ bl[190] br[190] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_193 
+ bl[191] br[191] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_194 
+ bl[192] br[192] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_195 
+ bl[193] br[193] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_196 
+ bl[194] br[194] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_197 
+ bl[195] br[195] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_198 
+ bl[196] br[196] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_199 
+ bl[197] br[197] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_200 
+ bl[198] br[198] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_201 
+ bl[199] br[199] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_202 
+ bl[200] br[200] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_203 
+ bl[201] br[201] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_204 
+ bl[202] br[202] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_205 
+ bl[203] br[203] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_206 
+ bl[204] br[204] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_207 
+ bl[205] br[205] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_208 
+ bl[206] br[206] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_209 
+ bl[207] br[207] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_210 
+ bl[208] br[208] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_211 
+ bl[209] br[209] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_212 
+ bl[210] br[210] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_213 
+ bl[211] br[211] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_214 
+ bl[212] br[212] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_215 
+ bl[213] br[213] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_216 
+ bl[214] br[214] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_217 
+ bl[215] br[215] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_218 
+ bl[216] br[216] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_219 
+ bl[217] br[217] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_220 
+ bl[218] br[218] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_221 
+ bl[219] br[219] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_222 
+ bl[220] br[220] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_223 
+ bl[221] br[221] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_224 
+ bl[222] br[222] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_225 
+ bl[223] br[223] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_226 
+ bl[224] br[224] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_227 
+ bl[225] br[225] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_228 
+ bl[226] br[226] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_229 
+ bl[227] br[227] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_230 
+ bl[228] br[228] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_231 
+ bl[229] br[229] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_232 
+ bl[230] br[230] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_233 
+ bl[231] br[231] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_234 
+ bl[232] br[232] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_235 
+ bl[233] br[233] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_236 
+ bl[234] br[234] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_237 
+ bl[235] br[235] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_238 
+ bl[236] br[236] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_239 
+ bl[237] br[237] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_240 
+ bl[238] br[238] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_241 
+ bl[239] br[239] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_242 
+ bl[240] br[240] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_243 
+ bl[241] br[241] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_244 
+ bl[242] br[242] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_245 
+ bl[243] br[243] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_246 
+ bl[244] br[244] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_247 
+ bl[245] br[245] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_248 
+ bl[246] br[246] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_249 
+ bl[247] br[247] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_250 
+ bl[248] br[248] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_251 
+ bl[249] br[249] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_252 
+ bl[250] br[250] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_253 
+ bl[251] br[251] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_254 
+ bl[252] br[252] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_255 
+ bl[253] br[253] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_256 
+ bl[254] br[254] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_257 
+ bl[255] br[255] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_258 
+ vdd vdd vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_259 
+ vdd vdd vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_0 
+ vdd vdd vss vdd vpb vnb wl[109] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_111_1 
+ rbl rbr vss vdd vpb vnb wl[109] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_111_2 
+ bl[0] br[0] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_3 
+ bl[1] br[1] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_4 
+ bl[2] br[2] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_5 
+ bl[3] br[3] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_6 
+ bl[4] br[4] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_7 
+ bl[5] br[5] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_8 
+ bl[6] br[6] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_9 
+ bl[7] br[7] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_10 
+ bl[8] br[8] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_11 
+ bl[9] br[9] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_12 
+ bl[10] br[10] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_13 
+ bl[11] br[11] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_14 
+ bl[12] br[12] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_15 
+ bl[13] br[13] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_16 
+ bl[14] br[14] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_17 
+ bl[15] br[15] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_18 
+ bl[16] br[16] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_19 
+ bl[17] br[17] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_20 
+ bl[18] br[18] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_21 
+ bl[19] br[19] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_22 
+ bl[20] br[20] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_23 
+ bl[21] br[21] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_24 
+ bl[22] br[22] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_25 
+ bl[23] br[23] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_26 
+ bl[24] br[24] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_27 
+ bl[25] br[25] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_28 
+ bl[26] br[26] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_29 
+ bl[27] br[27] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_30 
+ bl[28] br[28] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_31 
+ bl[29] br[29] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_32 
+ bl[30] br[30] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_33 
+ bl[31] br[31] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_34 
+ bl[32] br[32] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_35 
+ bl[33] br[33] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_36 
+ bl[34] br[34] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_37 
+ bl[35] br[35] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_38 
+ bl[36] br[36] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_39 
+ bl[37] br[37] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_40 
+ bl[38] br[38] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_41 
+ bl[39] br[39] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_42 
+ bl[40] br[40] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_43 
+ bl[41] br[41] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_44 
+ bl[42] br[42] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_45 
+ bl[43] br[43] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_46 
+ bl[44] br[44] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_47 
+ bl[45] br[45] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_48 
+ bl[46] br[46] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_49 
+ bl[47] br[47] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_50 
+ bl[48] br[48] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_51 
+ bl[49] br[49] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_52 
+ bl[50] br[50] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_53 
+ bl[51] br[51] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_54 
+ bl[52] br[52] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_55 
+ bl[53] br[53] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_56 
+ bl[54] br[54] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_57 
+ bl[55] br[55] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_58 
+ bl[56] br[56] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_59 
+ bl[57] br[57] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_60 
+ bl[58] br[58] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_61 
+ bl[59] br[59] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_62 
+ bl[60] br[60] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_63 
+ bl[61] br[61] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_64 
+ bl[62] br[62] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_65 
+ bl[63] br[63] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_66 
+ bl[64] br[64] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_67 
+ bl[65] br[65] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_68 
+ bl[66] br[66] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_69 
+ bl[67] br[67] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_70 
+ bl[68] br[68] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_71 
+ bl[69] br[69] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_72 
+ bl[70] br[70] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_73 
+ bl[71] br[71] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_74 
+ bl[72] br[72] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_75 
+ bl[73] br[73] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_76 
+ bl[74] br[74] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_77 
+ bl[75] br[75] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_78 
+ bl[76] br[76] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_79 
+ bl[77] br[77] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_80 
+ bl[78] br[78] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_81 
+ bl[79] br[79] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_82 
+ bl[80] br[80] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_83 
+ bl[81] br[81] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_84 
+ bl[82] br[82] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_85 
+ bl[83] br[83] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_86 
+ bl[84] br[84] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_87 
+ bl[85] br[85] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_88 
+ bl[86] br[86] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_89 
+ bl[87] br[87] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_90 
+ bl[88] br[88] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_91 
+ bl[89] br[89] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_92 
+ bl[90] br[90] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_93 
+ bl[91] br[91] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_94 
+ bl[92] br[92] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_95 
+ bl[93] br[93] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_96 
+ bl[94] br[94] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_97 
+ bl[95] br[95] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_98 
+ bl[96] br[96] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_99 
+ bl[97] br[97] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_100 
+ bl[98] br[98] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_101 
+ bl[99] br[99] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_102 
+ bl[100] br[100] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_103 
+ bl[101] br[101] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_104 
+ bl[102] br[102] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_105 
+ bl[103] br[103] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_106 
+ bl[104] br[104] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_107 
+ bl[105] br[105] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_108 
+ bl[106] br[106] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_109 
+ bl[107] br[107] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_110 
+ bl[108] br[108] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_111 
+ bl[109] br[109] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_112 
+ bl[110] br[110] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_113 
+ bl[111] br[111] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_114 
+ bl[112] br[112] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_115 
+ bl[113] br[113] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_116 
+ bl[114] br[114] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_117 
+ bl[115] br[115] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_118 
+ bl[116] br[116] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_119 
+ bl[117] br[117] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_120 
+ bl[118] br[118] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_121 
+ bl[119] br[119] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_122 
+ bl[120] br[120] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_123 
+ bl[121] br[121] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_124 
+ bl[122] br[122] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_125 
+ bl[123] br[123] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_126 
+ bl[124] br[124] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_127 
+ bl[125] br[125] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_128 
+ bl[126] br[126] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_129 
+ bl[127] br[127] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_130 
+ bl[128] br[128] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_131 
+ bl[129] br[129] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_132 
+ bl[130] br[130] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_133 
+ bl[131] br[131] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_134 
+ bl[132] br[132] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_135 
+ bl[133] br[133] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_136 
+ bl[134] br[134] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_137 
+ bl[135] br[135] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_138 
+ bl[136] br[136] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_139 
+ bl[137] br[137] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_140 
+ bl[138] br[138] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_141 
+ bl[139] br[139] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_142 
+ bl[140] br[140] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_143 
+ bl[141] br[141] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_144 
+ bl[142] br[142] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_145 
+ bl[143] br[143] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_146 
+ bl[144] br[144] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_147 
+ bl[145] br[145] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_148 
+ bl[146] br[146] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_149 
+ bl[147] br[147] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_150 
+ bl[148] br[148] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_151 
+ bl[149] br[149] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_152 
+ bl[150] br[150] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_153 
+ bl[151] br[151] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_154 
+ bl[152] br[152] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_155 
+ bl[153] br[153] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_156 
+ bl[154] br[154] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_157 
+ bl[155] br[155] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_158 
+ bl[156] br[156] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_159 
+ bl[157] br[157] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_160 
+ bl[158] br[158] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_161 
+ bl[159] br[159] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_162 
+ bl[160] br[160] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_163 
+ bl[161] br[161] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_164 
+ bl[162] br[162] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_165 
+ bl[163] br[163] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_166 
+ bl[164] br[164] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_167 
+ bl[165] br[165] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_168 
+ bl[166] br[166] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_169 
+ bl[167] br[167] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_170 
+ bl[168] br[168] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_171 
+ bl[169] br[169] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_172 
+ bl[170] br[170] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_173 
+ bl[171] br[171] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_174 
+ bl[172] br[172] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_175 
+ bl[173] br[173] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_176 
+ bl[174] br[174] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_177 
+ bl[175] br[175] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_178 
+ bl[176] br[176] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_179 
+ bl[177] br[177] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_180 
+ bl[178] br[178] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_181 
+ bl[179] br[179] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_182 
+ bl[180] br[180] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_183 
+ bl[181] br[181] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_184 
+ bl[182] br[182] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_185 
+ bl[183] br[183] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_186 
+ bl[184] br[184] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_187 
+ bl[185] br[185] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_188 
+ bl[186] br[186] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_189 
+ bl[187] br[187] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_190 
+ bl[188] br[188] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_191 
+ bl[189] br[189] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_192 
+ bl[190] br[190] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_193 
+ bl[191] br[191] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_194 
+ bl[192] br[192] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_195 
+ bl[193] br[193] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_196 
+ bl[194] br[194] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_197 
+ bl[195] br[195] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_198 
+ bl[196] br[196] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_199 
+ bl[197] br[197] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_200 
+ bl[198] br[198] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_201 
+ bl[199] br[199] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_202 
+ bl[200] br[200] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_203 
+ bl[201] br[201] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_204 
+ bl[202] br[202] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_205 
+ bl[203] br[203] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_206 
+ bl[204] br[204] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_207 
+ bl[205] br[205] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_208 
+ bl[206] br[206] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_209 
+ bl[207] br[207] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_210 
+ bl[208] br[208] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_211 
+ bl[209] br[209] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_212 
+ bl[210] br[210] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_213 
+ bl[211] br[211] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_214 
+ bl[212] br[212] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_215 
+ bl[213] br[213] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_216 
+ bl[214] br[214] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_217 
+ bl[215] br[215] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_218 
+ bl[216] br[216] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_219 
+ bl[217] br[217] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_220 
+ bl[218] br[218] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_221 
+ bl[219] br[219] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_222 
+ bl[220] br[220] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_223 
+ bl[221] br[221] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_224 
+ bl[222] br[222] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_225 
+ bl[223] br[223] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_226 
+ bl[224] br[224] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_227 
+ bl[225] br[225] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_228 
+ bl[226] br[226] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_229 
+ bl[227] br[227] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_230 
+ bl[228] br[228] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_231 
+ bl[229] br[229] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_232 
+ bl[230] br[230] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_233 
+ bl[231] br[231] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_234 
+ bl[232] br[232] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_235 
+ bl[233] br[233] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_236 
+ bl[234] br[234] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_237 
+ bl[235] br[235] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_238 
+ bl[236] br[236] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_239 
+ bl[237] br[237] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_240 
+ bl[238] br[238] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_241 
+ bl[239] br[239] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_242 
+ bl[240] br[240] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_243 
+ bl[241] br[241] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_244 
+ bl[242] br[242] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_245 
+ bl[243] br[243] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_246 
+ bl[244] br[244] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_247 
+ bl[245] br[245] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_248 
+ bl[246] br[246] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_249 
+ bl[247] br[247] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_250 
+ bl[248] br[248] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_251 
+ bl[249] br[249] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_252 
+ bl[250] br[250] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_253 
+ bl[251] br[251] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_254 
+ bl[252] br[252] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_255 
+ bl[253] br[253] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_256 
+ bl[254] br[254] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_257 
+ bl[255] br[255] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_258 
+ vdd vdd vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_259 
+ vdd vdd vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_0 
+ vdd vdd vss vdd vpb vnb wl[110] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_112_1 
+ rbl rbr vss vdd vpb vnb wl[110] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_112_2 
+ bl[0] br[0] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_3 
+ bl[1] br[1] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_4 
+ bl[2] br[2] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_5 
+ bl[3] br[3] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_6 
+ bl[4] br[4] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_7 
+ bl[5] br[5] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_8 
+ bl[6] br[6] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_9 
+ bl[7] br[7] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_10 
+ bl[8] br[8] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_11 
+ bl[9] br[9] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_12 
+ bl[10] br[10] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_13 
+ bl[11] br[11] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_14 
+ bl[12] br[12] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_15 
+ bl[13] br[13] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_16 
+ bl[14] br[14] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_17 
+ bl[15] br[15] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_18 
+ bl[16] br[16] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_19 
+ bl[17] br[17] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_20 
+ bl[18] br[18] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_21 
+ bl[19] br[19] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_22 
+ bl[20] br[20] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_23 
+ bl[21] br[21] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_24 
+ bl[22] br[22] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_25 
+ bl[23] br[23] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_26 
+ bl[24] br[24] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_27 
+ bl[25] br[25] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_28 
+ bl[26] br[26] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_29 
+ bl[27] br[27] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_30 
+ bl[28] br[28] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_31 
+ bl[29] br[29] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_32 
+ bl[30] br[30] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_33 
+ bl[31] br[31] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_34 
+ bl[32] br[32] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_35 
+ bl[33] br[33] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_36 
+ bl[34] br[34] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_37 
+ bl[35] br[35] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_38 
+ bl[36] br[36] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_39 
+ bl[37] br[37] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_40 
+ bl[38] br[38] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_41 
+ bl[39] br[39] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_42 
+ bl[40] br[40] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_43 
+ bl[41] br[41] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_44 
+ bl[42] br[42] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_45 
+ bl[43] br[43] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_46 
+ bl[44] br[44] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_47 
+ bl[45] br[45] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_48 
+ bl[46] br[46] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_49 
+ bl[47] br[47] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_50 
+ bl[48] br[48] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_51 
+ bl[49] br[49] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_52 
+ bl[50] br[50] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_53 
+ bl[51] br[51] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_54 
+ bl[52] br[52] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_55 
+ bl[53] br[53] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_56 
+ bl[54] br[54] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_57 
+ bl[55] br[55] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_58 
+ bl[56] br[56] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_59 
+ bl[57] br[57] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_60 
+ bl[58] br[58] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_61 
+ bl[59] br[59] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_62 
+ bl[60] br[60] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_63 
+ bl[61] br[61] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_64 
+ bl[62] br[62] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_65 
+ bl[63] br[63] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_66 
+ bl[64] br[64] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_67 
+ bl[65] br[65] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_68 
+ bl[66] br[66] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_69 
+ bl[67] br[67] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_70 
+ bl[68] br[68] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_71 
+ bl[69] br[69] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_72 
+ bl[70] br[70] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_73 
+ bl[71] br[71] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_74 
+ bl[72] br[72] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_75 
+ bl[73] br[73] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_76 
+ bl[74] br[74] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_77 
+ bl[75] br[75] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_78 
+ bl[76] br[76] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_79 
+ bl[77] br[77] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_80 
+ bl[78] br[78] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_81 
+ bl[79] br[79] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_82 
+ bl[80] br[80] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_83 
+ bl[81] br[81] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_84 
+ bl[82] br[82] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_85 
+ bl[83] br[83] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_86 
+ bl[84] br[84] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_87 
+ bl[85] br[85] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_88 
+ bl[86] br[86] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_89 
+ bl[87] br[87] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_90 
+ bl[88] br[88] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_91 
+ bl[89] br[89] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_92 
+ bl[90] br[90] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_93 
+ bl[91] br[91] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_94 
+ bl[92] br[92] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_95 
+ bl[93] br[93] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_96 
+ bl[94] br[94] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_97 
+ bl[95] br[95] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_98 
+ bl[96] br[96] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_99 
+ bl[97] br[97] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_100 
+ bl[98] br[98] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_101 
+ bl[99] br[99] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_102 
+ bl[100] br[100] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_103 
+ bl[101] br[101] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_104 
+ bl[102] br[102] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_105 
+ bl[103] br[103] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_106 
+ bl[104] br[104] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_107 
+ bl[105] br[105] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_108 
+ bl[106] br[106] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_109 
+ bl[107] br[107] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_110 
+ bl[108] br[108] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_111 
+ bl[109] br[109] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_112 
+ bl[110] br[110] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_113 
+ bl[111] br[111] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_114 
+ bl[112] br[112] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_115 
+ bl[113] br[113] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_116 
+ bl[114] br[114] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_117 
+ bl[115] br[115] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_118 
+ bl[116] br[116] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_119 
+ bl[117] br[117] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_120 
+ bl[118] br[118] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_121 
+ bl[119] br[119] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_122 
+ bl[120] br[120] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_123 
+ bl[121] br[121] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_124 
+ bl[122] br[122] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_125 
+ bl[123] br[123] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_126 
+ bl[124] br[124] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_127 
+ bl[125] br[125] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_128 
+ bl[126] br[126] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_129 
+ bl[127] br[127] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_130 
+ bl[128] br[128] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_131 
+ bl[129] br[129] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_132 
+ bl[130] br[130] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_133 
+ bl[131] br[131] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_134 
+ bl[132] br[132] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_135 
+ bl[133] br[133] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_136 
+ bl[134] br[134] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_137 
+ bl[135] br[135] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_138 
+ bl[136] br[136] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_139 
+ bl[137] br[137] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_140 
+ bl[138] br[138] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_141 
+ bl[139] br[139] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_142 
+ bl[140] br[140] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_143 
+ bl[141] br[141] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_144 
+ bl[142] br[142] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_145 
+ bl[143] br[143] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_146 
+ bl[144] br[144] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_147 
+ bl[145] br[145] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_148 
+ bl[146] br[146] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_149 
+ bl[147] br[147] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_150 
+ bl[148] br[148] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_151 
+ bl[149] br[149] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_152 
+ bl[150] br[150] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_153 
+ bl[151] br[151] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_154 
+ bl[152] br[152] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_155 
+ bl[153] br[153] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_156 
+ bl[154] br[154] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_157 
+ bl[155] br[155] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_158 
+ bl[156] br[156] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_159 
+ bl[157] br[157] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_160 
+ bl[158] br[158] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_161 
+ bl[159] br[159] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_162 
+ bl[160] br[160] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_163 
+ bl[161] br[161] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_164 
+ bl[162] br[162] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_165 
+ bl[163] br[163] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_166 
+ bl[164] br[164] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_167 
+ bl[165] br[165] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_168 
+ bl[166] br[166] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_169 
+ bl[167] br[167] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_170 
+ bl[168] br[168] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_171 
+ bl[169] br[169] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_172 
+ bl[170] br[170] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_173 
+ bl[171] br[171] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_174 
+ bl[172] br[172] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_175 
+ bl[173] br[173] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_176 
+ bl[174] br[174] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_177 
+ bl[175] br[175] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_178 
+ bl[176] br[176] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_179 
+ bl[177] br[177] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_180 
+ bl[178] br[178] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_181 
+ bl[179] br[179] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_182 
+ bl[180] br[180] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_183 
+ bl[181] br[181] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_184 
+ bl[182] br[182] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_185 
+ bl[183] br[183] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_186 
+ bl[184] br[184] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_187 
+ bl[185] br[185] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_188 
+ bl[186] br[186] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_189 
+ bl[187] br[187] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_190 
+ bl[188] br[188] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_191 
+ bl[189] br[189] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_192 
+ bl[190] br[190] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_193 
+ bl[191] br[191] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_194 
+ bl[192] br[192] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_195 
+ bl[193] br[193] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_196 
+ bl[194] br[194] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_197 
+ bl[195] br[195] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_198 
+ bl[196] br[196] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_199 
+ bl[197] br[197] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_200 
+ bl[198] br[198] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_201 
+ bl[199] br[199] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_202 
+ bl[200] br[200] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_203 
+ bl[201] br[201] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_204 
+ bl[202] br[202] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_205 
+ bl[203] br[203] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_206 
+ bl[204] br[204] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_207 
+ bl[205] br[205] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_208 
+ bl[206] br[206] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_209 
+ bl[207] br[207] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_210 
+ bl[208] br[208] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_211 
+ bl[209] br[209] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_212 
+ bl[210] br[210] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_213 
+ bl[211] br[211] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_214 
+ bl[212] br[212] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_215 
+ bl[213] br[213] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_216 
+ bl[214] br[214] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_217 
+ bl[215] br[215] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_218 
+ bl[216] br[216] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_219 
+ bl[217] br[217] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_220 
+ bl[218] br[218] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_221 
+ bl[219] br[219] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_222 
+ bl[220] br[220] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_223 
+ bl[221] br[221] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_224 
+ bl[222] br[222] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_225 
+ bl[223] br[223] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_226 
+ bl[224] br[224] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_227 
+ bl[225] br[225] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_228 
+ bl[226] br[226] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_229 
+ bl[227] br[227] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_230 
+ bl[228] br[228] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_231 
+ bl[229] br[229] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_232 
+ bl[230] br[230] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_233 
+ bl[231] br[231] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_234 
+ bl[232] br[232] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_235 
+ bl[233] br[233] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_236 
+ bl[234] br[234] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_237 
+ bl[235] br[235] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_238 
+ bl[236] br[236] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_239 
+ bl[237] br[237] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_240 
+ bl[238] br[238] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_241 
+ bl[239] br[239] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_242 
+ bl[240] br[240] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_243 
+ bl[241] br[241] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_244 
+ bl[242] br[242] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_245 
+ bl[243] br[243] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_246 
+ bl[244] br[244] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_247 
+ bl[245] br[245] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_248 
+ bl[246] br[246] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_249 
+ bl[247] br[247] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_250 
+ bl[248] br[248] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_251 
+ bl[249] br[249] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_252 
+ bl[250] br[250] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_253 
+ bl[251] br[251] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_254 
+ bl[252] br[252] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_255 
+ bl[253] br[253] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_256 
+ bl[254] br[254] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_257 
+ bl[255] br[255] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_258 
+ vdd vdd vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_259 
+ vdd vdd vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_0 
+ vdd vdd vss vdd vpb vnb wl[111] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_113_1 
+ rbl rbr vss vdd vpb vnb wl[111] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_113_2 
+ bl[0] br[0] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_3 
+ bl[1] br[1] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_4 
+ bl[2] br[2] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_5 
+ bl[3] br[3] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_6 
+ bl[4] br[4] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_7 
+ bl[5] br[5] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_8 
+ bl[6] br[6] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_9 
+ bl[7] br[7] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_10 
+ bl[8] br[8] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_11 
+ bl[9] br[9] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_12 
+ bl[10] br[10] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_13 
+ bl[11] br[11] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_14 
+ bl[12] br[12] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_15 
+ bl[13] br[13] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_16 
+ bl[14] br[14] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_17 
+ bl[15] br[15] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_18 
+ bl[16] br[16] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_19 
+ bl[17] br[17] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_20 
+ bl[18] br[18] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_21 
+ bl[19] br[19] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_22 
+ bl[20] br[20] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_23 
+ bl[21] br[21] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_24 
+ bl[22] br[22] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_25 
+ bl[23] br[23] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_26 
+ bl[24] br[24] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_27 
+ bl[25] br[25] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_28 
+ bl[26] br[26] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_29 
+ bl[27] br[27] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_30 
+ bl[28] br[28] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_31 
+ bl[29] br[29] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_32 
+ bl[30] br[30] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_33 
+ bl[31] br[31] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_34 
+ bl[32] br[32] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_35 
+ bl[33] br[33] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_36 
+ bl[34] br[34] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_37 
+ bl[35] br[35] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_38 
+ bl[36] br[36] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_39 
+ bl[37] br[37] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_40 
+ bl[38] br[38] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_41 
+ bl[39] br[39] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_42 
+ bl[40] br[40] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_43 
+ bl[41] br[41] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_44 
+ bl[42] br[42] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_45 
+ bl[43] br[43] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_46 
+ bl[44] br[44] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_47 
+ bl[45] br[45] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_48 
+ bl[46] br[46] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_49 
+ bl[47] br[47] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_50 
+ bl[48] br[48] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_51 
+ bl[49] br[49] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_52 
+ bl[50] br[50] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_53 
+ bl[51] br[51] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_54 
+ bl[52] br[52] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_55 
+ bl[53] br[53] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_56 
+ bl[54] br[54] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_57 
+ bl[55] br[55] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_58 
+ bl[56] br[56] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_59 
+ bl[57] br[57] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_60 
+ bl[58] br[58] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_61 
+ bl[59] br[59] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_62 
+ bl[60] br[60] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_63 
+ bl[61] br[61] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_64 
+ bl[62] br[62] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_65 
+ bl[63] br[63] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_66 
+ bl[64] br[64] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_67 
+ bl[65] br[65] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_68 
+ bl[66] br[66] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_69 
+ bl[67] br[67] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_70 
+ bl[68] br[68] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_71 
+ bl[69] br[69] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_72 
+ bl[70] br[70] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_73 
+ bl[71] br[71] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_74 
+ bl[72] br[72] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_75 
+ bl[73] br[73] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_76 
+ bl[74] br[74] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_77 
+ bl[75] br[75] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_78 
+ bl[76] br[76] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_79 
+ bl[77] br[77] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_80 
+ bl[78] br[78] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_81 
+ bl[79] br[79] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_82 
+ bl[80] br[80] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_83 
+ bl[81] br[81] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_84 
+ bl[82] br[82] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_85 
+ bl[83] br[83] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_86 
+ bl[84] br[84] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_87 
+ bl[85] br[85] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_88 
+ bl[86] br[86] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_89 
+ bl[87] br[87] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_90 
+ bl[88] br[88] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_91 
+ bl[89] br[89] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_92 
+ bl[90] br[90] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_93 
+ bl[91] br[91] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_94 
+ bl[92] br[92] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_95 
+ bl[93] br[93] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_96 
+ bl[94] br[94] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_97 
+ bl[95] br[95] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_98 
+ bl[96] br[96] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_99 
+ bl[97] br[97] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_100 
+ bl[98] br[98] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_101 
+ bl[99] br[99] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_102 
+ bl[100] br[100] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_103 
+ bl[101] br[101] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_104 
+ bl[102] br[102] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_105 
+ bl[103] br[103] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_106 
+ bl[104] br[104] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_107 
+ bl[105] br[105] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_108 
+ bl[106] br[106] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_109 
+ bl[107] br[107] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_110 
+ bl[108] br[108] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_111 
+ bl[109] br[109] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_112 
+ bl[110] br[110] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_113 
+ bl[111] br[111] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_114 
+ bl[112] br[112] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_115 
+ bl[113] br[113] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_116 
+ bl[114] br[114] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_117 
+ bl[115] br[115] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_118 
+ bl[116] br[116] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_119 
+ bl[117] br[117] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_120 
+ bl[118] br[118] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_121 
+ bl[119] br[119] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_122 
+ bl[120] br[120] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_123 
+ bl[121] br[121] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_124 
+ bl[122] br[122] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_125 
+ bl[123] br[123] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_126 
+ bl[124] br[124] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_127 
+ bl[125] br[125] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_128 
+ bl[126] br[126] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_129 
+ bl[127] br[127] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_130 
+ bl[128] br[128] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_131 
+ bl[129] br[129] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_132 
+ bl[130] br[130] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_133 
+ bl[131] br[131] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_134 
+ bl[132] br[132] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_135 
+ bl[133] br[133] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_136 
+ bl[134] br[134] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_137 
+ bl[135] br[135] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_138 
+ bl[136] br[136] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_139 
+ bl[137] br[137] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_140 
+ bl[138] br[138] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_141 
+ bl[139] br[139] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_142 
+ bl[140] br[140] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_143 
+ bl[141] br[141] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_144 
+ bl[142] br[142] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_145 
+ bl[143] br[143] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_146 
+ bl[144] br[144] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_147 
+ bl[145] br[145] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_148 
+ bl[146] br[146] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_149 
+ bl[147] br[147] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_150 
+ bl[148] br[148] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_151 
+ bl[149] br[149] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_152 
+ bl[150] br[150] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_153 
+ bl[151] br[151] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_154 
+ bl[152] br[152] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_155 
+ bl[153] br[153] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_156 
+ bl[154] br[154] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_157 
+ bl[155] br[155] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_158 
+ bl[156] br[156] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_159 
+ bl[157] br[157] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_160 
+ bl[158] br[158] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_161 
+ bl[159] br[159] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_162 
+ bl[160] br[160] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_163 
+ bl[161] br[161] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_164 
+ bl[162] br[162] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_165 
+ bl[163] br[163] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_166 
+ bl[164] br[164] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_167 
+ bl[165] br[165] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_168 
+ bl[166] br[166] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_169 
+ bl[167] br[167] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_170 
+ bl[168] br[168] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_171 
+ bl[169] br[169] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_172 
+ bl[170] br[170] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_173 
+ bl[171] br[171] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_174 
+ bl[172] br[172] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_175 
+ bl[173] br[173] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_176 
+ bl[174] br[174] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_177 
+ bl[175] br[175] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_178 
+ bl[176] br[176] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_179 
+ bl[177] br[177] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_180 
+ bl[178] br[178] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_181 
+ bl[179] br[179] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_182 
+ bl[180] br[180] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_183 
+ bl[181] br[181] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_184 
+ bl[182] br[182] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_185 
+ bl[183] br[183] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_186 
+ bl[184] br[184] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_187 
+ bl[185] br[185] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_188 
+ bl[186] br[186] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_189 
+ bl[187] br[187] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_190 
+ bl[188] br[188] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_191 
+ bl[189] br[189] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_192 
+ bl[190] br[190] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_193 
+ bl[191] br[191] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_194 
+ bl[192] br[192] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_195 
+ bl[193] br[193] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_196 
+ bl[194] br[194] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_197 
+ bl[195] br[195] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_198 
+ bl[196] br[196] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_199 
+ bl[197] br[197] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_200 
+ bl[198] br[198] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_201 
+ bl[199] br[199] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_202 
+ bl[200] br[200] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_203 
+ bl[201] br[201] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_204 
+ bl[202] br[202] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_205 
+ bl[203] br[203] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_206 
+ bl[204] br[204] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_207 
+ bl[205] br[205] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_208 
+ bl[206] br[206] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_209 
+ bl[207] br[207] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_210 
+ bl[208] br[208] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_211 
+ bl[209] br[209] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_212 
+ bl[210] br[210] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_213 
+ bl[211] br[211] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_214 
+ bl[212] br[212] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_215 
+ bl[213] br[213] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_216 
+ bl[214] br[214] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_217 
+ bl[215] br[215] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_218 
+ bl[216] br[216] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_219 
+ bl[217] br[217] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_220 
+ bl[218] br[218] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_221 
+ bl[219] br[219] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_222 
+ bl[220] br[220] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_223 
+ bl[221] br[221] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_224 
+ bl[222] br[222] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_225 
+ bl[223] br[223] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_226 
+ bl[224] br[224] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_227 
+ bl[225] br[225] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_228 
+ bl[226] br[226] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_229 
+ bl[227] br[227] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_230 
+ bl[228] br[228] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_231 
+ bl[229] br[229] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_232 
+ bl[230] br[230] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_233 
+ bl[231] br[231] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_234 
+ bl[232] br[232] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_235 
+ bl[233] br[233] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_236 
+ bl[234] br[234] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_237 
+ bl[235] br[235] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_238 
+ bl[236] br[236] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_239 
+ bl[237] br[237] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_240 
+ bl[238] br[238] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_241 
+ bl[239] br[239] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_242 
+ bl[240] br[240] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_243 
+ bl[241] br[241] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_244 
+ bl[242] br[242] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_245 
+ bl[243] br[243] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_246 
+ bl[244] br[244] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_247 
+ bl[245] br[245] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_248 
+ bl[246] br[246] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_249 
+ bl[247] br[247] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_250 
+ bl[248] br[248] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_251 
+ bl[249] br[249] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_252 
+ bl[250] br[250] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_253 
+ bl[251] br[251] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_254 
+ bl[252] br[252] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_255 
+ bl[253] br[253] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_256 
+ bl[254] br[254] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_257 
+ bl[255] br[255] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_258 
+ vdd vdd vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_259 
+ vdd vdd vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_0 
+ vdd vdd vss vdd vpb vnb wl[112] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_114_1 
+ rbl rbr vss vdd vpb vnb wl[112] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_114_2 
+ bl[0] br[0] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_3 
+ bl[1] br[1] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_4 
+ bl[2] br[2] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_5 
+ bl[3] br[3] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_6 
+ bl[4] br[4] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_7 
+ bl[5] br[5] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_8 
+ bl[6] br[6] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_9 
+ bl[7] br[7] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_10 
+ bl[8] br[8] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_11 
+ bl[9] br[9] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_12 
+ bl[10] br[10] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_13 
+ bl[11] br[11] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_14 
+ bl[12] br[12] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_15 
+ bl[13] br[13] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_16 
+ bl[14] br[14] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_17 
+ bl[15] br[15] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_18 
+ bl[16] br[16] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_19 
+ bl[17] br[17] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_20 
+ bl[18] br[18] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_21 
+ bl[19] br[19] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_22 
+ bl[20] br[20] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_23 
+ bl[21] br[21] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_24 
+ bl[22] br[22] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_25 
+ bl[23] br[23] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_26 
+ bl[24] br[24] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_27 
+ bl[25] br[25] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_28 
+ bl[26] br[26] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_29 
+ bl[27] br[27] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_30 
+ bl[28] br[28] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_31 
+ bl[29] br[29] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_32 
+ bl[30] br[30] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_33 
+ bl[31] br[31] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_34 
+ bl[32] br[32] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_35 
+ bl[33] br[33] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_36 
+ bl[34] br[34] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_37 
+ bl[35] br[35] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_38 
+ bl[36] br[36] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_39 
+ bl[37] br[37] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_40 
+ bl[38] br[38] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_41 
+ bl[39] br[39] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_42 
+ bl[40] br[40] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_43 
+ bl[41] br[41] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_44 
+ bl[42] br[42] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_45 
+ bl[43] br[43] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_46 
+ bl[44] br[44] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_47 
+ bl[45] br[45] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_48 
+ bl[46] br[46] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_49 
+ bl[47] br[47] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_50 
+ bl[48] br[48] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_51 
+ bl[49] br[49] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_52 
+ bl[50] br[50] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_53 
+ bl[51] br[51] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_54 
+ bl[52] br[52] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_55 
+ bl[53] br[53] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_56 
+ bl[54] br[54] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_57 
+ bl[55] br[55] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_58 
+ bl[56] br[56] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_59 
+ bl[57] br[57] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_60 
+ bl[58] br[58] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_61 
+ bl[59] br[59] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_62 
+ bl[60] br[60] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_63 
+ bl[61] br[61] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_64 
+ bl[62] br[62] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_65 
+ bl[63] br[63] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_66 
+ bl[64] br[64] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_67 
+ bl[65] br[65] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_68 
+ bl[66] br[66] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_69 
+ bl[67] br[67] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_70 
+ bl[68] br[68] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_71 
+ bl[69] br[69] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_72 
+ bl[70] br[70] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_73 
+ bl[71] br[71] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_74 
+ bl[72] br[72] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_75 
+ bl[73] br[73] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_76 
+ bl[74] br[74] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_77 
+ bl[75] br[75] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_78 
+ bl[76] br[76] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_79 
+ bl[77] br[77] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_80 
+ bl[78] br[78] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_81 
+ bl[79] br[79] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_82 
+ bl[80] br[80] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_83 
+ bl[81] br[81] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_84 
+ bl[82] br[82] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_85 
+ bl[83] br[83] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_86 
+ bl[84] br[84] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_87 
+ bl[85] br[85] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_88 
+ bl[86] br[86] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_89 
+ bl[87] br[87] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_90 
+ bl[88] br[88] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_91 
+ bl[89] br[89] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_92 
+ bl[90] br[90] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_93 
+ bl[91] br[91] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_94 
+ bl[92] br[92] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_95 
+ bl[93] br[93] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_96 
+ bl[94] br[94] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_97 
+ bl[95] br[95] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_98 
+ bl[96] br[96] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_99 
+ bl[97] br[97] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_100 
+ bl[98] br[98] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_101 
+ bl[99] br[99] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_102 
+ bl[100] br[100] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_103 
+ bl[101] br[101] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_104 
+ bl[102] br[102] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_105 
+ bl[103] br[103] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_106 
+ bl[104] br[104] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_107 
+ bl[105] br[105] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_108 
+ bl[106] br[106] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_109 
+ bl[107] br[107] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_110 
+ bl[108] br[108] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_111 
+ bl[109] br[109] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_112 
+ bl[110] br[110] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_113 
+ bl[111] br[111] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_114 
+ bl[112] br[112] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_115 
+ bl[113] br[113] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_116 
+ bl[114] br[114] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_117 
+ bl[115] br[115] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_118 
+ bl[116] br[116] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_119 
+ bl[117] br[117] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_120 
+ bl[118] br[118] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_121 
+ bl[119] br[119] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_122 
+ bl[120] br[120] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_123 
+ bl[121] br[121] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_124 
+ bl[122] br[122] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_125 
+ bl[123] br[123] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_126 
+ bl[124] br[124] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_127 
+ bl[125] br[125] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_128 
+ bl[126] br[126] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_129 
+ bl[127] br[127] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_130 
+ bl[128] br[128] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_131 
+ bl[129] br[129] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_132 
+ bl[130] br[130] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_133 
+ bl[131] br[131] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_134 
+ bl[132] br[132] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_135 
+ bl[133] br[133] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_136 
+ bl[134] br[134] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_137 
+ bl[135] br[135] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_138 
+ bl[136] br[136] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_139 
+ bl[137] br[137] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_140 
+ bl[138] br[138] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_141 
+ bl[139] br[139] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_142 
+ bl[140] br[140] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_143 
+ bl[141] br[141] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_144 
+ bl[142] br[142] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_145 
+ bl[143] br[143] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_146 
+ bl[144] br[144] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_147 
+ bl[145] br[145] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_148 
+ bl[146] br[146] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_149 
+ bl[147] br[147] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_150 
+ bl[148] br[148] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_151 
+ bl[149] br[149] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_152 
+ bl[150] br[150] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_153 
+ bl[151] br[151] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_154 
+ bl[152] br[152] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_155 
+ bl[153] br[153] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_156 
+ bl[154] br[154] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_157 
+ bl[155] br[155] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_158 
+ bl[156] br[156] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_159 
+ bl[157] br[157] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_160 
+ bl[158] br[158] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_161 
+ bl[159] br[159] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_162 
+ bl[160] br[160] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_163 
+ bl[161] br[161] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_164 
+ bl[162] br[162] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_165 
+ bl[163] br[163] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_166 
+ bl[164] br[164] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_167 
+ bl[165] br[165] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_168 
+ bl[166] br[166] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_169 
+ bl[167] br[167] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_170 
+ bl[168] br[168] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_171 
+ bl[169] br[169] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_172 
+ bl[170] br[170] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_173 
+ bl[171] br[171] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_174 
+ bl[172] br[172] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_175 
+ bl[173] br[173] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_176 
+ bl[174] br[174] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_177 
+ bl[175] br[175] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_178 
+ bl[176] br[176] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_179 
+ bl[177] br[177] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_180 
+ bl[178] br[178] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_181 
+ bl[179] br[179] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_182 
+ bl[180] br[180] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_183 
+ bl[181] br[181] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_184 
+ bl[182] br[182] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_185 
+ bl[183] br[183] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_186 
+ bl[184] br[184] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_187 
+ bl[185] br[185] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_188 
+ bl[186] br[186] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_189 
+ bl[187] br[187] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_190 
+ bl[188] br[188] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_191 
+ bl[189] br[189] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_192 
+ bl[190] br[190] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_193 
+ bl[191] br[191] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_194 
+ bl[192] br[192] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_195 
+ bl[193] br[193] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_196 
+ bl[194] br[194] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_197 
+ bl[195] br[195] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_198 
+ bl[196] br[196] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_199 
+ bl[197] br[197] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_200 
+ bl[198] br[198] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_201 
+ bl[199] br[199] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_202 
+ bl[200] br[200] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_203 
+ bl[201] br[201] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_204 
+ bl[202] br[202] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_205 
+ bl[203] br[203] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_206 
+ bl[204] br[204] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_207 
+ bl[205] br[205] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_208 
+ bl[206] br[206] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_209 
+ bl[207] br[207] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_210 
+ bl[208] br[208] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_211 
+ bl[209] br[209] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_212 
+ bl[210] br[210] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_213 
+ bl[211] br[211] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_214 
+ bl[212] br[212] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_215 
+ bl[213] br[213] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_216 
+ bl[214] br[214] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_217 
+ bl[215] br[215] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_218 
+ bl[216] br[216] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_219 
+ bl[217] br[217] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_220 
+ bl[218] br[218] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_221 
+ bl[219] br[219] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_222 
+ bl[220] br[220] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_223 
+ bl[221] br[221] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_224 
+ bl[222] br[222] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_225 
+ bl[223] br[223] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_226 
+ bl[224] br[224] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_227 
+ bl[225] br[225] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_228 
+ bl[226] br[226] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_229 
+ bl[227] br[227] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_230 
+ bl[228] br[228] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_231 
+ bl[229] br[229] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_232 
+ bl[230] br[230] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_233 
+ bl[231] br[231] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_234 
+ bl[232] br[232] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_235 
+ bl[233] br[233] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_236 
+ bl[234] br[234] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_237 
+ bl[235] br[235] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_238 
+ bl[236] br[236] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_239 
+ bl[237] br[237] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_240 
+ bl[238] br[238] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_241 
+ bl[239] br[239] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_242 
+ bl[240] br[240] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_243 
+ bl[241] br[241] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_244 
+ bl[242] br[242] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_245 
+ bl[243] br[243] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_246 
+ bl[244] br[244] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_247 
+ bl[245] br[245] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_248 
+ bl[246] br[246] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_249 
+ bl[247] br[247] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_250 
+ bl[248] br[248] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_251 
+ bl[249] br[249] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_252 
+ bl[250] br[250] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_253 
+ bl[251] br[251] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_254 
+ bl[252] br[252] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_255 
+ bl[253] br[253] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_256 
+ bl[254] br[254] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_257 
+ bl[255] br[255] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_258 
+ vdd vdd vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_259 
+ vdd vdd vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_0 
+ vdd vdd vss vdd vpb vnb wl[113] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_115_1 
+ rbl rbr vss vdd vpb vnb wl[113] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_115_2 
+ bl[0] br[0] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_3 
+ bl[1] br[1] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_4 
+ bl[2] br[2] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_5 
+ bl[3] br[3] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_6 
+ bl[4] br[4] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_7 
+ bl[5] br[5] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_8 
+ bl[6] br[6] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_9 
+ bl[7] br[7] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_10 
+ bl[8] br[8] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_11 
+ bl[9] br[9] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_12 
+ bl[10] br[10] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_13 
+ bl[11] br[11] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_14 
+ bl[12] br[12] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_15 
+ bl[13] br[13] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_16 
+ bl[14] br[14] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_17 
+ bl[15] br[15] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_18 
+ bl[16] br[16] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_19 
+ bl[17] br[17] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_20 
+ bl[18] br[18] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_21 
+ bl[19] br[19] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_22 
+ bl[20] br[20] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_23 
+ bl[21] br[21] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_24 
+ bl[22] br[22] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_25 
+ bl[23] br[23] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_26 
+ bl[24] br[24] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_27 
+ bl[25] br[25] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_28 
+ bl[26] br[26] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_29 
+ bl[27] br[27] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_30 
+ bl[28] br[28] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_31 
+ bl[29] br[29] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_32 
+ bl[30] br[30] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_33 
+ bl[31] br[31] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_34 
+ bl[32] br[32] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_35 
+ bl[33] br[33] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_36 
+ bl[34] br[34] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_37 
+ bl[35] br[35] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_38 
+ bl[36] br[36] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_39 
+ bl[37] br[37] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_40 
+ bl[38] br[38] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_41 
+ bl[39] br[39] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_42 
+ bl[40] br[40] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_43 
+ bl[41] br[41] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_44 
+ bl[42] br[42] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_45 
+ bl[43] br[43] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_46 
+ bl[44] br[44] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_47 
+ bl[45] br[45] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_48 
+ bl[46] br[46] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_49 
+ bl[47] br[47] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_50 
+ bl[48] br[48] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_51 
+ bl[49] br[49] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_52 
+ bl[50] br[50] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_53 
+ bl[51] br[51] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_54 
+ bl[52] br[52] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_55 
+ bl[53] br[53] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_56 
+ bl[54] br[54] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_57 
+ bl[55] br[55] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_58 
+ bl[56] br[56] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_59 
+ bl[57] br[57] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_60 
+ bl[58] br[58] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_61 
+ bl[59] br[59] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_62 
+ bl[60] br[60] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_63 
+ bl[61] br[61] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_64 
+ bl[62] br[62] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_65 
+ bl[63] br[63] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_66 
+ bl[64] br[64] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_67 
+ bl[65] br[65] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_68 
+ bl[66] br[66] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_69 
+ bl[67] br[67] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_70 
+ bl[68] br[68] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_71 
+ bl[69] br[69] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_72 
+ bl[70] br[70] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_73 
+ bl[71] br[71] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_74 
+ bl[72] br[72] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_75 
+ bl[73] br[73] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_76 
+ bl[74] br[74] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_77 
+ bl[75] br[75] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_78 
+ bl[76] br[76] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_79 
+ bl[77] br[77] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_80 
+ bl[78] br[78] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_81 
+ bl[79] br[79] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_82 
+ bl[80] br[80] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_83 
+ bl[81] br[81] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_84 
+ bl[82] br[82] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_85 
+ bl[83] br[83] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_86 
+ bl[84] br[84] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_87 
+ bl[85] br[85] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_88 
+ bl[86] br[86] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_89 
+ bl[87] br[87] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_90 
+ bl[88] br[88] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_91 
+ bl[89] br[89] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_92 
+ bl[90] br[90] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_93 
+ bl[91] br[91] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_94 
+ bl[92] br[92] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_95 
+ bl[93] br[93] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_96 
+ bl[94] br[94] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_97 
+ bl[95] br[95] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_98 
+ bl[96] br[96] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_99 
+ bl[97] br[97] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_100 
+ bl[98] br[98] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_101 
+ bl[99] br[99] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_102 
+ bl[100] br[100] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_103 
+ bl[101] br[101] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_104 
+ bl[102] br[102] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_105 
+ bl[103] br[103] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_106 
+ bl[104] br[104] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_107 
+ bl[105] br[105] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_108 
+ bl[106] br[106] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_109 
+ bl[107] br[107] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_110 
+ bl[108] br[108] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_111 
+ bl[109] br[109] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_112 
+ bl[110] br[110] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_113 
+ bl[111] br[111] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_114 
+ bl[112] br[112] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_115 
+ bl[113] br[113] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_116 
+ bl[114] br[114] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_117 
+ bl[115] br[115] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_118 
+ bl[116] br[116] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_119 
+ bl[117] br[117] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_120 
+ bl[118] br[118] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_121 
+ bl[119] br[119] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_122 
+ bl[120] br[120] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_123 
+ bl[121] br[121] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_124 
+ bl[122] br[122] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_125 
+ bl[123] br[123] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_126 
+ bl[124] br[124] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_127 
+ bl[125] br[125] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_128 
+ bl[126] br[126] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_129 
+ bl[127] br[127] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_130 
+ bl[128] br[128] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_131 
+ bl[129] br[129] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_132 
+ bl[130] br[130] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_133 
+ bl[131] br[131] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_134 
+ bl[132] br[132] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_135 
+ bl[133] br[133] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_136 
+ bl[134] br[134] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_137 
+ bl[135] br[135] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_138 
+ bl[136] br[136] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_139 
+ bl[137] br[137] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_140 
+ bl[138] br[138] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_141 
+ bl[139] br[139] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_142 
+ bl[140] br[140] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_143 
+ bl[141] br[141] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_144 
+ bl[142] br[142] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_145 
+ bl[143] br[143] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_146 
+ bl[144] br[144] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_147 
+ bl[145] br[145] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_148 
+ bl[146] br[146] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_149 
+ bl[147] br[147] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_150 
+ bl[148] br[148] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_151 
+ bl[149] br[149] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_152 
+ bl[150] br[150] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_153 
+ bl[151] br[151] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_154 
+ bl[152] br[152] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_155 
+ bl[153] br[153] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_156 
+ bl[154] br[154] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_157 
+ bl[155] br[155] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_158 
+ bl[156] br[156] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_159 
+ bl[157] br[157] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_160 
+ bl[158] br[158] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_161 
+ bl[159] br[159] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_162 
+ bl[160] br[160] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_163 
+ bl[161] br[161] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_164 
+ bl[162] br[162] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_165 
+ bl[163] br[163] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_166 
+ bl[164] br[164] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_167 
+ bl[165] br[165] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_168 
+ bl[166] br[166] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_169 
+ bl[167] br[167] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_170 
+ bl[168] br[168] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_171 
+ bl[169] br[169] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_172 
+ bl[170] br[170] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_173 
+ bl[171] br[171] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_174 
+ bl[172] br[172] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_175 
+ bl[173] br[173] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_176 
+ bl[174] br[174] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_177 
+ bl[175] br[175] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_178 
+ bl[176] br[176] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_179 
+ bl[177] br[177] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_180 
+ bl[178] br[178] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_181 
+ bl[179] br[179] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_182 
+ bl[180] br[180] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_183 
+ bl[181] br[181] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_184 
+ bl[182] br[182] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_185 
+ bl[183] br[183] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_186 
+ bl[184] br[184] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_187 
+ bl[185] br[185] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_188 
+ bl[186] br[186] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_189 
+ bl[187] br[187] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_190 
+ bl[188] br[188] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_191 
+ bl[189] br[189] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_192 
+ bl[190] br[190] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_193 
+ bl[191] br[191] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_194 
+ bl[192] br[192] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_195 
+ bl[193] br[193] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_196 
+ bl[194] br[194] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_197 
+ bl[195] br[195] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_198 
+ bl[196] br[196] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_199 
+ bl[197] br[197] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_200 
+ bl[198] br[198] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_201 
+ bl[199] br[199] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_202 
+ bl[200] br[200] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_203 
+ bl[201] br[201] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_204 
+ bl[202] br[202] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_205 
+ bl[203] br[203] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_206 
+ bl[204] br[204] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_207 
+ bl[205] br[205] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_208 
+ bl[206] br[206] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_209 
+ bl[207] br[207] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_210 
+ bl[208] br[208] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_211 
+ bl[209] br[209] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_212 
+ bl[210] br[210] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_213 
+ bl[211] br[211] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_214 
+ bl[212] br[212] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_215 
+ bl[213] br[213] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_216 
+ bl[214] br[214] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_217 
+ bl[215] br[215] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_218 
+ bl[216] br[216] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_219 
+ bl[217] br[217] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_220 
+ bl[218] br[218] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_221 
+ bl[219] br[219] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_222 
+ bl[220] br[220] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_223 
+ bl[221] br[221] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_224 
+ bl[222] br[222] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_225 
+ bl[223] br[223] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_226 
+ bl[224] br[224] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_227 
+ bl[225] br[225] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_228 
+ bl[226] br[226] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_229 
+ bl[227] br[227] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_230 
+ bl[228] br[228] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_231 
+ bl[229] br[229] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_232 
+ bl[230] br[230] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_233 
+ bl[231] br[231] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_234 
+ bl[232] br[232] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_235 
+ bl[233] br[233] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_236 
+ bl[234] br[234] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_237 
+ bl[235] br[235] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_238 
+ bl[236] br[236] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_239 
+ bl[237] br[237] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_240 
+ bl[238] br[238] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_241 
+ bl[239] br[239] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_242 
+ bl[240] br[240] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_243 
+ bl[241] br[241] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_244 
+ bl[242] br[242] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_245 
+ bl[243] br[243] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_246 
+ bl[244] br[244] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_247 
+ bl[245] br[245] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_248 
+ bl[246] br[246] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_249 
+ bl[247] br[247] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_250 
+ bl[248] br[248] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_251 
+ bl[249] br[249] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_252 
+ bl[250] br[250] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_253 
+ bl[251] br[251] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_254 
+ bl[252] br[252] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_255 
+ bl[253] br[253] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_256 
+ bl[254] br[254] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_257 
+ bl[255] br[255] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_258 
+ vdd vdd vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_259 
+ vdd vdd vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_0 
+ vdd vdd vss vdd vpb vnb wl[114] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_116_1 
+ rbl rbr vss vdd vpb vnb wl[114] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_116_2 
+ bl[0] br[0] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_3 
+ bl[1] br[1] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_4 
+ bl[2] br[2] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_5 
+ bl[3] br[3] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_6 
+ bl[4] br[4] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_7 
+ bl[5] br[5] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_8 
+ bl[6] br[6] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_9 
+ bl[7] br[7] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_10 
+ bl[8] br[8] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_11 
+ bl[9] br[9] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_12 
+ bl[10] br[10] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_13 
+ bl[11] br[11] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_14 
+ bl[12] br[12] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_15 
+ bl[13] br[13] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_16 
+ bl[14] br[14] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_17 
+ bl[15] br[15] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_18 
+ bl[16] br[16] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_19 
+ bl[17] br[17] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_20 
+ bl[18] br[18] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_21 
+ bl[19] br[19] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_22 
+ bl[20] br[20] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_23 
+ bl[21] br[21] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_24 
+ bl[22] br[22] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_25 
+ bl[23] br[23] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_26 
+ bl[24] br[24] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_27 
+ bl[25] br[25] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_28 
+ bl[26] br[26] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_29 
+ bl[27] br[27] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_30 
+ bl[28] br[28] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_31 
+ bl[29] br[29] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_32 
+ bl[30] br[30] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_33 
+ bl[31] br[31] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_34 
+ bl[32] br[32] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_35 
+ bl[33] br[33] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_36 
+ bl[34] br[34] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_37 
+ bl[35] br[35] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_38 
+ bl[36] br[36] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_39 
+ bl[37] br[37] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_40 
+ bl[38] br[38] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_41 
+ bl[39] br[39] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_42 
+ bl[40] br[40] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_43 
+ bl[41] br[41] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_44 
+ bl[42] br[42] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_45 
+ bl[43] br[43] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_46 
+ bl[44] br[44] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_47 
+ bl[45] br[45] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_48 
+ bl[46] br[46] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_49 
+ bl[47] br[47] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_50 
+ bl[48] br[48] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_51 
+ bl[49] br[49] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_52 
+ bl[50] br[50] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_53 
+ bl[51] br[51] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_54 
+ bl[52] br[52] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_55 
+ bl[53] br[53] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_56 
+ bl[54] br[54] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_57 
+ bl[55] br[55] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_58 
+ bl[56] br[56] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_59 
+ bl[57] br[57] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_60 
+ bl[58] br[58] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_61 
+ bl[59] br[59] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_62 
+ bl[60] br[60] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_63 
+ bl[61] br[61] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_64 
+ bl[62] br[62] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_65 
+ bl[63] br[63] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_66 
+ bl[64] br[64] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_67 
+ bl[65] br[65] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_68 
+ bl[66] br[66] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_69 
+ bl[67] br[67] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_70 
+ bl[68] br[68] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_71 
+ bl[69] br[69] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_72 
+ bl[70] br[70] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_73 
+ bl[71] br[71] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_74 
+ bl[72] br[72] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_75 
+ bl[73] br[73] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_76 
+ bl[74] br[74] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_77 
+ bl[75] br[75] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_78 
+ bl[76] br[76] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_79 
+ bl[77] br[77] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_80 
+ bl[78] br[78] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_81 
+ bl[79] br[79] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_82 
+ bl[80] br[80] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_83 
+ bl[81] br[81] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_84 
+ bl[82] br[82] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_85 
+ bl[83] br[83] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_86 
+ bl[84] br[84] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_87 
+ bl[85] br[85] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_88 
+ bl[86] br[86] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_89 
+ bl[87] br[87] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_90 
+ bl[88] br[88] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_91 
+ bl[89] br[89] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_92 
+ bl[90] br[90] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_93 
+ bl[91] br[91] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_94 
+ bl[92] br[92] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_95 
+ bl[93] br[93] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_96 
+ bl[94] br[94] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_97 
+ bl[95] br[95] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_98 
+ bl[96] br[96] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_99 
+ bl[97] br[97] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_100 
+ bl[98] br[98] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_101 
+ bl[99] br[99] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_102 
+ bl[100] br[100] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_103 
+ bl[101] br[101] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_104 
+ bl[102] br[102] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_105 
+ bl[103] br[103] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_106 
+ bl[104] br[104] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_107 
+ bl[105] br[105] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_108 
+ bl[106] br[106] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_109 
+ bl[107] br[107] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_110 
+ bl[108] br[108] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_111 
+ bl[109] br[109] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_112 
+ bl[110] br[110] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_113 
+ bl[111] br[111] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_114 
+ bl[112] br[112] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_115 
+ bl[113] br[113] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_116 
+ bl[114] br[114] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_117 
+ bl[115] br[115] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_118 
+ bl[116] br[116] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_119 
+ bl[117] br[117] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_120 
+ bl[118] br[118] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_121 
+ bl[119] br[119] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_122 
+ bl[120] br[120] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_123 
+ bl[121] br[121] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_124 
+ bl[122] br[122] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_125 
+ bl[123] br[123] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_126 
+ bl[124] br[124] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_127 
+ bl[125] br[125] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_128 
+ bl[126] br[126] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_129 
+ bl[127] br[127] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_130 
+ bl[128] br[128] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_131 
+ bl[129] br[129] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_132 
+ bl[130] br[130] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_133 
+ bl[131] br[131] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_134 
+ bl[132] br[132] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_135 
+ bl[133] br[133] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_136 
+ bl[134] br[134] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_137 
+ bl[135] br[135] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_138 
+ bl[136] br[136] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_139 
+ bl[137] br[137] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_140 
+ bl[138] br[138] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_141 
+ bl[139] br[139] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_142 
+ bl[140] br[140] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_143 
+ bl[141] br[141] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_144 
+ bl[142] br[142] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_145 
+ bl[143] br[143] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_146 
+ bl[144] br[144] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_147 
+ bl[145] br[145] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_148 
+ bl[146] br[146] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_149 
+ bl[147] br[147] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_150 
+ bl[148] br[148] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_151 
+ bl[149] br[149] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_152 
+ bl[150] br[150] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_153 
+ bl[151] br[151] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_154 
+ bl[152] br[152] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_155 
+ bl[153] br[153] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_156 
+ bl[154] br[154] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_157 
+ bl[155] br[155] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_158 
+ bl[156] br[156] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_159 
+ bl[157] br[157] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_160 
+ bl[158] br[158] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_161 
+ bl[159] br[159] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_162 
+ bl[160] br[160] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_163 
+ bl[161] br[161] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_164 
+ bl[162] br[162] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_165 
+ bl[163] br[163] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_166 
+ bl[164] br[164] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_167 
+ bl[165] br[165] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_168 
+ bl[166] br[166] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_169 
+ bl[167] br[167] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_170 
+ bl[168] br[168] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_171 
+ bl[169] br[169] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_172 
+ bl[170] br[170] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_173 
+ bl[171] br[171] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_174 
+ bl[172] br[172] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_175 
+ bl[173] br[173] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_176 
+ bl[174] br[174] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_177 
+ bl[175] br[175] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_178 
+ bl[176] br[176] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_179 
+ bl[177] br[177] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_180 
+ bl[178] br[178] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_181 
+ bl[179] br[179] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_182 
+ bl[180] br[180] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_183 
+ bl[181] br[181] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_184 
+ bl[182] br[182] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_185 
+ bl[183] br[183] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_186 
+ bl[184] br[184] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_187 
+ bl[185] br[185] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_188 
+ bl[186] br[186] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_189 
+ bl[187] br[187] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_190 
+ bl[188] br[188] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_191 
+ bl[189] br[189] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_192 
+ bl[190] br[190] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_193 
+ bl[191] br[191] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_194 
+ bl[192] br[192] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_195 
+ bl[193] br[193] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_196 
+ bl[194] br[194] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_197 
+ bl[195] br[195] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_198 
+ bl[196] br[196] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_199 
+ bl[197] br[197] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_200 
+ bl[198] br[198] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_201 
+ bl[199] br[199] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_202 
+ bl[200] br[200] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_203 
+ bl[201] br[201] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_204 
+ bl[202] br[202] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_205 
+ bl[203] br[203] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_206 
+ bl[204] br[204] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_207 
+ bl[205] br[205] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_208 
+ bl[206] br[206] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_209 
+ bl[207] br[207] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_210 
+ bl[208] br[208] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_211 
+ bl[209] br[209] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_212 
+ bl[210] br[210] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_213 
+ bl[211] br[211] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_214 
+ bl[212] br[212] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_215 
+ bl[213] br[213] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_216 
+ bl[214] br[214] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_217 
+ bl[215] br[215] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_218 
+ bl[216] br[216] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_219 
+ bl[217] br[217] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_220 
+ bl[218] br[218] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_221 
+ bl[219] br[219] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_222 
+ bl[220] br[220] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_223 
+ bl[221] br[221] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_224 
+ bl[222] br[222] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_225 
+ bl[223] br[223] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_226 
+ bl[224] br[224] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_227 
+ bl[225] br[225] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_228 
+ bl[226] br[226] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_229 
+ bl[227] br[227] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_230 
+ bl[228] br[228] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_231 
+ bl[229] br[229] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_232 
+ bl[230] br[230] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_233 
+ bl[231] br[231] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_234 
+ bl[232] br[232] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_235 
+ bl[233] br[233] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_236 
+ bl[234] br[234] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_237 
+ bl[235] br[235] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_238 
+ bl[236] br[236] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_239 
+ bl[237] br[237] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_240 
+ bl[238] br[238] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_241 
+ bl[239] br[239] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_242 
+ bl[240] br[240] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_243 
+ bl[241] br[241] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_244 
+ bl[242] br[242] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_245 
+ bl[243] br[243] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_246 
+ bl[244] br[244] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_247 
+ bl[245] br[245] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_248 
+ bl[246] br[246] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_249 
+ bl[247] br[247] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_250 
+ bl[248] br[248] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_251 
+ bl[249] br[249] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_252 
+ bl[250] br[250] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_253 
+ bl[251] br[251] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_254 
+ bl[252] br[252] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_255 
+ bl[253] br[253] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_256 
+ bl[254] br[254] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_257 
+ bl[255] br[255] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_258 
+ vdd vdd vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_259 
+ vdd vdd vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_0 
+ vdd vdd vss vdd vpb vnb wl[115] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_117_1 
+ rbl rbr vss vdd vpb vnb wl[115] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_117_2 
+ bl[0] br[0] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_3 
+ bl[1] br[1] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_4 
+ bl[2] br[2] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_5 
+ bl[3] br[3] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_6 
+ bl[4] br[4] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_7 
+ bl[5] br[5] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_8 
+ bl[6] br[6] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_9 
+ bl[7] br[7] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_10 
+ bl[8] br[8] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_11 
+ bl[9] br[9] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_12 
+ bl[10] br[10] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_13 
+ bl[11] br[11] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_14 
+ bl[12] br[12] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_15 
+ bl[13] br[13] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_16 
+ bl[14] br[14] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_17 
+ bl[15] br[15] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_18 
+ bl[16] br[16] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_19 
+ bl[17] br[17] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_20 
+ bl[18] br[18] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_21 
+ bl[19] br[19] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_22 
+ bl[20] br[20] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_23 
+ bl[21] br[21] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_24 
+ bl[22] br[22] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_25 
+ bl[23] br[23] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_26 
+ bl[24] br[24] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_27 
+ bl[25] br[25] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_28 
+ bl[26] br[26] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_29 
+ bl[27] br[27] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_30 
+ bl[28] br[28] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_31 
+ bl[29] br[29] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_32 
+ bl[30] br[30] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_33 
+ bl[31] br[31] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_34 
+ bl[32] br[32] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_35 
+ bl[33] br[33] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_36 
+ bl[34] br[34] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_37 
+ bl[35] br[35] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_38 
+ bl[36] br[36] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_39 
+ bl[37] br[37] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_40 
+ bl[38] br[38] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_41 
+ bl[39] br[39] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_42 
+ bl[40] br[40] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_43 
+ bl[41] br[41] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_44 
+ bl[42] br[42] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_45 
+ bl[43] br[43] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_46 
+ bl[44] br[44] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_47 
+ bl[45] br[45] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_48 
+ bl[46] br[46] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_49 
+ bl[47] br[47] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_50 
+ bl[48] br[48] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_51 
+ bl[49] br[49] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_52 
+ bl[50] br[50] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_53 
+ bl[51] br[51] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_54 
+ bl[52] br[52] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_55 
+ bl[53] br[53] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_56 
+ bl[54] br[54] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_57 
+ bl[55] br[55] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_58 
+ bl[56] br[56] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_59 
+ bl[57] br[57] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_60 
+ bl[58] br[58] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_61 
+ bl[59] br[59] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_62 
+ bl[60] br[60] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_63 
+ bl[61] br[61] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_64 
+ bl[62] br[62] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_65 
+ bl[63] br[63] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_66 
+ bl[64] br[64] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_67 
+ bl[65] br[65] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_68 
+ bl[66] br[66] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_69 
+ bl[67] br[67] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_70 
+ bl[68] br[68] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_71 
+ bl[69] br[69] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_72 
+ bl[70] br[70] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_73 
+ bl[71] br[71] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_74 
+ bl[72] br[72] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_75 
+ bl[73] br[73] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_76 
+ bl[74] br[74] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_77 
+ bl[75] br[75] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_78 
+ bl[76] br[76] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_79 
+ bl[77] br[77] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_80 
+ bl[78] br[78] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_81 
+ bl[79] br[79] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_82 
+ bl[80] br[80] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_83 
+ bl[81] br[81] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_84 
+ bl[82] br[82] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_85 
+ bl[83] br[83] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_86 
+ bl[84] br[84] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_87 
+ bl[85] br[85] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_88 
+ bl[86] br[86] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_89 
+ bl[87] br[87] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_90 
+ bl[88] br[88] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_91 
+ bl[89] br[89] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_92 
+ bl[90] br[90] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_93 
+ bl[91] br[91] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_94 
+ bl[92] br[92] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_95 
+ bl[93] br[93] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_96 
+ bl[94] br[94] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_97 
+ bl[95] br[95] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_98 
+ bl[96] br[96] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_99 
+ bl[97] br[97] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_100 
+ bl[98] br[98] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_101 
+ bl[99] br[99] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_102 
+ bl[100] br[100] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_103 
+ bl[101] br[101] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_104 
+ bl[102] br[102] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_105 
+ bl[103] br[103] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_106 
+ bl[104] br[104] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_107 
+ bl[105] br[105] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_108 
+ bl[106] br[106] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_109 
+ bl[107] br[107] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_110 
+ bl[108] br[108] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_111 
+ bl[109] br[109] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_112 
+ bl[110] br[110] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_113 
+ bl[111] br[111] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_114 
+ bl[112] br[112] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_115 
+ bl[113] br[113] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_116 
+ bl[114] br[114] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_117 
+ bl[115] br[115] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_118 
+ bl[116] br[116] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_119 
+ bl[117] br[117] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_120 
+ bl[118] br[118] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_121 
+ bl[119] br[119] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_122 
+ bl[120] br[120] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_123 
+ bl[121] br[121] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_124 
+ bl[122] br[122] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_125 
+ bl[123] br[123] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_126 
+ bl[124] br[124] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_127 
+ bl[125] br[125] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_128 
+ bl[126] br[126] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_129 
+ bl[127] br[127] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_130 
+ bl[128] br[128] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_131 
+ bl[129] br[129] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_132 
+ bl[130] br[130] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_133 
+ bl[131] br[131] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_134 
+ bl[132] br[132] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_135 
+ bl[133] br[133] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_136 
+ bl[134] br[134] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_137 
+ bl[135] br[135] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_138 
+ bl[136] br[136] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_139 
+ bl[137] br[137] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_140 
+ bl[138] br[138] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_141 
+ bl[139] br[139] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_142 
+ bl[140] br[140] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_143 
+ bl[141] br[141] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_144 
+ bl[142] br[142] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_145 
+ bl[143] br[143] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_146 
+ bl[144] br[144] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_147 
+ bl[145] br[145] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_148 
+ bl[146] br[146] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_149 
+ bl[147] br[147] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_150 
+ bl[148] br[148] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_151 
+ bl[149] br[149] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_152 
+ bl[150] br[150] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_153 
+ bl[151] br[151] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_154 
+ bl[152] br[152] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_155 
+ bl[153] br[153] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_156 
+ bl[154] br[154] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_157 
+ bl[155] br[155] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_158 
+ bl[156] br[156] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_159 
+ bl[157] br[157] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_160 
+ bl[158] br[158] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_161 
+ bl[159] br[159] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_162 
+ bl[160] br[160] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_163 
+ bl[161] br[161] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_164 
+ bl[162] br[162] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_165 
+ bl[163] br[163] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_166 
+ bl[164] br[164] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_167 
+ bl[165] br[165] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_168 
+ bl[166] br[166] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_169 
+ bl[167] br[167] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_170 
+ bl[168] br[168] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_171 
+ bl[169] br[169] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_172 
+ bl[170] br[170] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_173 
+ bl[171] br[171] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_174 
+ bl[172] br[172] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_175 
+ bl[173] br[173] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_176 
+ bl[174] br[174] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_177 
+ bl[175] br[175] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_178 
+ bl[176] br[176] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_179 
+ bl[177] br[177] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_180 
+ bl[178] br[178] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_181 
+ bl[179] br[179] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_182 
+ bl[180] br[180] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_183 
+ bl[181] br[181] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_184 
+ bl[182] br[182] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_185 
+ bl[183] br[183] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_186 
+ bl[184] br[184] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_187 
+ bl[185] br[185] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_188 
+ bl[186] br[186] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_189 
+ bl[187] br[187] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_190 
+ bl[188] br[188] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_191 
+ bl[189] br[189] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_192 
+ bl[190] br[190] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_193 
+ bl[191] br[191] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_194 
+ bl[192] br[192] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_195 
+ bl[193] br[193] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_196 
+ bl[194] br[194] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_197 
+ bl[195] br[195] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_198 
+ bl[196] br[196] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_199 
+ bl[197] br[197] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_200 
+ bl[198] br[198] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_201 
+ bl[199] br[199] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_202 
+ bl[200] br[200] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_203 
+ bl[201] br[201] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_204 
+ bl[202] br[202] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_205 
+ bl[203] br[203] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_206 
+ bl[204] br[204] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_207 
+ bl[205] br[205] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_208 
+ bl[206] br[206] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_209 
+ bl[207] br[207] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_210 
+ bl[208] br[208] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_211 
+ bl[209] br[209] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_212 
+ bl[210] br[210] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_213 
+ bl[211] br[211] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_214 
+ bl[212] br[212] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_215 
+ bl[213] br[213] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_216 
+ bl[214] br[214] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_217 
+ bl[215] br[215] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_218 
+ bl[216] br[216] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_219 
+ bl[217] br[217] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_220 
+ bl[218] br[218] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_221 
+ bl[219] br[219] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_222 
+ bl[220] br[220] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_223 
+ bl[221] br[221] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_224 
+ bl[222] br[222] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_225 
+ bl[223] br[223] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_226 
+ bl[224] br[224] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_227 
+ bl[225] br[225] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_228 
+ bl[226] br[226] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_229 
+ bl[227] br[227] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_230 
+ bl[228] br[228] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_231 
+ bl[229] br[229] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_232 
+ bl[230] br[230] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_233 
+ bl[231] br[231] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_234 
+ bl[232] br[232] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_235 
+ bl[233] br[233] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_236 
+ bl[234] br[234] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_237 
+ bl[235] br[235] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_238 
+ bl[236] br[236] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_239 
+ bl[237] br[237] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_240 
+ bl[238] br[238] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_241 
+ bl[239] br[239] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_242 
+ bl[240] br[240] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_243 
+ bl[241] br[241] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_244 
+ bl[242] br[242] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_245 
+ bl[243] br[243] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_246 
+ bl[244] br[244] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_247 
+ bl[245] br[245] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_248 
+ bl[246] br[246] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_249 
+ bl[247] br[247] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_250 
+ bl[248] br[248] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_251 
+ bl[249] br[249] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_252 
+ bl[250] br[250] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_253 
+ bl[251] br[251] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_254 
+ bl[252] br[252] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_255 
+ bl[253] br[253] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_256 
+ bl[254] br[254] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_257 
+ bl[255] br[255] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_258 
+ vdd vdd vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_259 
+ vdd vdd vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_0 
+ vdd vdd vss vdd vpb vnb wl[116] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_118_1 
+ rbl rbr vss vdd vpb vnb wl[116] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_118_2 
+ bl[0] br[0] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_3 
+ bl[1] br[1] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_4 
+ bl[2] br[2] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_5 
+ bl[3] br[3] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_6 
+ bl[4] br[4] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_7 
+ bl[5] br[5] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_8 
+ bl[6] br[6] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_9 
+ bl[7] br[7] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_10 
+ bl[8] br[8] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_11 
+ bl[9] br[9] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_12 
+ bl[10] br[10] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_13 
+ bl[11] br[11] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_14 
+ bl[12] br[12] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_15 
+ bl[13] br[13] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_16 
+ bl[14] br[14] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_17 
+ bl[15] br[15] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_18 
+ bl[16] br[16] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_19 
+ bl[17] br[17] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_20 
+ bl[18] br[18] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_21 
+ bl[19] br[19] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_22 
+ bl[20] br[20] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_23 
+ bl[21] br[21] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_24 
+ bl[22] br[22] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_25 
+ bl[23] br[23] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_26 
+ bl[24] br[24] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_27 
+ bl[25] br[25] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_28 
+ bl[26] br[26] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_29 
+ bl[27] br[27] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_30 
+ bl[28] br[28] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_31 
+ bl[29] br[29] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_32 
+ bl[30] br[30] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_33 
+ bl[31] br[31] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_34 
+ bl[32] br[32] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_35 
+ bl[33] br[33] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_36 
+ bl[34] br[34] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_37 
+ bl[35] br[35] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_38 
+ bl[36] br[36] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_39 
+ bl[37] br[37] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_40 
+ bl[38] br[38] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_41 
+ bl[39] br[39] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_42 
+ bl[40] br[40] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_43 
+ bl[41] br[41] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_44 
+ bl[42] br[42] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_45 
+ bl[43] br[43] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_46 
+ bl[44] br[44] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_47 
+ bl[45] br[45] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_48 
+ bl[46] br[46] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_49 
+ bl[47] br[47] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_50 
+ bl[48] br[48] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_51 
+ bl[49] br[49] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_52 
+ bl[50] br[50] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_53 
+ bl[51] br[51] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_54 
+ bl[52] br[52] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_55 
+ bl[53] br[53] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_56 
+ bl[54] br[54] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_57 
+ bl[55] br[55] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_58 
+ bl[56] br[56] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_59 
+ bl[57] br[57] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_60 
+ bl[58] br[58] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_61 
+ bl[59] br[59] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_62 
+ bl[60] br[60] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_63 
+ bl[61] br[61] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_64 
+ bl[62] br[62] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_65 
+ bl[63] br[63] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_66 
+ bl[64] br[64] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_67 
+ bl[65] br[65] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_68 
+ bl[66] br[66] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_69 
+ bl[67] br[67] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_70 
+ bl[68] br[68] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_71 
+ bl[69] br[69] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_72 
+ bl[70] br[70] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_73 
+ bl[71] br[71] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_74 
+ bl[72] br[72] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_75 
+ bl[73] br[73] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_76 
+ bl[74] br[74] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_77 
+ bl[75] br[75] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_78 
+ bl[76] br[76] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_79 
+ bl[77] br[77] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_80 
+ bl[78] br[78] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_81 
+ bl[79] br[79] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_82 
+ bl[80] br[80] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_83 
+ bl[81] br[81] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_84 
+ bl[82] br[82] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_85 
+ bl[83] br[83] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_86 
+ bl[84] br[84] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_87 
+ bl[85] br[85] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_88 
+ bl[86] br[86] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_89 
+ bl[87] br[87] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_90 
+ bl[88] br[88] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_91 
+ bl[89] br[89] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_92 
+ bl[90] br[90] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_93 
+ bl[91] br[91] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_94 
+ bl[92] br[92] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_95 
+ bl[93] br[93] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_96 
+ bl[94] br[94] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_97 
+ bl[95] br[95] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_98 
+ bl[96] br[96] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_99 
+ bl[97] br[97] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_100 
+ bl[98] br[98] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_101 
+ bl[99] br[99] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_102 
+ bl[100] br[100] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_103 
+ bl[101] br[101] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_104 
+ bl[102] br[102] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_105 
+ bl[103] br[103] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_106 
+ bl[104] br[104] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_107 
+ bl[105] br[105] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_108 
+ bl[106] br[106] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_109 
+ bl[107] br[107] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_110 
+ bl[108] br[108] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_111 
+ bl[109] br[109] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_112 
+ bl[110] br[110] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_113 
+ bl[111] br[111] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_114 
+ bl[112] br[112] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_115 
+ bl[113] br[113] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_116 
+ bl[114] br[114] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_117 
+ bl[115] br[115] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_118 
+ bl[116] br[116] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_119 
+ bl[117] br[117] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_120 
+ bl[118] br[118] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_121 
+ bl[119] br[119] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_122 
+ bl[120] br[120] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_123 
+ bl[121] br[121] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_124 
+ bl[122] br[122] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_125 
+ bl[123] br[123] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_126 
+ bl[124] br[124] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_127 
+ bl[125] br[125] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_128 
+ bl[126] br[126] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_129 
+ bl[127] br[127] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_130 
+ bl[128] br[128] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_131 
+ bl[129] br[129] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_132 
+ bl[130] br[130] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_133 
+ bl[131] br[131] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_134 
+ bl[132] br[132] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_135 
+ bl[133] br[133] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_136 
+ bl[134] br[134] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_137 
+ bl[135] br[135] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_138 
+ bl[136] br[136] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_139 
+ bl[137] br[137] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_140 
+ bl[138] br[138] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_141 
+ bl[139] br[139] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_142 
+ bl[140] br[140] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_143 
+ bl[141] br[141] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_144 
+ bl[142] br[142] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_145 
+ bl[143] br[143] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_146 
+ bl[144] br[144] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_147 
+ bl[145] br[145] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_148 
+ bl[146] br[146] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_149 
+ bl[147] br[147] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_150 
+ bl[148] br[148] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_151 
+ bl[149] br[149] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_152 
+ bl[150] br[150] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_153 
+ bl[151] br[151] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_154 
+ bl[152] br[152] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_155 
+ bl[153] br[153] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_156 
+ bl[154] br[154] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_157 
+ bl[155] br[155] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_158 
+ bl[156] br[156] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_159 
+ bl[157] br[157] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_160 
+ bl[158] br[158] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_161 
+ bl[159] br[159] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_162 
+ bl[160] br[160] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_163 
+ bl[161] br[161] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_164 
+ bl[162] br[162] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_165 
+ bl[163] br[163] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_166 
+ bl[164] br[164] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_167 
+ bl[165] br[165] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_168 
+ bl[166] br[166] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_169 
+ bl[167] br[167] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_170 
+ bl[168] br[168] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_171 
+ bl[169] br[169] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_172 
+ bl[170] br[170] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_173 
+ bl[171] br[171] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_174 
+ bl[172] br[172] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_175 
+ bl[173] br[173] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_176 
+ bl[174] br[174] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_177 
+ bl[175] br[175] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_178 
+ bl[176] br[176] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_179 
+ bl[177] br[177] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_180 
+ bl[178] br[178] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_181 
+ bl[179] br[179] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_182 
+ bl[180] br[180] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_183 
+ bl[181] br[181] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_184 
+ bl[182] br[182] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_185 
+ bl[183] br[183] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_186 
+ bl[184] br[184] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_187 
+ bl[185] br[185] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_188 
+ bl[186] br[186] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_189 
+ bl[187] br[187] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_190 
+ bl[188] br[188] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_191 
+ bl[189] br[189] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_192 
+ bl[190] br[190] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_193 
+ bl[191] br[191] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_194 
+ bl[192] br[192] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_195 
+ bl[193] br[193] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_196 
+ bl[194] br[194] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_197 
+ bl[195] br[195] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_198 
+ bl[196] br[196] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_199 
+ bl[197] br[197] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_200 
+ bl[198] br[198] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_201 
+ bl[199] br[199] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_202 
+ bl[200] br[200] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_203 
+ bl[201] br[201] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_204 
+ bl[202] br[202] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_205 
+ bl[203] br[203] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_206 
+ bl[204] br[204] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_207 
+ bl[205] br[205] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_208 
+ bl[206] br[206] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_209 
+ bl[207] br[207] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_210 
+ bl[208] br[208] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_211 
+ bl[209] br[209] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_212 
+ bl[210] br[210] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_213 
+ bl[211] br[211] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_214 
+ bl[212] br[212] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_215 
+ bl[213] br[213] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_216 
+ bl[214] br[214] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_217 
+ bl[215] br[215] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_218 
+ bl[216] br[216] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_219 
+ bl[217] br[217] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_220 
+ bl[218] br[218] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_221 
+ bl[219] br[219] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_222 
+ bl[220] br[220] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_223 
+ bl[221] br[221] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_224 
+ bl[222] br[222] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_225 
+ bl[223] br[223] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_226 
+ bl[224] br[224] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_227 
+ bl[225] br[225] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_228 
+ bl[226] br[226] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_229 
+ bl[227] br[227] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_230 
+ bl[228] br[228] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_231 
+ bl[229] br[229] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_232 
+ bl[230] br[230] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_233 
+ bl[231] br[231] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_234 
+ bl[232] br[232] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_235 
+ bl[233] br[233] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_236 
+ bl[234] br[234] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_237 
+ bl[235] br[235] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_238 
+ bl[236] br[236] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_239 
+ bl[237] br[237] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_240 
+ bl[238] br[238] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_241 
+ bl[239] br[239] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_242 
+ bl[240] br[240] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_243 
+ bl[241] br[241] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_244 
+ bl[242] br[242] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_245 
+ bl[243] br[243] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_246 
+ bl[244] br[244] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_247 
+ bl[245] br[245] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_248 
+ bl[246] br[246] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_249 
+ bl[247] br[247] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_250 
+ bl[248] br[248] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_251 
+ bl[249] br[249] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_252 
+ bl[250] br[250] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_253 
+ bl[251] br[251] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_254 
+ bl[252] br[252] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_255 
+ bl[253] br[253] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_256 
+ bl[254] br[254] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_257 
+ bl[255] br[255] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_258 
+ vdd vdd vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_259 
+ vdd vdd vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_0 
+ vdd vdd vss vdd vpb vnb wl[117] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_119_1 
+ rbl rbr vss vdd vpb vnb wl[117] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_119_2 
+ bl[0] br[0] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_3 
+ bl[1] br[1] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_4 
+ bl[2] br[2] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_5 
+ bl[3] br[3] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_6 
+ bl[4] br[4] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_7 
+ bl[5] br[5] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_8 
+ bl[6] br[6] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_9 
+ bl[7] br[7] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_10 
+ bl[8] br[8] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_11 
+ bl[9] br[9] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_12 
+ bl[10] br[10] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_13 
+ bl[11] br[11] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_14 
+ bl[12] br[12] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_15 
+ bl[13] br[13] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_16 
+ bl[14] br[14] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_17 
+ bl[15] br[15] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_18 
+ bl[16] br[16] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_19 
+ bl[17] br[17] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_20 
+ bl[18] br[18] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_21 
+ bl[19] br[19] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_22 
+ bl[20] br[20] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_23 
+ bl[21] br[21] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_24 
+ bl[22] br[22] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_25 
+ bl[23] br[23] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_26 
+ bl[24] br[24] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_27 
+ bl[25] br[25] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_28 
+ bl[26] br[26] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_29 
+ bl[27] br[27] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_30 
+ bl[28] br[28] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_31 
+ bl[29] br[29] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_32 
+ bl[30] br[30] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_33 
+ bl[31] br[31] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_34 
+ bl[32] br[32] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_35 
+ bl[33] br[33] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_36 
+ bl[34] br[34] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_37 
+ bl[35] br[35] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_38 
+ bl[36] br[36] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_39 
+ bl[37] br[37] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_40 
+ bl[38] br[38] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_41 
+ bl[39] br[39] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_42 
+ bl[40] br[40] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_43 
+ bl[41] br[41] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_44 
+ bl[42] br[42] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_45 
+ bl[43] br[43] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_46 
+ bl[44] br[44] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_47 
+ bl[45] br[45] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_48 
+ bl[46] br[46] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_49 
+ bl[47] br[47] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_50 
+ bl[48] br[48] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_51 
+ bl[49] br[49] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_52 
+ bl[50] br[50] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_53 
+ bl[51] br[51] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_54 
+ bl[52] br[52] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_55 
+ bl[53] br[53] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_56 
+ bl[54] br[54] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_57 
+ bl[55] br[55] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_58 
+ bl[56] br[56] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_59 
+ bl[57] br[57] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_60 
+ bl[58] br[58] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_61 
+ bl[59] br[59] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_62 
+ bl[60] br[60] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_63 
+ bl[61] br[61] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_64 
+ bl[62] br[62] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_65 
+ bl[63] br[63] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_66 
+ bl[64] br[64] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_67 
+ bl[65] br[65] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_68 
+ bl[66] br[66] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_69 
+ bl[67] br[67] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_70 
+ bl[68] br[68] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_71 
+ bl[69] br[69] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_72 
+ bl[70] br[70] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_73 
+ bl[71] br[71] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_74 
+ bl[72] br[72] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_75 
+ bl[73] br[73] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_76 
+ bl[74] br[74] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_77 
+ bl[75] br[75] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_78 
+ bl[76] br[76] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_79 
+ bl[77] br[77] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_80 
+ bl[78] br[78] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_81 
+ bl[79] br[79] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_82 
+ bl[80] br[80] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_83 
+ bl[81] br[81] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_84 
+ bl[82] br[82] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_85 
+ bl[83] br[83] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_86 
+ bl[84] br[84] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_87 
+ bl[85] br[85] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_88 
+ bl[86] br[86] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_89 
+ bl[87] br[87] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_90 
+ bl[88] br[88] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_91 
+ bl[89] br[89] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_92 
+ bl[90] br[90] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_93 
+ bl[91] br[91] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_94 
+ bl[92] br[92] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_95 
+ bl[93] br[93] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_96 
+ bl[94] br[94] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_97 
+ bl[95] br[95] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_98 
+ bl[96] br[96] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_99 
+ bl[97] br[97] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_100 
+ bl[98] br[98] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_101 
+ bl[99] br[99] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_102 
+ bl[100] br[100] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_103 
+ bl[101] br[101] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_104 
+ bl[102] br[102] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_105 
+ bl[103] br[103] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_106 
+ bl[104] br[104] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_107 
+ bl[105] br[105] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_108 
+ bl[106] br[106] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_109 
+ bl[107] br[107] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_110 
+ bl[108] br[108] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_111 
+ bl[109] br[109] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_112 
+ bl[110] br[110] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_113 
+ bl[111] br[111] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_114 
+ bl[112] br[112] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_115 
+ bl[113] br[113] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_116 
+ bl[114] br[114] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_117 
+ bl[115] br[115] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_118 
+ bl[116] br[116] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_119 
+ bl[117] br[117] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_120 
+ bl[118] br[118] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_121 
+ bl[119] br[119] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_122 
+ bl[120] br[120] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_123 
+ bl[121] br[121] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_124 
+ bl[122] br[122] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_125 
+ bl[123] br[123] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_126 
+ bl[124] br[124] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_127 
+ bl[125] br[125] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_128 
+ bl[126] br[126] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_129 
+ bl[127] br[127] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_130 
+ bl[128] br[128] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_131 
+ bl[129] br[129] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_132 
+ bl[130] br[130] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_133 
+ bl[131] br[131] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_134 
+ bl[132] br[132] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_135 
+ bl[133] br[133] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_136 
+ bl[134] br[134] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_137 
+ bl[135] br[135] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_138 
+ bl[136] br[136] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_139 
+ bl[137] br[137] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_140 
+ bl[138] br[138] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_141 
+ bl[139] br[139] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_142 
+ bl[140] br[140] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_143 
+ bl[141] br[141] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_144 
+ bl[142] br[142] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_145 
+ bl[143] br[143] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_146 
+ bl[144] br[144] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_147 
+ bl[145] br[145] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_148 
+ bl[146] br[146] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_149 
+ bl[147] br[147] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_150 
+ bl[148] br[148] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_151 
+ bl[149] br[149] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_152 
+ bl[150] br[150] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_153 
+ bl[151] br[151] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_154 
+ bl[152] br[152] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_155 
+ bl[153] br[153] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_156 
+ bl[154] br[154] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_157 
+ bl[155] br[155] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_158 
+ bl[156] br[156] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_159 
+ bl[157] br[157] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_160 
+ bl[158] br[158] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_161 
+ bl[159] br[159] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_162 
+ bl[160] br[160] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_163 
+ bl[161] br[161] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_164 
+ bl[162] br[162] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_165 
+ bl[163] br[163] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_166 
+ bl[164] br[164] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_167 
+ bl[165] br[165] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_168 
+ bl[166] br[166] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_169 
+ bl[167] br[167] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_170 
+ bl[168] br[168] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_171 
+ bl[169] br[169] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_172 
+ bl[170] br[170] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_173 
+ bl[171] br[171] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_174 
+ bl[172] br[172] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_175 
+ bl[173] br[173] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_176 
+ bl[174] br[174] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_177 
+ bl[175] br[175] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_178 
+ bl[176] br[176] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_179 
+ bl[177] br[177] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_180 
+ bl[178] br[178] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_181 
+ bl[179] br[179] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_182 
+ bl[180] br[180] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_183 
+ bl[181] br[181] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_184 
+ bl[182] br[182] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_185 
+ bl[183] br[183] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_186 
+ bl[184] br[184] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_187 
+ bl[185] br[185] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_188 
+ bl[186] br[186] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_189 
+ bl[187] br[187] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_190 
+ bl[188] br[188] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_191 
+ bl[189] br[189] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_192 
+ bl[190] br[190] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_193 
+ bl[191] br[191] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_194 
+ bl[192] br[192] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_195 
+ bl[193] br[193] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_196 
+ bl[194] br[194] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_197 
+ bl[195] br[195] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_198 
+ bl[196] br[196] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_199 
+ bl[197] br[197] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_200 
+ bl[198] br[198] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_201 
+ bl[199] br[199] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_202 
+ bl[200] br[200] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_203 
+ bl[201] br[201] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_204 
+ bl[202] br[202] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_205 
+ bl[203] br[203] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_206 
+ bl[204] br[204] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_207 
+ bl[205] br[205] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_208 
+ bl[206] br[206] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_209 
+ bl[207] br[207] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_210 
+ bl[208] br[208] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_211 
+ bl[209] br[209] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_212 
+ bl[210] br[210] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_213 
+ bl[211] br[211] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_214 
+ bl[212] br[212] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_215 
+ bl[213] br[213] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_216 
+ bl[214] br[214] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_217 
+ bl[215] br[215] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_218 
+ bl[216] br[216] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_219 
+ bl[217] br[217] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_220 
+ bl[218] br[218] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_221 
+ bl[219] br[219] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_222 
+ bl[220] br[220] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_223 
+ bl[221] br[221] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_224 
+ bl[222] br[222] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_225 
+ bl[223] br[223] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_226 
+ bl[224] br[224] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_227 
+ bl[225] br[225] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_228 
+ bl[226] br[226] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_229 
+ bl[227] br[227] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_230 
+ bl[228] br[228] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_231 
+ bl[229] br[229] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_232 
+ bl[230] br[230] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_233 
+ bl[231] br[231] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_234 
+ bl[232] br[232] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_235 
+ bl[233] br[233] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_236 
+ bl[234] br[234] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_237 
+ bl[235] br[235] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_238 
+ bl[236] br[236] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_239 
+ bl[237] br[237] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_240 
+ bl[238] br[238] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_241 
+ bl[239] br[239] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_242 
+ bl[240] br[240] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_243 
+ bl[241] br[241] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_244 
+ bl[242] br[242] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_245 
+ bl[243] br[243] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_246 
+ bl[244] br[244] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_247 
+ bl[245] br[245] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_248 
+ bl[246] br[246] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_249 
+ bl[247] br[247] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_250 
+ bl[248] br[248] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_251 
+ bl[249] br[249] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_252 
+ bl[250] br[250] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_253 
+ bl[251] br[251] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_254 
+ bl[252] br[252] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_255 
+ bl[253] br[253] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_256 
+ bl[254] br[254] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_257 
+ bl[255] br[255] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_258 
+ vdd vdd vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_259 
+ vdd vdd vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_0 
+ vdd vdd vss vdd vpb vnb wl[118] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_120_1 
+ rbl rbr vss vdd vpb vnb wl[118] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_120_2 
+ bl[0] br[0] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_3 
+ bl[1] br[1] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_4 
+ bl[2] br[2] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_5 
+ bl[3] br[3] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_6 
+ bl[4] br[4] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_7 
+ bl[5] br[5] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_8 
+ bl[6] br[6] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_9 
+ bl[7] br[7] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_10 
+ bl[8] br[8] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_11 
+ bl[9] br[9] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_12 
+ bl[10] br[10] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_13 
+ bl[11] br[11] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_14 
+ bl[12] br[12] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_15 
+ bl[13] br[13] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_16 
+ bl[14] br[14] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_17 
+ bl[15] br[15] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_18 
+ bl[16] br[16] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_19 
+ bl[17] br[17] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_20 
+ bl[18] br[18] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_21 
+ bl[19] br[19] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_22 
+ bl[20] br[20] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_23 
+ bl[21] br[21] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_24 
+ bl[22] br[22] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_25 
+ bl[23] br[23] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_26 
+ bl[24] br[24] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_27 
+ bl[25] br[25] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_28 
+ bl[26] br[26] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_29 
+ bl[27] br[27] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_30 
+ bl[28] br[28] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_31 
+ bl[29] br[29] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_32 
+ bl[30] br[30] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_33 
+ bl[31] br[31] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_34 
+ bl[32] br[32] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_35 
+ bl[33] br[33] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_36 
+ bl[34] br[34] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_37 
+ bl[35] br[35] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_38 
+ bl[36] br[36] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_39 
+ bl[37] br[37] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_40 
+ bl[38] br[38] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_41 
+ bl[39] br[39] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_42 
+ bl[40] br[40] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_43 
+ bl[41] br[41] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_44 
+ bl[42] br[42] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_45 
+ bl[43] br[43] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_46 
+ bl[44] br[44] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_47 
+ bl[45] br[45] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_48 
+ bl[46] br[46] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_49 
+ bl[47] br[47] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_50 
+ bl[48] br[48] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_51 
+ bl[49] br[49] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_52 
+ bl[50] br[50] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_53 
+ bl[51] br[51] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_54 
+ bl[52] br[52] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_55 
+ bl[53] br[53] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_56 
+ bl[54] br[54] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_57 
+ bl[55] br[55] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_58 
+ bl[56] br[56] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_59 
+ bl[57] br[57] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_60 
+ bl[58] br[58] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_61 
+ bl[59] br[59] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_62 
+ bl[60] br[60] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_63 
+ bl[61] br[61] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_64 
+ bl[62] br[62] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_65 
+ bl[63] br[63] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_66 
+ bl[64] br[64] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_67 
+ bl[65] br[65] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_68 
+ bl[66] br[66] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_69 
+ bl[67] br[67] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_70 
+ bl[68] br[68] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_71 
+ bl[69] br[69] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_72 
+ bl[70] br[70] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_73 
+ bl[71] br[71] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_74 
+ bl[72] br[72] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_75 
+ bl[73] br[73] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_76 
+ bl[74] br[74] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_77 
+ bl[75] br[75] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_78 
+ bl[76] br[76] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_79 
+ bl[77] br[77] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_80 
+ bl[78] br[78] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_81 
+ bl[79] br[79] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_82 
+ bl[80] br[80] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_83 
+ bl[81] br[81] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_84 
+ bl[82] br[82] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_85 
+ bl[83] br[83] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_86 
+ bl[84] br[84] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_87 
+ bl[85] br[85] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_88 
+ bl[86] br[86] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_89 
+ bl[87] br[87] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_90 
+ bl[88] br[88] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_91 
+ bl[89] br[89] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_92 
+ bl[90] br[90] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_93 
+ bl[91] br[91] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_94 
+ bl[92] br[92] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_95 
+ bl[93] br[93] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_96 
+ bl[94] br[94] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_97 
+ bl[95] br[95] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_98 
+ bl[96] br[96] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_99 
+ bl[97] br[97] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_100 
+ bl[98] br[98] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_101 
+ bl[99] br[99] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_102 
+ bl[100] br[100] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_103 
+ bl[101] br[101] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_104 
+ bl[102] br[102] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_105 
+ bl[103] br[103] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_106 
+ bl[104] br[104] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_107 
+ bl[105] br[105] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_108 
+ bl[106] br[106] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_109 
+ bl[107] br[107] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_110 
+ bl[108] br[108] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_111 
+ bl[109] br[109] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_112 
+ bl[110] br[110] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_113 
+ bl[111] br[111] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_114 
+ bl[112] br[112] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_115 
+ bl[113] br[113] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_116 
+ bl[114] br[114] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_117 
+ bl[115] br[115] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_118 
+ bl[116] br[116] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_119 
+ bl[117] br[117] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_120 
+ bl[118] br[118] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_121 
+ bl[119] br[119] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_122 
+ bl[120] br[120] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_123 
+ bl[121] br[121] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_124 
+ bl[122] br[122] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_125 
+ bl[123] br[123] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_126 
+ bl[124] br[124] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_127 
+ bl[125] br[125] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_128 
+ bl[126] br[126] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_129 
+ bl[127] br[127] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_130 
+ bl[128] br[128] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_131 
+ bl[129] br[129] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_132 
+ bl[130] br[130] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_133 
+ bl[131] br[131] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_134 
+ bl[132] br[132] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_135 
+ bl[133] br[133] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_136 
+ bl[134] br[134] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_137 
+ bl[135] br[135] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_138 
+ bl[136] br[136] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_139 
+ bl[137] br[137] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_140 
+ bl[138] br[138] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_141 
+ bl[139] br[139] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_142 
+ bl[140] br[140] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_143 
+ bl[141] br[141] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_144 
+ bl[142] br[142] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_145 
+ bl[143] br[143] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_146 
+ bl[144] br[144] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_147 
+ bl[145] br[145] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_148 
+ bl[146] br[146] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_149 
+ bl[147] br[147] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_150 
+ bl[148] br[148] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_151 
+ bl[149] br[149] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_152 
+ bl[150] br[150] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_153 
+ bl[151] br[151] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_154 
+ bl[152] br[152] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_155 
+ bl[153] br[153] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_156 
+ bl[154] br[154] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_157 
+ bl[155] br[155] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_158 
+ bl[156] br[156] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_159 
+ bl[157] br[157] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_160 
+ bl[158] br[158] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_161 
+ bl[159] br[159] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_162 
+ bl[160] br[160] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_163 
+ bl[161] br[161] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_164 
+ bl[162] br[162] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_165 
+ bl[163] br[163] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_166 
+ bl[164] br[164] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_167 
+ bl[165] br[165] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_168 
+ bl[166] br[166] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_169 
+ bl[167] br[167] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_170 
+ bl[168] br[168] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_171 
+ bl[169] br[169] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_172 
+ bl[170] br[170] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_173 
+ bl[171] br[171] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_174 
+ bl[172] br[172] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_175 
+ bl[173] br[173] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_176 
+ bl[174] br[174] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_177 
+ bl[175] br[175] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_178 
+ bl[176] br[176] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_179 
+ bl[177] br[177] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_180 
+ bl[178] br[178] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_181 
+ bl[179] br[179] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_182 
+ bl[180] br[180] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_183 
+ bl[181] br[181] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_184 
+ bl[182] br[182] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_185 
+ bl[183] br[183] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_186 
+ bl[184] br[184] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_187 
+ bl[185] br[185] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_188 
+ bl[186] br[186] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_189 
+ bl[187] br[187] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_190 
+ bl[188] br[188] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_191 
+ bl[189] br[189] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_192 
+ bl[190] br[190] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_193 
+ bl[191] br[191] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_194 
+ bl[192] br[192] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_195 
+ bl[193] br[193] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_196 
+ bl[194] br[194] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_197 
+ bl[195] br[195] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_198 
+ bl[196] br[196] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_199 
+ bl[197] br[197] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_200 
+ bl[198] br[198] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_201 
+ bl[199] br[199] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_202 
+ bl[200] br[200] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_203 
+ bl[201] br[201] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_204 
+ bl[202] br[202] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_205 
+ bl[203] br[203] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_206 
+ bl[204] br[204] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_207 
+ bl[205] br[205] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_208 
+ bl[206] br[206] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_209 
+ bl[207] br[207] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_210 
+ bl[208] br[208] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_211 
+ bl[209] br[209] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_212 
+ bl[210] br[210] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_213 
+ bl[211] br[211] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_214 
+ bl[212] br[212] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_215 
+ bl[213] br[213] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_216 
+ bl[214] br[214] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_217 
+ bl[215] br[215] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_218 
+ bl[216] br[216] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_219 
+ bl[217] br[217] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_220 
+ bl[218] br[218] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_221 
+ bl[219] br[219] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_222 
+ bl[220] br[220] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_223 
+ bl[221] br[221] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_224 
+ bl[222] br[222] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_225 
+ bl[223] br[223] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_226 
+ bl[224] br[224] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_227 
+ bl[225] br[225] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_228 
+ bl[226] br[226] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_229 
+ bl[227] br[227] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_230 
+ bl[228] br[228] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_231 
+ bl[229] br[229] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_232 
+ bl[230] br[230] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_233 
+ bl[231] br[231] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_234 
+ bl[232] br[232] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_235 
+ bl[233] br[233] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_236 
+ bl[234] br[234] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_237 
+ bl[235] br[235] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_238 
+ bl[236] br[236] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_239 
+ bl[237] br[237] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_240 
+ bl[238] br[238] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_241 
+ bl[239] br[239] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_242 
+ bl[240] br[240] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_243 
+ bl[241] br[241] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_244 
+ bl[242] br[242] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_245 
+ bl[243] br[243] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_246 
+ bl[244] br[244] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_247 
+ bl[245] br[245] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_248 
+ bl[246] br[246] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_249 
+ bl[247] br[247] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_250 
+ bl[248] br[248] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_251 
+ bl[249] br[249] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_252 
+ bl[250] br[250] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_253 
+ bl[251] br[251] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_254 
+ bl[252] br[252] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_255 
+ bl[253] br[253] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_256 
+ bl[254] br[254] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_257 
+ bl[255] br[255] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_258 
+ vdd vdd vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_259 
+ vdd vdd vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_0 
+ vdd vdd vss vdd vpb vnb wl[119] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_121_1 
+ rbl rbr vss vdd vpb vnb wl[119] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_121_2 
+ bl[0] br[0] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_3 
+ bl[1] br[1] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_4 
+ bl[2] br[2] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_5 
+ bl[3] br[3] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_6 
+ bl[4] br[4] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_7 
+ bl[5] br[5] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_8 
+ bl[6] br[6] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_9 
+ bl[7] br[7] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_10 
+ bl[8] br[8] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_11 
+ bl[9] br[9] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_12 
+ bl[10] br[10] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_13 
+ bl[11] br[11] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_14 
+ bl[12] br[12] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_15 
+ bl[13] br[13] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_16 
+ bl[14] br[14] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_17 
+ bl[15] br[15] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_18 
+ bl[16] br[16] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_19 
+ bl[17] br[17] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_20 
+ bl[18] br[18] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_21 
+ bl[19] br[19] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_22 
+ bl[20] br[20] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_23 
+ bl[21] br[21] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_24 
+ bl[22] br[22] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_25 
+ bl[23] br[23] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_26 
+ bl[24] br[24] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_27 
+ bl[25] br[25] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_28 
+ bl[26] br[26] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_29 
+ bl[27] br[27] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_30 
+ bl[28] br[28] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_31 
+ bl[29] br[29] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_32 
+ bl[30] br[30] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_33 
+ bl[31] br[31] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_34 
+ bl[32] br[32] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_35 
+ bl[33] br[33] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_36 
+ bl[34] br[34] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_37 
+ bl[35] br[35] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_38 
+ bl[36] br[36] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_39 
+ bl[37] br[37] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_40 
+ bl[38] br[38] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_41 
+ bl[39] br[39] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_42 
+ bl[40] br[40] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_43 
+ bl[41] br[41] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_44 
+ bl[42] br[42] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_45 
+ bl[43] br[43] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_46 
+ bl[44] br[44] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_47 
+ bl[45] br[45] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_48 
+ bl[46] br[46] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_49 
+ bl[47] br[47] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_50 
+ bl[48] br[48] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_51 
+ bl[49] br[49] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_52 
+ bl[50] br[50] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_53 
+ bl[51] br[51] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_54 
+ bl[52] br[52] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_55 
+ bl[53] br[53] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_56 
+ bl[54] br[54] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_57 
+ bl[55] br[55] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_58 
+ bl[56] br[56] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_59 
+ bl[57] br[57] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_60 
+ bl[58] br[58] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_61 
+ bl[59] br[59] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_62 
+ bl[60] br[60] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_63 
+ bl[61] br[61] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_64 
+ bl[62] br[62] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_65 
+ bl[63] br[63] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_66 
+ bl[64] br[64] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_67 
+ bl[65] br[65] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_68 
+ bl[66] br[66] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_69 
+ bl[67] br[67] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_70 
+ bl[68] br[68] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_71 
+ bl[69] br[69] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_72 
+ bl[70] br[70] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_73 
+ bl[71] br[71] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_74 
+ bl[72] br[72] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_75 
+ bl[73] br[73] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_76 
+ bl[74] br[74] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_77 
+ bl[75] br[75] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_78 
+ bl[76] br[76] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_79 
+ bl[77] br[77] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_80 
+ bl[78] br[78] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_81 
+ bl[79] br[79] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_82 
+ bl[80] br[80] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_83 
+ bl[81] br[81] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_84 
+ bl[82] br[82] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_85 
+ bl[83] br[83] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_86 
+ bl[84] br[84] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_87 
+ bl[85] br[85] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_88 
+ bl[86] br[86] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_89 
+ bl[87] br[87] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_90 
+ bl[88] br[88] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_91 
+ bl[89] br[89] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_92 
+ bl[90] br[90] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_93 
+ bl[91] br[91] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_94 
+ bl[92] br[92] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_95 
+ bl[93] br[93] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_96 
+ bl[94] br[94] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_97 
+ bl[95] br[95] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_98 
+ bl[96] br[96] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_99 
+ bl[97] br[97] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_100 
+ bl[98] br[98] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_101 
+ bl[99] br[99] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_102 
+ bl[100] br[100] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_103 
+ bl[101] br[101] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_104 
+ bl[102] br[102] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_105 
+ bl[103] br[103] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_106 
+ bl[104] br[104] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_107 
+ bl[105] br[105] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_108 
+ bl[106] br[106] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_109 
+ bl[107] br[107] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_110 
+ bl[108] br[108] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_111 
+ bl[109] br[109] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_112 
+ bl[110] br[110] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_113 
+ bl[111] br[111] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_114 
+ bl[112] br[112] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_115 
+ bl[113] br[113] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_116 
+ bl[114] br[114] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_117 
+ bl[115] br[115] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_118 
+ bl[116] br[116] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_119 
+ bl[117] br[117] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_120 
+ bl[118] br[118] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_121 
+ bl[119] br[119] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_122 
+ bl[120] br[120] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_123 
+ bl[121] br[121] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_124 
+ bl[122] br[122] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_125 
+ bl[123] br[123] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_126 
+ bl[124] br[124] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_127 
+ bl[125] br[125] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_128 
+ bl[126] br[126] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_129 
+ bl[127] br[127] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_130 
+ bl[128] br[128] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_131 
+ bl[129] br[129] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_132 
+ bl[130] br[130] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_133 
+ bl[131] br[131] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_134 
+ bl[132] br[132] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_135 
+ bl[133] br[133] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_136 
+ bl[134] br[134] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_137 
+ bl[135] br[135] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_138 
+ bl[136] br[136] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_139 
+ bl[137] br[137] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_140 
+ bl[138] br[138] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_141 
+ bl[139] br[139] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_142 
+ bl[140] br[140] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_143 
+ bl[141] br[141] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_144 
+ bl[142] br[142] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_145 
+ bl[143] br[143] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_146 
+ bl[144] br[144] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_147 
+ bl[145] br[145] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_148 
+ bl[146] br[146] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_149 
+ bl[147] br[147] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_150 
+ bl[148] br[148] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_151 
+ bl[149] br[149] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_152 
+ bl[150] br[150] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_153 
+ bl[151] br[151] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_154 
+ bl[152] br[152] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_155 
+ bl[153] br[153] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_156 
+ bl[154] br[154] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_157 
+ bl[155] br[155] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_158 
+ bl[156] br[156] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_159 
+ bl[157] br[157] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_160 
+ bl[158] br[158] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_161 
+ bl[159] br[159] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_162 
+ bl[160] br[160] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_163 
+ bl[161] br[161] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_164 
+ bl[162] br[162] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_165 
+ bl[163] br[163] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_166 
+ bl[164] br[164] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_167 
+ bl[165] br[165] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_168 
+ bl[166] br[166] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_169 
+ bl[167] br[167] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_170 
+ bl[168] br[168] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_171 
+ bl[169] br[169] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_172 
+ bl[170] br[170] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_173 
+ bl[171] br[171] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_174 
+ bl[172] br[172] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_175 
+ bl[173] br[173] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_176 
+ bl[174] br[174] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_177 
+ bl[175] br[175] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_178 
+ bl[176] br[176] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_179 
+ bl[177] br[177] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_180 
+ bl[178] br[178] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_181 
+ bl[179] br[179] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_182 
+ bl[180] br[180] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_183 
+ bl[181] br[181] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_184 
+ bl[182] br[182] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_185 
+ bl[183] br[183] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_186 
+ bl[184] br[184] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_187 
+ bl[185] br[185] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_188 
+ bl[186] br[186] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_189 
+ bl[187] br[187] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_190 
+ bl[188] br[188] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_191 
+ bl[189] br[189] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_192 
+ bl[190] br[190] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_193 
+ bl[191] br[191] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_194 
+ bl[192] br[192] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_195 
+ bl[193] br[193] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_196 
+ bl[194] br[194] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_197 
+ bl[195] br[195] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_198 
+ bl[196] br[196] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_199 
+ bl[197] br[197] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_200 
+ bl[198] br[198] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_201 
+ bl[199] br[199] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_202 
+ bl[200] br[200] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_203 
+ bl[201] br[201] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_204 
+ bl[202] br[202] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_205 
+ bl[203] br[203] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_206 
+ bl[204] br[204] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_207 
+ bl[205] br[205] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_208 
+ bl[206] br[206] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_209 
+ bl[207] br[207] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_210 
+ bl[208] br[208] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_211 
+ bl[209] br[209] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_212 
+ bl[210] br[210] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_213 
+ bl[211] br[211] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_214 
+ bl[212] br[212] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_215 
+ bl[213] br[213] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_216 
+ bl[214] br[214] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_217 
+ bl[215] br[215] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_218 
+ bl[216] br[216] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_219 
+ bl[217] br[217] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_220 
+ bl[218] br[218] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_221 
+ bl[219] br[219] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_222 
+ bl[220] br[220] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_223 
+ bl[221] br[221] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_224 
+ bl[222] br[222] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_225 
+ bl[223] br[223] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_226 
+ bl[224] br[224] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_227 
+ bl[225] br[225] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_228 
+ bl[226] br[226] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_229 
+ bl[227] br[227] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_230 
+ bl[228] br[228] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_231 
+ bl[229] br[229] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_232 
+ bl[230] br[230] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_233 
+ bl[231] br[231] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_234 
+ bl[232] br[232] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_235 
+ bl[233] br[233] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_236 
+ bl[234] br[234] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_237 
+ bl[235] br[235] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_238 
+ bl[236] br[236] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_239 
+ bl[237] br[237] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_240 
+ bl[238] br[238] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_241 
+ bl[239] br[239] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_242 
+ bl[240] br[240] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_243 
+ bl[241] br[241] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_244 
+ bl[242] br[242] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_245 
+ bl[243] br[243] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_246 
+ bl[244] br[244] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_247 
+ bl[245] br[245] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_248 
+ bl[246] br[246] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_249 
+ bl[247] br[247] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_250 
+ bl[248] br[248] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_251 
+ bl[249] br[249] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_252 
+ bl[250] br[250] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_253 
+ bl[251] br[251] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_254 
+ bl[252] br[252] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_255 
+ bl[253] br[253] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_256 
+ bl[254] br[254] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_257 
+ bl[255] br[255] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_258 
+ vdd vdd vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_259 
+ vdd vdd vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_0 
+ vdd vdd vss vdd vpb vnb wl[120] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_122_1 
+ rbl rbr vss vdd vpb vnb wl[120] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_122_2 
+ bl[0] br[0] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_3 
+ bl[1] br[1] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_4 
+ bl[2] br[2] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_5 
+ bl[3] br[3] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_6 
+ bl[4] br[4] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_7 
+ bl[5] br[5] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_8 
+ bl[6] br[6] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_9 
+ bl[7] br[7] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_10 
+ bl[8] br[8] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_11 
+ bl[9] br[9] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_12 
+ bl[10] br[10] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_13 
+ bl[11] br[11] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_14 
+ bl[12] br[12] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_15 
+ bl[13] br[13] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_16 
+ bl[14] br[14] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_17 
+ bl[15] br[15] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_18 
+ bl[16] br[16] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_19 
+ bl[17] br[17] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_20 
+ bl[18] br[18] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_21 
+ bl[19] br[19] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_22 
+ bl[20] br[20] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_23 
+ bl[21] br[21] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_24 
+ bl[22] br[22] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_25 
+ bl[23] br[23] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_26 
+ bl[24] br[24] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_27 
+ bl[25] br[25] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_28 
+ bl[26] br[26] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_29 
+ bl[27] br[27] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_30 
+ bl[28] br[28] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_31 
+ bl[29] br[29] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_32 
+ bl[30] br[30] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_33 
+ bl[31] br[31] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_34 
+ bl[32] br[32] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_35 
+ bl[33] br[33] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_36 
+ bl[34] br[34] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_37 
+ bl[35] br[35] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_38 
+ bl[36] br[36] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_39 
+ bl[37] br[37] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_40 
+ bl[38] br[38] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_41 
+ bl[39] br[39] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_42 
+ bl[40] br[40] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_43 
+ bl[41] br[41] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_44 
+ bl[42] br[42] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_45 
+ bl[43] br[43] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_46 
+ bl[44] br[44] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_47 
+ bl[45] br[45] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_48 
+ bl[46] br[46] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_49 
+ bl[47] br[47] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_50 
+ bl[48] br[48] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_51 
+ bl[49] br[49] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_52 
+ bl[50] br[50] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_53 
+ bl[51] br[51] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_54 
+ bl[52] br[52] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_55 
+ bl[53] br[53] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_56 
+ bl[54] br[54] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_57 
+ bl[55] br[55] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_58 
+ bl[56] br[56] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_59 
+ bl[57] br[57] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_60 
+ bl[58] br[58] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_61 
+ bl[59] br[59] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_62 
+ bl[60] br[60] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_63 
+ bl[61] br[61] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_64 
+ bl[62] br[62] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_65 
+ bl[63] br[63] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_66 
+ bl[64] br[64] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_67 
+ bl[65] br[65] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_68 
+ bl[66] br[66] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_69 
+ bl[67] br[67] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_70 
+ bl[68] br[68] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_71 
+ bl[69] br[69] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_72 
+ bl[70] br[70] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_73 
+ bl[71] br[71] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_74 
+ bl[72] br[72] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_75 
+ bl[73] br[73] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_76 
+ bl[74] br[74] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_77 
+ bl[75] br[75] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_78 
+ bl[76] br[76] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_79 
+ bl[77] br[77] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_80 
+ bl[78] br[78] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_81 
+ bl[79] br[79] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_82 
+ bl[80] br[80] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_83 
+ bl[81] br[81] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_84 
+ bl[82] br[82] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_85 
+ bl[83] br[83] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_86 
+ bl[84] br[84] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_87 
+ bl[85] br[85] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_88 
+ bl[86] br[86] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_89 
+ bl[87] br[87] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_90 
+ bl[88] br[88] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_91 
+ bl[89] br[89] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_92 
+ bl[90] br[90] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_93 
+ bl[91] br[91] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_94 
+ bl[92] br[92] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_95 
+ bl[93] br[93] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_96 
+ bl[94] br[94] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_97 
+ bl[95] br[95] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_98 
+ bl[96] br[96] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_99 
+ bl[97] br[97] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_100 
+ bl[98] br[98] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_101 
+ bl[99] br[99] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_102 
+ bl[100] br[100] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_103 
+ bl[101] br[101] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_104 
+ bl[102] br[102] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_105 
+ bl[103] br[103] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_106 
+ bl[104] br[104] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_107 
+ bl[105] br[105] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_108 
+ bl[106] br[106] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_109 
+ bl[107] br[107] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_110 
+ bl[108] br[108] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_111 
+ bl[109] br[109] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_112 
+ bl[110] br[110] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_113 
+ bl[111] br[111] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_114 
+ bl[112] br[112] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_115 
+ bl[113] br[113] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_116 
+ bl[114] br[114] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_117 
+ bl[115] br[115] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_118 
+ bl[116] br[116] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_119 
+ bl[117] br[117] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_120 
+ bl[118] br[118] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_121 
+ bl[119] br[119] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_122 
+ bl[120] br[120] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_123 
+ bl[121] br[121] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_124 
+ bl[122] br[122] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_125 
+ bl[123] br[123] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_126 
+ bl[124] br[124] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_127 
+ bl[125] br[125] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_128 
+ bl[126] br[126] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_129 
+ bl[127] br[127] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_130 
+ bl[128] br[128] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_131 
+ bl[129] br[129] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_132 
+ bl[130] br[130] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_133 
+ bl[131] br[131] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_134 
+ bl[132] br[132] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_135 
+ bl[133] br[133] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_136 
+ bl[134] br[134] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_137 
+ bl[135] br[135] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_138 
+ bl[136] br[136] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_139 
+ bl[137] br[137] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_140 
+ bl[138] br[138] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_141 
+ bl[139] br[139] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_142 
+ bl[140] br[140] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_143 
+ bl[141] br[141] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_144 
+ bl[142] br[142] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_145 
+ bl[143] br[143] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_146 
+ bl[144] br[144] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_147 
+ bl[145] br[145] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_148 
+ bl[146] br[146] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_149 
+ bl[147] br[147] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_150 
+ bl[148] br[148] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_151 
+ bl[149] br[149] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_152 
+ bl[150] br[150] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_153 
+ bl[151] br[151] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_154 
+ bl[152] br[152] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_155 
+ bl[153] br[153] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_156 
+ bl[154] br[154] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_157 
+ bl[155] br[155] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_158 
+ bl[156] br[156] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_159 
+ bl[157] br[157] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_160 
+ bl[158] br[158] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_161 
+ bl[159] br[159] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_162 
+ bl[160] br[160] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_163 
+ bl[161] br[161] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_164 
+ bl[162] br[162] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_165 
+ bl[163] br[163] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_166 
+ bl[164] br[164] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_167 
+ bl[165] br[165] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_168 
+ bl[166] br[166] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_169 
+ bl[167] br[167] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_170 
+ bl[168] br[168] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_171 
+ bl[169] br[169] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_172 
+ bl[170] br[170] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_173 
+ bl[171] br[171] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_174 
+ bl[172] br[172] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_175 
+ bl[173] br[173] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_176 
+ bl[174] br[174] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_177 
+ bl[175] br[175] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_178 
+ bl[176] br[176] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_179 
+ bl[177] br[177] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_180 
+ bl[178] br[178] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_181 
+ bl[179] br[179] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_182 
+ bl[180] br[180] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_183 
+ bl[181] br[181] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_184 
+ bl[182] br[182] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_185 
+ bl[183] br[183] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_186 
+ bl[184] br[184] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_187 
+ bl[185] br[185] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_188 
+ bl[186] br[186] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_189 
+ bl[187] br[187] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_190 
+ bl[188] br[188] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_191 
+ bl[189] br[189] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_192 
+ bl[190] br[190] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_193 
+ bl[191] br[191] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_194 
+ bl[192] br[192] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_195 
+ bl[193] br[193] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_196 
+ bl[194] br[194] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_197 
+ bl[195] br[195] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_198 
+ bl[196] br[196] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_199 
+ bl[197] br[197] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_200 
+ bl[198] br[198] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_201 
+ bl[199] br[199] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_202 
+ bl[200] br[200] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_203 
+ bl[201] br[201] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_204 
+ bl[202] br[202] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_205 
+ bl[203] br[203] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_206 
+ bl[204] br[204] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_207 
+ bl[205] br[205] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_208 
+ bl[206] br[206] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_209 
+ bl[207] br[207] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_210 
+ bl[208] br[208] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_211 
+ bl[209] br[209] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_212 
+ bl[210] br[210] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_213 
+ bl[211] br[211] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_214 
+ bl[212] br[212] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_215 
+ bl[213] br[213] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_216 
+ bl[214] br[214] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_217 
+ bl[215] br[215] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_218 
+ bl[216] br[216] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_219 
+ bl[217] br[217] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_220 
+ bl[218] br[218] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_221 
+ bl[219] br[219] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_222 
+ bl[220] br[220] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_223 
+ bl[221] br[221] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_224 
+ bl[222] br[222] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_225 
+ bl[223] br[223] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_226 
+ bl[224] br[224] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_227 
+ bl[225] br[225] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_228 
+ bl[226] br[226] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_229 
+ bl[227] br[227] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_230 
+ bl[228] br[228] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_231 
+ bl[229] br[229] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_232 
+ bl[230] br[230] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_233 
+ bl[231] br[231] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_234 
+ bl[232] br[232] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_235 
+ bl[233] br[233] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_236 
+ bl[234] br[234] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_237 
+ bl[235] br[235] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_238 
+ bl[236] br[236] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_239 
+ bl[237] br[237] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_240 
+ bl[238] br[238] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_241 
+ bl[239] br[239] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_242 
+ bl[240] br[240] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_243 
+ bl[241] br[241] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_244 
+ bl[242] br[242] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_245 
+ bl[243] br[243] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_246 
+ bl[244] br[244] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_247 
+ bl[245] br[245] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_248 
+ bl[246] br[246] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_249 
+ bl[247] br[247] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_250 
+ bl[248] br[248] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_251 
+ bl[249] br[249] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_252 
+ bl[250] br[250] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_253 
+ bl[251] br[251] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_254 
+ bl[252] br[252] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_255 
+ bl[253] br[253] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_256 
+ bl[254] br[254] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_257 
+ bl[255] br[255] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_258 
+ vdd vdd vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_259 
+ vdd vdd vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_0 
+ vdd vdd vss vdd vpb vnb wl[121] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_123_1 
+ rbl rbr vss vdd vpb vnb wl[121] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_123_2 
+ bl[0] br[0] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_3 
+ bl[1] br[1] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_4 
+ bl[2] br[2] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_5 
+ bl[3] br[3] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_6 
+ bl[4] br[4] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_7 
+ bl[5] br[5] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_8 
+ bl[6] br[6] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_9 
+ bl[7] br[7] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_10 
+ bl[8] br[8] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_11 
+ bl[9] br[9] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_12 
+ bl[10] br[10] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_13 
+ bl[11] br[11] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_14 
+ bl[12] br[12] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_15 
+ bl[13] br[13] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_16 
+ bl[14] br[14] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_17 
+ bl[15] br[15] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_18 
+ bl[16] br[16] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_19 
+ bl[17] br[17] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_20 
+ bl[18] br[18] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_21 
+ bl[19] br[19] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_22 
+ bl[20] br[20] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_23 
+ bl[21] br[21] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_24 
+ bl[22] br[22] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_25 
+ bl[23] br[23] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_26 
+ bl[24] br[24] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_27 
+ bl[25] br[25] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_28 
+ bl[26] br[26] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_29 
+ bl[27] br[27] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_30 
+ bl[28] br[28] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_31 
+ bl[29] br[29] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_32 
+ bl[30] br[30] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_33 
+ bl[31] br[31] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_34 
+ bl[32] br[32] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_35 
+ bl[33] br[33] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_36 
+ bl[34] br[34] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_37 
+ bl[35] br[35] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_38 
+ bl[36] br[36] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_39 
+ bl[37] br[37] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_40 
+ bl[38] br[38] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_41 
+ bl[39] br[39] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_42 
+ bl[40] br[40] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_43 
+ bl[41] br[41] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_44 
+ bl[42] br[42] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_45 
+ bl[43] br[43] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_46 
+ bl[44] br[44] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_47 
+ bl[45] br[45] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_48 
+ bl[46] br[46] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_49 
+ bl[47] br[47] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_50 
+ bl[48] br[48] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_51 
+ bl[49] br[49] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_52 
+ bl[50] br[50] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_53 
+ bl[51] br[51] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_54 
+ bl[52] br[52] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_55 
+ bl[53] br[53] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_56 
+ bl[54] br[54] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_57 
+ bl[55] br[55] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_58 
+ bl[56] br[56] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_59 
+ bl[57] br[57] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_60 
+ bl[58] br[58] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_61 
+ bl[59] br[59] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_62 
+ bl[60] br[60] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_63 
+ bl[61] br[61] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_64 
+ bl[62] br[62] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_65 
+ bl[63] br[63] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_66 
+ bl[64] br[64] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_67 
+ bl[65] br[65] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_68 
+ bl[66] br[66] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_69 
+ bl[67] br[67] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_70 
+ bl[68] br[68] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_71 
+ bl[69] br[69] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_72 
+ bl[70] br[70] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_73 
+ bl[71] br[71] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_74 
+ bl[72] br[72] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_75 
+ bl[73] br[73] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_76 
+ bl[74] br[74] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_77 
+ bl[75] br[75] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_78 
+ bl[76] br[76] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_79 
+ bl[77] br[77] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_80 
+ bl[78] br[78] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_81 
+ bl[79] br[79] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_82 
+ bl[80] br[80] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_83 
+ bl[81] br[81] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_84 
+ bl[82] br[82] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_85 
+ bl[83] br[83] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_86 
+ bl[84] br[84] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_87 
+ bl[85] br[85] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_88 
+ bl[86] br[86] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_89 
+ bl[87] br[87] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_90 
+ bl[88] br[88] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_91 
+ bl[89] br[89] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_92 
+ bl[90] br[90] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_93 
+ bl[91] br[91] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_94 
+ bl[92] br[92] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_95 
+ bl[93] br[93] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_96 
+ bl[94] br[94] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_97 
+ bl[95] br[95] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_98 
+ bl[96] br[96] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_99 
+ bl[97] br[97] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_100 
+ bl[98] br[98] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_101 
+ bl[99] br[99] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_102 
+ bl[100] br[100] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_103 
+ bl[101] br[101] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_104 
+ bl[102] br[102] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_105 
+ bl[103] br[103] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_106 
+ bl[104] br[104] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_107 
+ bl[105] br[105] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_108 
+ bl[106] br[106] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_109 
+ bl[107] br[107] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_110 
+ bl[108] br[108] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_111 
+ bl[109] br[109] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_112 
+ bl[110] br[110] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_113 
+ bl[111] br[111] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_114 
+ bl[112] br[112] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_115 
+ bl[113] br[113] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_116 
+ bl[114] br[114] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_117 
+ bl[115] br[115] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_118 
+ bl[116] br[116] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_119 
+ bl[117] br[117] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_120 
+ bl[118] br[118] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_121 
+ bl[119] br[119] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_122 
+ bl[120] br[120] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_123 
+ bl[121] br[121] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_124 
+ bl[122] br[122] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_125 
+ bl[123] br[123] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_126 
+ bl[124] br[124] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_127 
+ bl[125] br[125] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_128 
+ bl[126] br[126] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_129 
+ bl[127] br[127] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_130 
+ bl[128] br[128] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_131 
+ bl[129] br[129] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_132 
+ bl[130] br[130] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_133 
+ bl[131] br[131] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_134 
+ bl[132] br[132] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_135 
+ bl[133] br[133] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_136 
+ bl[134] br[134] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_137 
+ bl[135] br[135] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_138 
+ bl[136] br[136] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_139 
+ bl[137] br[137] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_140 
+ bl[138] br[138] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_141 
+ bl[139] br[139] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_142 
+ bl[140] br[140] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_143 
+ bl[141] br[141] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_144 
+ bl[142] br[142] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_145 
+ bl[143] br[143] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_146 
+ bl[144] br[144] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_147 
+ bl[145] br[145] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_148 
+ bl[146] br[146] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_149 
+ bl[147] br[147] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_150 
+ bl[148] br[148] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_151 
+ bl[149] br[149] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_152 
+ bl[150] br[150] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_153 
+ bl[151] br[151] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_154 
+ bl[152] br[152] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_155 
+ bl[153] br[153] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_156 
+ bl[154] br[154] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_157 
+ bl[155] br[155] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_158 
+ bl[156] br[156] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_159 
+ bl[157] br[157] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_160 
+ bl[158] br[158] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_161 
+ bl[159] br[159] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_162 
+ bl[160] br[160] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_163 
+ bl[161] br[161] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_164 
+ bl[162] br[162] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_165 
+ bl[163] br[163] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_166 
+ bl[164] br[164] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_167 
+ bl[165] br[165] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_168 
+ bl[166] br[166] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_169 
+ bl[167] br[167] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_170 
+ bl[168] br[168] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_171 
+ bl[169] br[169] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_172 
+ bl[170] br[170] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_173 
+ bl[171] br[171] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_174 
+ bl[172] br[172] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_175 
+ bl[173] br[173] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_176 
+ bl[174] br[174] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_177 
+ bl[175] br[175] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_178 
+ bl[176] br[176] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_179 
+ bl[177] br[177] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_180 
+ bl[178] br[178] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_181 
+ bl[179] br[179] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_182 
+ bl[180] br[180] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_183 
+ bl[181] br[181] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_184 
+ bl[182] br[182] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_185 
+ bl[183] br[183] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_186 
+ bl[184] br[184] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_187 
+ bl[185] br[185] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_188 
+ bl[186] br[186] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_189 
+ bl[187] br[187] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_190 
+ bl[188] br[188] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_191 
+ bl[189] br[189] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_192 
+ bl[190] br[190] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_193 
+ bl[191] br[191] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_194 
+ bl[192] br[192] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_195 
+ bl[193] br[193] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_196 
+ bl[194] br[194] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_197 
+ bl[195] br[195] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_198 
+ bl[196] br[196] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_199 
+ bl[197] br[197] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_200 
+ bl[198] br[198] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_201 
+ bl[199] br[199] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_202 
+ bl[200] br[200] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_203 
+ bl[201] br[201] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_204 
+ bl[202] br[202] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_205 
+ bl[203] br[203] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_206 
+ bl[204] br[204] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_207 
+ bl[205] br[205] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_208 
+ bl[206] br[206] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_209 
+ bl[207] br[207] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_210 
+ bl[208] br[208] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_211 
+ bl[209] br[209] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_212 
+ bl[210] br[210] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_213 
+ bl[211] br[211] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_214 
+ bl[212] br[212] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_215 
+ bl[213] br[213] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_216 
+ bl[214] br[214] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_217 
+ bl[215] br[215] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_218 
+ bl[216] br[216] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_219 
+ bl[217] br[217] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_220 
+ bl[218] br[218] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_221 
+ bl[219] br[219] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_222 
+ bl[220] br[220] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_223 
+ bl[221] br[221] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_224 
+ bl[222] br[222] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_225 
+ bl[223] br[223] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_226 
+ bl[224] br[224] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_227 
+ bl[225] br[225] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_228 
+ bl[226] br[226] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_229 
+ bl[227] br[227] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_230 
+ bl[228] br[228] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_231 
+ bl[229] br[229] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_232 
+ bl[230] br[230] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_233 
+ bl[231] br[231] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_234 
+ bl[232] br[232] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_235 
+ bl[233] br[233] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_236 
+ bl[234] br[234] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_237 
+ bl[235] br[235] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_238 
+ bl[236] br[236] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_239 
+ bl[237] br[237] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_240 
+ bl[238] br[238] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_241 
+ bl[239] br[239] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_242 
+ bl[240] br[240] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_243 
+ bl[241] br[241] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_244 
+ bl[242] br[242] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_245 
+ bl[243] br[243] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_246 
+ bl[244] br[244] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_247 
+ bl[245] br[245] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_248 
+ bl[246] br[246] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_249 
+ bl[247] br[247] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_250 
+ bl[248] br[248] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_251 
+ bl[249] br[249] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_252 
+ bl[250] br[250] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_253 
+ bl[251] br[251] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_254 
+ bl[252] br[252] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_255 
+ bl[253] br[253] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_256 
+ bl[254] br[254] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_257 
+ bl[255] br[255] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_258 
+ vdd vdd vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_259 
+ vdd vdd vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_0 
+ vdd vdd vss vdd vpb vnb wl[122] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_124_1 
+ rbl rbr vss vdd vpb vnb wl[122] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_124_2 
+ bl[0] br[0] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_3 
+ bl[1] br[1] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_4 
+ bl[2] br[2] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_5 
+ bl[3] br[3] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_6 
+ bl[4] br[4] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_7 
+ bl[5] br[5] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_8 
+ bl[6] br[6] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_9 
+ bl[7] br[7] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_10 
+ bl[8] br[8] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_11 
+ bl[9] br[9] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_12 
+ bl[10] br[10] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_13 
+ bl[11] br[11] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_14 
+ bl[12] br[12] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_15 
+ bl[13] br[13] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_16 
+ bl[14] br[14] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_17 
+ bl[15] br[15] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_18 
+ bl[16] br[16] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_19 
+ bl[17] br[17] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_20 
+ bl[18] br[18] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_21 
+ bl[19] br[19] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_22 
+ bl[20] br[20] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_23 
+ bl[21] br[21] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_24 
+ bl[22] br[22] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_25 
+ bl[23] br[23] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_26 
+ bl[24] br[24] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_27 
+ bl[25] br[25] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_28 
+ bl[26] br[26] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_29 
+ bl[27] br[27] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_30 
+ bl[28] br[28] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_31 
+ bl[29] br[29] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_32 
+ bl[30] br[30] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_33 
+ bl[31] br[31] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_34 
+ bl[32] br[32] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_35 
+ bl[33] br[33] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_36 
+ bl[34] br[34] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_37 
+ bl[35] br[35] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_38 
+ bl[36] br[36] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_39 
+ bl[37] br[37] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_40 
+ bl[38] br[38] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_41 
+ bl[39] br[39] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_42 
+ bl[40] br[40] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_43 
+ bl[41] br[41] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_44 
+ bl[42] br[42] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_45 
+ bl[43] br[43] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_46 
+ bl[44] br[44] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_47 
+ bl[45] br[45] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_48 
+ bl[46] br[46] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_49 
+ bl[47] br[47] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_50 
+ bl[48] br[48] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_51 
+ bl[49] br[49] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_52 
+ bl[50] br[50] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_53 
+ bl[51] br[51] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_54 
+ bl[52] br[52] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_55 
+ bl[53] br[53] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_56 
+ bl[54] br[54] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_57 
+ bl[55] br[55] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_58 
+ bl[56] br[56] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_59 
+ bl[57] br[57] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_60 
+ bl[58] br[58] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_61 
+ bl[59] br[59] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_62 
+ bl[60] br[60] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_63 
+ bl[61] br[61] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_64 
+ bl[62] br[62] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_65 
+ bl[63] br[63] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_66 
+ bl[64] br[64] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_67 
+ bl[65] br[65] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_68 
+ bl[66] br[66] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_69 
+ bl[67] br[67] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_70 
+ bl[68] br[68] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_71 
+ bl[69] br[69] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_72 
+ bl[70] br[70] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_73 
+ bl[71] br[71] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_74 
+ bl[72] br[72] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_75 
+ bl[73] br[73] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_76 
+ bl[74] br[74] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_77 
+ bl[75] br[75] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_78 
+ bl[76] br[76] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_79 
+ bl[77] br[77] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_80 
+ bl[78] br[78] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_81 
+ bl[79] br[79] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_82 
+ bl[80] br[80] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_83 
+ bl[81] br[81] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_84 
+ bl[82] br[82] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_85 
+ bl[83] br[83] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_86 
+ bl[84] br[84] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_87 
+ bl[85] br[85] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_88 
+ bl[86] br[86] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_89 
+ bl[87] br[87] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_90 
+ bl[88] br[88] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_91 
+ bl[89] br[89] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_92 
+ bl[90] br[90] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_93 
+ bl[91] br[91] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_94 
+ bl[92] br[92] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_95 
+ bl[93] br[93] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_96 
+ bl[94] br[94] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_97 
+ bl[95] br[95] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_98 
+ bl[96] br[96] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_99 
+ bl[97] br[97] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_100 
+ bl[98] br[98] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_101 
+ bl[99] br[99] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_102 
+ bl[100] br[100] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_103 
+ bl[101] br[101] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_104 
+ bl[102] br[102] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_105 
+ bl[103] br[103] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_106 
+ bl[104] br[104] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_107 
+ bl[105] br[105] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_108 
+ bl[106] br[106] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_109 
+ bl[107] br[107] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_110 
+ bl[108] br[108] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_111 
+ bl[109] br[109] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_112 
+ bl[110] br[110] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_113 
+ bl[111] br[111] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_114 
+ bl[112] br[112] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_115 
+ bl[113] br[113] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_116 
+ bl[114] br[114] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_117 
+ bl[115] br[115] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_118 
+ bl[116] br[116] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_119 
+ bl[117] br[117] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_120 
+ bl[118] br[118] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_121 
+ bl[119] br[119] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_122 
+ bl[120] br[120] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_123 
+ bl[121] br[121] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_124 
+ bl[122] br[122] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_125 
+ bl[123] br[123] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_126 
+ bl[124] br[124] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_127 
+ bl[125] br[125] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_128 
+ bl[126] br[126] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_129 
+ bl[127] br[127] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_130 
+ bl[128] br[128] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_131 
+ bl[129] br[129] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_132 
+ bl[130] br[130] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_133 
+ bl[131] br[131] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_134 
+ bl[132] br[132] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_135 
+ bl[133] br[133] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_136 
+ bl[134] br[134] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_137 
+ bl[135] br[135] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_138 
+ bl[136] br[136] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_139 
+ bl[137] br[137] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_140 
+ bl[138] br[138] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_141 
+ bl[139] br[139] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_142 
+ bl[140] br[140] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_143 
+ bl[141] br[141] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_144 
+ bl[142] br[142] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_145 
+ bl[143] br[143] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_146 
+ bl[144] br[144] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_147 
+ bl[145] br[145] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_148 
+ bl[146] br[146] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_149 
+ bl[147] br[147] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_150 
+ bl[148] br[148] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_151 
+ bl[149] br[149] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_152 
+ bl[150] br[150] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_153 
+ bl[151] br[151] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_154 
+ bl[152] br[152] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_155 
+ bl[153] br[153] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_156 
+ bl[154] br[154] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_157 
+ bl[155] br[155] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_158 
+ bl[156] br[156] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_159 
+ bl[157] br[157] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_160 
+ bl[158] br[158] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_161 
+ bl[159] br[159] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_162 
+ bl[160] br[160] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_163 
+ bl[161] br[161] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_164 
+ bl[162] br[162] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_165 
+ bl[163] br[163] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_166 
+ bl[164] br[164] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_167 
+ bl[165] br[165] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_168 
+ bl[166] br[166] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_169 
+ bl[167] br[167] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_170 
+ bl[168] br[168] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_171 
+ bl[169] br[169] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_172 
+ bl[170] br[170] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_173 
+ bl[171] br[171] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_174 
+ bl[172] br[172] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_175 
+ bl[173] br[173] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_176 
+ bl[174] br[174] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_177 
+ bl[175] br[175] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_178 
+ bl[176] br[176] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_179 
+ bl[177] br[177] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_180 
+ bl[178] br[178] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_181 
+ bl[179] br[179] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_182 
+ bl[180] br[180] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_183 
+ bl[181] br[181] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_184 
+ bl[182] br[182] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_185 
+ bl[183] br[183] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_186 
+ bl[184] br[184] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_187 
+ bl[185] br[185] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_188 
+ bl[186] br[186] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_189 
+ bl[187] br[187] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_190 
+ bl[188] br[188] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_191 
+ bl[189] br[189] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_192 
+ bl[190] br[190] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_193 
+ bl[191] br[191] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_194 
+ bl[192] br[192] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_195 
+ bl[193] br[193] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_196 
+ bl[194] br[194] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_197 
+ bl[195] br[195] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_198 
+ bl[196] br[196] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_199 
+ bl[197] br[197] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_200 
+ bl[198] br[198] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_201 
+ bl[199] br[199] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_202 
+ bl[200] br[200] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_203 
+ bl[201] br[201] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_204 
+ bl[202] br[202] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_205 
+ bl[203] br[203] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_206 
+ bl[204] br[204] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_207 
+ bl[205] br[205] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_208 
+ bl[206] br[206] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_209 
+ bl[207] br[207] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_210 
+ bl[208] br[208] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_211 
+ bl[209] br[209] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_212 
+ bl[210] br[210] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_213 
+ bl[211] br[211] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_214 
+ bl[212] br[212] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_215 
+ bl[213] br[213] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_216 
+ bl[214] br[214] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_217 
+ bl[215] br[215] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_218 
+ bl[216] br[216] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_219 
+ bl[217] br[217] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_220 
+ bl[218] br[218] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_221 
+ bl[219] br[219] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_222 
+ bl[220] br[220] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_223 
+ bl[221] br[221] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_224 
+ bl[222] br[222] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_225 
+ bl[223] br[223] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_226 
+ bl[224] br[224] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_227 
+ bl[225] br[225] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_228 
+ bl[226] br[226] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_229 
+ bl[227] br[227] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_230 
+ bl[228] br[228] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_231 
+ bl[229] br[229] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_232 
+ bl[230] br[230] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_233 
+ bl[231] br[231] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_234 
+ bl[232] br[232] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_235 
+ bl[233] br[233] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_236 
+ bl[234] br[234] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_237 
+ bl[235] br[235] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_238 
+ bl[236] br[236] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_239 
+ bl[237] br[237] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_240 
+ bl[238] br[238] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_241 
+ bl[239] br[239] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_242 
+ bl[240] br[240] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_243 
+ bl[241] br[241] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_244 
+ bl[242] br[242] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_245 
+ bl[243] br[243] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_246 
+ bl[244] br[244] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_247 
+ bl[245] br[245] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_248 
+ bl[246] br[246] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_249 
+ bl[247] br[247] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_250 
+ bl[248] br[248] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_251 
+ bl[249] br[249] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_252 
+ bl[250] br[250] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_253 
+ bl[251] br[251] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_254 
+ bl[252] br[252] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_255 
+ bl[253] br[253] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_256 
+ bl[254] br[254] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_257 
+ bl[255] br[255] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_258 
+ vdd vdd vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_259 
+ vdd vdd vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_0 
+ vdd vdd vss vdd vpb vnb wl[123] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_125_1 
+ rbl rbr vss vdd vpb vnb wl[123] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_125_2 
+ bl[0] br[0] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_3 
+ bl[1] br[1] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_4 
+ bl[2] br[2] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_5 
+ bl[3] br[3] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_6 
+ bl[4] br[4] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_7 
+ bl[5] br[5] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_8 
+ bl[6] br[6] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_9 
+ bl[7] br[7] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_10 
+ bl[8] br[8] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_11 
+ bl[9] br[9] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_12 
+ bl[10] br[10] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_13 
+ bl[11] br[11] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_14 
+ bl[12] br[12] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_15 
+ bl[13] br[13] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_16 
+ bl[14] br[14] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_17 
+ bl[15] br[15] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_18 
+ bl[16] br[16] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_19 
+ bl[17] br[17] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_20 
+ bl[18] br[18] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_21 
+ bl[19] br[19] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_22 
+ bl[20] br[20] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_23 
+ bl[21] br[21] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_24 
+ bl[22] br[22] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_25 
+ bl[23] br[23] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_26 
+ bl[24] br[24] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_27 
+ bl[25] br[25] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_28 
+ bl[26] br[26] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_29 
+ bl[27] br[27] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_30 
+ bl[28] br[28] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_31 
+ bl[29] br[29] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_32 
+ bl[30] br[30] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_33 
+ bl[31] br[31] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_34 
+ bl[32] br[32] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_35 
+ bl[33] br[33] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_36 
+ bl[34] br[34] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_37 
+ bl[35] br[35] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_38 
+ bl[36] br[36] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_39 
+ bl[37] br[37] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_40 
+ bl[38] br[38] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_41 
+ bl[39] br[39] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_42 
+ bl[40] br[40] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_43 
+ bl[41] br[41] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_44 
+ bl[42] br[42] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_45 
+ bl[43] br[43] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_46 
+ bl[44] br[44] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_47 
+ bl[45] br[45] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_48 
+ bl[46] br[46] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_49 
+ bl[47] br[47] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_50 
+ bl[48] br[48] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_51 
+ bl[49] br[49] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_52 
+ bl[50] br[50] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_53 
+ bl[51] br[51] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_54 
+ bl[52] br[52] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_55 
+ bl[53] br[53] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_56 
+ bl[54] br[54] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_57 
+ bl[55] br[55] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_58 
+ bl[56] br[56] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_59 
+ bl[57] br[57] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_60 
+ bl[58] br[58] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_61 
+ bl[59] br[59] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_62 
+ bl[60] br[60] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_63 
+ bl[61] br[61] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_64 
+ bl[62] br[62] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_65 
+ bl[63] br[63] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_66 
+ bl[64] br[64] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_67 
+ bl[65] br[65] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_68 
+ bl[66] br[66] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_69 
+ bl[67] br[67] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_70 
+ bl[68] br[68] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_71 
+ bl[69] br[69] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_72 
+ bl[70] br[70] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_73 
+ bl[71] br[71] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_74 
+ bl[72] br[72] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_75 
+ bl[73] br[73] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_76 
+ bl[74] br[74] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_77 
+ bl[75] br[75] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_78 
+ bl[76] br[76] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_79 
+ bl[77] br[77] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_80 
+ bl[78] br[78] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_81 
+ bl[79] br[79] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_82 
+ bl[80] br[80] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_83 
+ bl[81] br[81] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_84 
+ bl[82] br[82] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_85 
+ bl[83] br[83] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_86 
+ bl[84] br[84] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_87 
+ bl[85] br[85] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_88 
+ bl[86] br[86] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_89 
+ bl[87] br[87] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_90 
+ bl[88] br[88] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_91 
+ bl[89] br[89] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_92 
+ bl[90] br[90] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_93 
+ bl[91] br[91] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_94 
+ bl[92] br[92] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_95 
+ bl[93] br[93] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_96 
+ bl[94] br[94] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_97 
+ bl[95] br[95] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_98 
+ bl[96] br[96] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_99 
+ bl[97] br[97] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_100 
+ bl[98] br[98] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_101 
+ bl[99] br[99] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_102 
+ bl[100] br[100] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_103 
+ bl[101] br[101] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_104 
+ bl[102] br[102] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_105 
+ bl[103] br[103] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_106 
+ bl[104] br[104] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_107 
+ bl[105] br[105] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_108 
+ bl[106] br[106] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_109 
+ bl[107] br[107] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_110 
+ bl[108] br[108] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_111 
+ bl[109] br[109] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_112 
+ bl[110] br[110] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_113 
+ bl[111] br[111] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_114 
+ bl[112] br[112] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_115 
+ bl[113] br[113] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_116 
+ bl[114] br[114] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_117 
+ bl[115] br[115] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_118 
+ bl[116] br[116] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_119 
+ bl[117] br[117] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_120 
+ bl[118] br[118] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_121 
+ bl[119] br[119] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_122 
+ bl[120] br[120] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_123 
+ bl[121] br[121] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_124 
+ bl[122] br[122] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_125 
+ bl[123] br[123] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_126 
+ bl[124] br[124] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_127 
+ bl[125] br[125] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_128 
+ bl[126] br[126] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_129 
+ bl[127] br[127] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_130 
+ bl[128] br[128] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_131 
+ bl[129] br[129] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_132 
+ bl[130] br[130] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_133 
+ bl[131] br[131] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_134 
+ bl[132] br[132] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_135 
+ bl[133] br[133] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_136 
+ bl[134] br[134] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_137 
+ bl[135] br[135] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_138 
+ bl[136] br[136] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_139 
+ bl[137] br[137] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_140 
+ bl[138] br[138] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_141 
+ bl[139] br[139] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_142 
+ bl[140] br[140] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_143 
+ bl[141] br[141] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_144 
+ bl[142] br[142] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_145 
+ bl[143] br[143] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_146 
+ bl[144] br[144] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_147 
+ bl[145] br[145] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_148 
+ bl[146] br[146] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_149 
+ bl[147] br[147] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_150 
+ bl[148] br[148] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_151 
+ bl[149] br[149] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_152 
+ bl[150] br[150] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_153 
+ bl[151] br[151] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_154 
+ bl[152] br[152] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_155 
+ bl[153] br[153] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_156 
+ bl[154] br[154] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_157 
+ bl[155] br[155] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_158 
+ bl[156] br[156] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_159 
+ bl[157] br[157] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_160 
+ bl[158] br[158] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_161 
+ bl[159] br[159] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_162 
+ bl[160] br[160] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_163 
+ bl[161] br[161] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_164 
+ bl[162] br[162] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_165 
+ bl[163] br[163] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_166 
+ bl[164] br[164] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_167 
+ bl[165] br[165] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_168 
+ bl[166] br[166] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_169 
+ bl[167] br[167] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_170 
+ bl[168] br[168] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_171 
+ bl[169] br[169] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_172 
+ bl[170] br[170] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_173 
+ bl[171] br[171] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_174 
+ bl[172] br[172] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_175 
+ bl[173] br[173] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_176 
+ bl[174] br[174] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_177 
+ bl[175] br[175] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_178 
+ bl[176] br[176] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_179 
+ bl[177] br[177] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_180 
+ bl[178] br[178] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_181 
+ bl[179] br[179] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_182 
+ bl[180] br[180] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_183 
+ bl[181] br[181] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_184 
+ bl[182] br[182] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_185 
+ bl[183] br[183] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_186 
+ bl[184] br[184] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_187 
+ bl[185] br[185] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_188 
+ bl[186] br[186] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_189 
+ bl[187] br[187] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_190 
+ bl[188] br[188] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_191 
+ bl[189] br[189] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_192 
+ bl[190] br[190] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_193 
+ bl[191] br[191] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_194 
+ bl[192] br[192] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_195 
+ bl[193] br[193] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_196 
+ bl[194] br[194] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_197 
+ bl[195] br[195] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_198 
+ bl[196] br[196] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_199 
+ bl[197] br[197] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_200 
+ bl[198] br[198] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_201 
+ bl[199] br[199] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_202 
+ bl[200] br[200] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_203 
+ bl[201] br[201] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_204 
+ bl[202] br[202] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_205 
+ bl[203] br[203] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_206 
+ bl[204] br[204] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_207 
+ bl[205] br[205] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_208 
+ bl[206] br[206] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_209 
+ bl[207] br[207] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_210 
+ bl[208] br[208] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_211 
+ bl[209] br[209] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_212 
+ bl[210] br[210] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_213 
+ bl[211] br[211] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_214 
+ bl[212] br[212] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_215 
+ bl[213] br[213] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_216 
+ bl[214] br[214] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_217 
+ bl[215] br[215] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_218 
+ bl[216] br[216] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_219 
+ bl[217] br[217] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_220 
+ bl[218] br[218] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_221 
+ bl[219] br[219] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_222 
+ bl[220] br[220] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_223 
+ bl[221] br[221] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_224 
+ bl[222] br[222] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_225 
+ bl[223] br[223] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_226 
+ bl[224] br[224] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_227 
+ bl[225] br[225] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_228 
+ bl[226] br[226] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_229 
+ bl[227] br[227] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_230 
+ bl[228] br[228] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_231 
+ bl[229] br[229] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_232 
+ bl[230] br[230] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_233 
+ bl[231] br[231] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_234 
+ bl[232] br[232] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_235 
+ bl[233] br[233] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_236 
+ bl[234] br[234] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_237 
+ bl[235] br[235] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_238 
+ bl[236] br[236] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_239 
+ bl[237] br[237] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_240 
+ bl[238] br[238] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_241 
+ bl[239] br[239] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_242 
+ bl[240] br[240] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_243 
+ bl[241] br[241] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_244 
+ bl[242] br[242] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_245 
+ bl[243] br[243] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_246 
+ bl[244] br[244] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_247 
+ bl[245] br[245] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_248 
+ bl[246] br[246] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_249 
+ bl[247] br[247] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_250 
+ bl[248] br[248] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_251 
+ bl[249] br[249] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_252 
+ bl[250] br[250] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_253 
+ bl[251] br[251] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_254 
+ bl[252] br[252] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_255 
+ bl[253] br[253] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_256 
+ bl[254] br[254] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_257 
+ bl[255] br[255] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_258 
+ vdd vdd vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_259 
+ vdd vdd vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_0 
+ vdd vdd vss vdd vpb vnb wl[124] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_126_1 
+ rbl rbr vss vdd vpb vnb wl[124] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_126_2 
+ bl[0] br[0] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_3 
+ bl[1] br[1] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_4 
+ bl[2] br[2] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_5 
+ bl[3] br[3] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_6 
+ bl[4] br[4] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_7 
+ bl[5] br[5] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_8 
+ bl[6] br[6] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_9 
+ bl[7] br[7] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_10 
+ bl[8] br[8] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_11 
+ bl[9] br[9] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_12 
+ bl[10] br[10] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_13 
+ bl[11] br[11] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_14 
+ bl[12] br[12] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_15 
+ bl[13] br[13] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_16 
+ bl[14] br[14] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_17 
+ bl[15] br[15] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_18 
+ bl[16] br[16] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_19 
+ bl[17] br[17] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_20 
+ bl[18] br[18] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_21 
+ bl[19] br[19] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_22 
+ bl[20] br[20] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_23 
+ bl[21] br[21] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_24 
+ bl[22] br[22] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_25 
+ bl[23] br[23] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_26 
+ bl[24] br[24] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_27 
+ bl[25] br[25] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_28 
+ bl[26] br[26] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_29 
+ bl[27] br[27] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_30 
+ bl[28] br[28] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_31 
+ bl[29] br[29] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_32 
+ bl[30] br[30] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_33 
+ bl[31] br[31] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_34 
+ bl[32] br[32] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_35 
+ bl[33] br[33] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_36 
+ bl[34] br[34] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_37 
+ bl[35] br[35] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_38 
+ bl[36] br[36] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_39 
+ bl[37] br[37] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_40 
+ bl[38] br[38] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_41 
+ bl[39] br[39] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_42 
+ bl[40] br[40] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_43 
+ bl[41] br[41] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_44 
+ bl[42] br[42] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_45 
+ bl[43] br[43] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_46 
+ bl[44] br[44] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_47 
+ bl[45] br[45] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_48 
+ bl[46] br[46] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_49 
+ bl[47] br[47] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_50 
+ bl[48] br[48] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_51 
+ bl[49] br[49] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_52 
+ bl[50] br[50] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_53 
+ bl[51] br[51] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_54 
+ bl[52] br[52] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_55 
+ bl[53] br[53] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_56 
+ bl[54] br[54] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_57 
+ bl[55] br[55] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_58 
+ bl[56] br[56] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_59 
+ bl[57] br[57] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_60 
+ bl[58] br[58] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_61 
+ bl[59] br[59] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_62 
+ bl[60] br[60] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_63 
+ bl[61] br[61] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_64 
+ bl[62] br[62] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_65 
+ bl[63] br[63] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_66 
+ bl[64] br[64] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_67 
+ bl[65] br[65] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_68 
+ bl[66] br[66] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_69 
+ bl[67] br[67] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_70 
+ bl[68] br[68] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_71 
+ bl[69] br[69] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_72 
+ bl[70] br[70] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_73 
+ bl[71] br[71] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_74 
+ bl[72] br[72] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_75 
+ bl[73] br[73] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_76 
+ bl[74] br[74] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_77 
+ bl[75] br[75] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_78 
+ bl[76] br[76] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_79 
+ bl[77] br[77] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_80 
+ bl[78] br[78] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_81 
+ bl[79] br[79] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_82 
+ bl[80] br[80] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_83 
+ bl[81] br[81] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_84 
+ bl[82] br[82] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_85 
+ bl[83] br[83] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_86 
+ bl[84] br[84] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_87 
+ bl[85] br[85] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_88 
+ bl[86] br[86] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_89 
+ bl[87] br[87] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_90 
+ bl[88] br[88] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_91 
+ bl[89] br[89] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_92 
+ bl[90] br[90] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_93 
+ bl[91] br[91] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_94 
+ bl[92] br[92] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_95 
+ bl[93] br[93] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_96 
+ bl[94] br[94] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_97 
+ bl[95] br[95] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_98 
+ bl[96] br[96] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_99 
+ bl[97] br[97] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_100 
+ bl[98] br[98] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_101 
+ bl[99] br[99] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_102 
+ bl[100] br[100] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_103 
+ bl[101] br[101] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_104 
+ bl[102] br[102] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_105 
+ bl[103] br[103] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_106 
+ bl[104] br[104] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_107 
+ bl[105] br[105] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_108 
+ bl[106] br[106] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_109 
+ bl[107] br[107] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_110 
+ bl[108] br[108] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_111 
+ bl[109] br[109] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_112 
+ bl[110] br[110] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_113 
+ bl[111] br[111] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_114 
+ bl[112] br[112] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_115 
+ bl[113] br[113] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_116 
+ bl[114] br[114] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_117 
+ bl[115] br[115] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_118 
+ bl[116] br[116] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_119 
+ bl[117] br[117] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_120 
+ bl[118] br[118] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_121 
+ bl[119] br[119] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_122 
+ bl[120] br[120] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_123 
+ bl[121] br[121] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_124 
+ bl[122] br[122] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_125 
+ bl[123] br[123] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_126 
+ bl[124] br[124] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_127 
+ bl[125] br[125] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_128 
+ bl[126] br[126] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_129 
+ bl[127] br[127] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_130 
+ bl[128] br[128] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_131 
+ bl[129] br[129] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_132 
+ bl[130] br[130] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_133 
+ bl[131] br[131] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_134 
+ bl[132] br[132] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_135 
+ bl[133] br[133] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_136 
+ bl[134] br[134] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_137 
+ bl[135] br[135] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_138 
+ bl[136] br[136] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_139 
+ bl[137] br[137] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_140 
+ bl[138] br[138] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_141 
+ bl[139] br[139] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_142 
+ bl[140] br[140] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_143 
+ bl[141] br[141] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_144 
+ bl[142] br[142] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_145 
+ bl[143] br[143] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_146 
+ bl[144] br[144] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_147 
+ bl[145] br[145] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_148 
+ bl[146] br[146] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_149 
+ bl[147] br[147] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_150 
+ bl[148] br[148] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_151 
+ bl[149] br[149] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_152 
+ bl[150] br[150] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_153 
+ bl[151] br[151] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_154 
+ bl[152] br[152] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_155 
+ bl[153] br[153] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_156 
+ bl[154] br[154] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_157 
+ bl[155] br[155] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_158 
+ bl[156] br[156] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_159 
+ bl[157] br[157] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_160 
+ bl[158] br[158] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_161 
+ bl[159] br[159] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_162 
+ bl[160] br[160] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_163 
+ bl[161] br[161] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_164 
+ bl[162] br[162] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_165 
+ bl[163] br[163] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_166 
+ bl[164] br[164] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_167 
+ bl[165] br[165] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_168 
+ bl[166] br[166] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_169 
+ bl[167] br[167] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_170 
+ bl[168] br[168] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_171 
+ bl[169] br[169] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_172 
+ bl[170] br[170] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_173 
+ bl[171] br[171] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_174 
+ bl[172] br[172] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_175 
+ bl[173] br[173] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_176 
+ bl[174] br[174] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_177 
+ bl[175] br[175] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_178 
+ bl[176] br[176] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_179 
+ bl[177] br[177] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_180 
+ bl[178] br[178] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_181 
+ bl[179] br[179] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_182 
+ bl[180] br[180] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_183 
+ bl[181] br[181] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_184 
+ bl[182] br[182] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_185 
+ bl[183] br[183] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_186 
+ bl[184] br[184] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_187 
+ bl[185] br[185] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_188 
+ bl[186] br[186] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_189 
+ bl[187] br[187] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_190 
+ bl[188] br[188] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_191 
+ bl[189] br[189] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_192 
+ bl[190] br[190] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_193 
+ bl[191] br[191] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_194 
+ bl[192] br[192] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_195 
+ bl[193] br[193] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_196 
+ bl[194] br[194] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_197 
+ bl[195] br[195] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_198 
+ bl[196] br[196] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_199 
+ bl[197] br[197] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_200 
+ bl[198] br[198] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_201 
+ bl[199] br[199] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_202 
+ bl[200] br[200] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_203 
+ bl[201] br[201] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_204 
+ bl[202] br[202] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_205 
+ bl[203] br[203] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_206 
+ bl[204] br[204] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_207 
+ bl[205] br[205] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_208 
+ bl[206] br[206] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_209 
+ bl[207] br[207] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_210 
+ bl[208] br[208] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_211 
+ bl[209] br[209] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_212 
+ bl[210] br[210] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_213 
+ bl[211] br[211] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_214 
+ bl[212] br[212] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_215 
+ bl[213] br[213] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_216 
+ bl[214] br[214] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_217 
+ bl[215] br[215] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_218 
+ bl[216] br[216] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_219 
+ bl[217] br[217] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_220 
+ bl[218] br[218] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_221 
+ bl[219] br[219] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_222 
+ bl[220] br[220] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_223 
+ bl[221] br[221] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_224 
+ bl[222] br[222] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_225 
+ bl[223] br[223] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_226 
+ bl[224] br[224] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_227 
+ bl[225] br[225] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_228 
+ bl[226] br[226] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_229 
+ bl[227] br[227] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_230 
+ bl[228] br[228] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_231 
+ bl[229] br[229] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_232 
+ bl[230] br[230] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_233 
+ bl[231] br[231] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_234 
+ bl[232] br[232] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_235 
+ bl[233] br[233] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_236 
+ bl[234] br[234] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_237 
+ bl[235] br[235] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_238 
+ bl[236] br[236] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_239 
+ bl[237] br[237] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_240 
+ bl[238] br[238] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_241 
+ bl[239] br[239] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_242 
+ bl[240] br[240] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_243 
+ bl[241] br[241] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_244 
+ bl[242] br[242] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_245 
+ bl[243] br[243] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_246 
+ bl[244] br[244] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_247 
+ bl[245] br[245] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_248 
+ bl[246] br[246] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_249 
+ bl[247] br[247] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_250 
+ bl[248] br[248] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_251 
+ bl[249] br[249] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_252 
+ bl[250] br[250] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_253 
+ bl[251] br[251] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_254 
+ bl[252] br[252] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_255 
+ bl[253] br[253] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_256 
+ bl[254] br[254] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_257 
+ bl[255] br[255] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_258 
+ vdd vdd vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_259 
+ vdd vdd vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_0 
+ vdd vdd vss vdd vpb vnb wl[125] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_127_1 
+ rbl rbr vss vdd vpb vnb wl[125] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_127_2 
+ bl[0] br[0] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_3 
+ bl[1] br[1] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_4 
+ bl[2] br[2] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_5 
+ bl[3] br[3] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_6 
+ bl[4] br[4] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_7 
+ bl[5] br[5] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_8 
+ bl[6] br[6] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_9 
+ bl[7] br[7] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_10 
+ bl[8] br[8] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_11 
+ bl[9] br[9] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_12 
+ bl[10] br[10] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_13 
+ bl[11] br[11] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_14 
+ bl[12] br[12] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_15 
+ bl[13] br[13] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_16 
+ bl[14] br[14] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_17 
+ bl[15] br[15] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_18 
+ bl[16] br[16] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_19 
+ bl[17] br[17] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_20 
+ bl[18] br[18] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_21 
+ bl[19] br[19] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_22 
+ bl[20] br[20] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_23 
+ bl[21] br[21] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_24 
+ bl[22] br[22] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_25 
+ bl[23] br[23] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_26 
+ bl[24] br[24] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_27 
+ bl[25] br[25] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_28 
+ bl[26] br[26] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_29 
+ bl[27] br[27] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_30 
+ bl[28] br[28] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_31 
+ bl[29] br[29] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_32 
+ bl[30] br[30] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_33 
+ bl[31] br[31] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_34 
+ bl[32] br[32] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_35 
+ bl[33] br[33] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_36 
+ bl[34] br[34] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_37 
+ bl[35] br[35] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_38 
+ bl[36] br[36] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_39 
+ bl[37] br[37] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_40 
+ bl[38] br[38] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_41 
+ bl[39] br[39] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_42 
+ bl[40] br[40] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_43 
+ bl[41] br[41] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_44 
+ bl[42] br[42] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_45 
+ bl[43] br[43] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_46 
+ bl[44] br[44] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_47 
+ bl[45] br[45] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_48 
+ bl[46] br[46] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_49 
+ bl[47] br[47] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_50 
+ bl[48] br[48] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_51 
+ bl[49] br[49] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_52 
+ bl[50] br[50] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_53 
+ bl[51] br[51] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_54 
+ bl[52] br[52] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_55 
+ bl[53] br[53] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_56 
+ bl[54] br[54] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_57 
+ bl[55] br[55] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_58 
+ bl[56] br[56] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_59 
+ bl[57] br[57] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_60 
+ bl[58] br[58] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_61 
+ bl[59] br[59] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_62 
+ bl[60] br[60] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_63 
+ bl[61] br[61] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_64 
+ bl[62] br[62] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_65 
+ bl[63] br[63] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_66 
+ bl[64] br[64] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_67 
+ bl[65] br[65] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_68 
+ bl[66] br[66] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_69 
+ bl[67] br[67] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_70 
+ bl[68] br[68] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_71 
+ bl[69] br[69] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_72 
+ bl[70] br[70] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_73 
+ bl[71] br[71] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_74 
+ bl[72] br[72] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_75 
+ bl[73] br[73] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_76 
+ bl[74] br[74] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_77 
+ bl[75] br[75] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_78 
+ bl[76] br[76] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_79 
+ bl[77] br[77] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_80 
+ bl[78] br[78] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_81 
+ bl[79] br[79] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_82 
+ bl[80] br[80] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_83 
+ bl[81] br[81] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_84 
+ bl[82] br[82] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_85 
+ bl[83] br[83] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_86 
+ bl[84] br[84] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_87 
+ bl[85] br[85] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_88 
+ bl[86] br[86] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_89 
+ bl[87] br[87] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_90 
+ bl[88] br[88] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_91 
+ bl[89] br[89] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_92 
+ bl[90] br[90] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_93 
+ bl[91] br[91] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_94 
+ bl[92] br[92] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_95 
+ bl[93] br[93] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_96 
+ bl[94] br[94] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_97 
+ bl[95] br[95] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_98 
+ bl[96] br[96] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_99 
+ bl[97] br[97] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_100 
+ bl[98] br[98] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_101 
+ bl[99] br[99] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_102 
+ bl[100] br[100] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_103 
+ bl[101] br[101] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_104 
+ bl[102] br[102] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_105 
+ bl[103] br[103] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_106 
+ bl[104] br[104] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_107 
+ bl[105] br[105] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_108 
+ bl[106] br[106] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_109 
+ bl[107] br[107] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_110 
+ bl[108] br[108] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_111 
+ bl[109] br[109] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_112 
+ bl[110] br[110] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_113 
+ bl[111] br[111] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_114 
+ bl[112] br[112] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_115 
+ bl[113] br[113] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_116 
+ bl[114] br[114] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_117 
+ bl[115] br[115] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_118 
+ bl[116] br[116] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_119 
+ bl[117] br[117] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_120 
+ bl[118] br[118] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_121 
+ bl[119] br[119] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_122 
+ bl[120] br[120] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_123 
+ bl[121] br[121] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_124 
+ bl[122] br[122] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_125 
+ bl[123] br[123] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_126 
+ bl[124] br[124] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_127 
+ bl[125] br[125] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_128 
+ bl[126] br[126] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_129 
+ bl[127] br[127] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_130 
+ bl[128] br[128] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_131 
+ bl[129] br[129] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_132 
+ bl[130] br[130] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_133 
+ bl[131] br[131] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_134 
+ bl[132] br[132] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_135 
+ bl[133] br[133] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_136 
+ bl[134] br[134] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_137 
+ bl[135] br[135] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_138 
+ bl[136] br[136] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_139 
+ bl[137] br[137] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_140 
+ bl[138] br[138] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_141 
+ bl[139] br[139] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_142 
+ bl[140] br[140] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_143 
+ bl[141] br[141] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_144 
+ bl[142] br[142] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_145 
+ bl[143] br[143] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_146 
+ bl[144] br[144] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_147 
+ bl[145] br[145] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_148 
+ bl[146] br[146] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_149 
+ bl[147] br[147] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_150 
+ bl[148] br[148] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_151 
+ bl[149] br[149] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_152 
+ bl[150] br[150] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_153 
+ bl[151] br[151] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_154 
+ bl[152] br[152] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_155 
+ bl[153] br[153] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_156 
+ bl[154] br[154] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_157 
+ bl[155] br[155] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_158 
+ bl[156] br[156] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_159 
+ bl[157] br[157] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_160 
+ bl[158] br[158] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_161 
+ bl[159] br[159] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_162 
+ bl[160] br[160] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_163 
+ bl[161] br[161] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_164 
+ bl[162] br[162] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_165 
+ bl[163] br[163] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_166 
+ bl[164] br[164] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_167 
+ bl[165] br[165] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_168 
+ bl[166] br[166] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_169 
+ bl[167] br[167] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_170 
+ bl[168] br[168] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_171 
+ bl[169] br[169] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_172 
+ bl[170] br[170] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_173 
+ bl[171] br[171] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_174 
+ bl[172] br[172] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_175 
+ bl[173] br[173] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_176 
+ bl[174] br[174] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_177 
+ bl[175] br[175] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_178 
+ bl[176] br[176] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_179 
+ bl[177] br[177] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_180 
+ bl[178] br[178] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_181 
+ bl[179] br[179] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_182 
+ bl[180] br[180] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_183 
+ bl[181] br[181] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_184 
+ bl[182] br[182] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_185 
+ bl[183] br[183] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_186 
+ bl[184] br[184] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_187 
+ bl[185] br[185] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_188 
+ bl[186] br[186] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_189 
+ bl[187] br[187] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_190 
+ bl[188] br[188] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_191 
+ bl[189] br[189] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_192 
+ bl[190] br[190] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_193 
+ bl[191] br[191] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_194 
+ bl[192] br[192] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_195 
+ bl[193] br[193] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_196 
+ bl[194] br[194] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_197 
+ bl[195] br[195] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_198 
+ bl[196] br[196] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_199 
+ bl[197] br[197] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_200 
+ bl[198] br[198] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_201 
+ bl[199] br[199] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_202 
+ bl[200] br[200] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_203 
+ bl[201] br[201] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_204 
+ bl[202] br[202] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_205 
+ bl[203] br[203] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_206 
+ bl[204] br[204] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_207 
+ bl[205] br[205] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_208 
+ bl[206] br[206] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_209 
+ bl[207] br[207] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_210 
+ bl[208] br[208] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_211 
+ bl[209] br[209] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_212 
+ bl[210] br[210] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_213 
+ bl[211] br[211] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_214 
+ bl[212] br[212] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_215 
+ bl[213] br[213] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_216 
+ bl[214] br[214] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_217 
+ bl[215] br[215] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_218 
+ bl[216] br[216] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_219 
+ bl[217] br[217] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_220 
+ bl[218] br[218] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_221 
+ bl[219] br[219] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_222 
+ bl[220] br[220] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_223 
+ bl[221] br[221] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_224 
+ bl[222] br[222] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_225 
+ bl[223] br[223] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_226 
+ bl[224] br[224] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_227 
+ bl[225] br[225] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_228 
+ bl[226] br[226] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_229 
+ bl[227] br[227] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_230 
+ bl[228] br[228] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_231 
+ bl[229] br[229] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_232 
+ bl[230] br[230] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_233 
+ bl[231] br[231] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_234 
+ bl[232] br[232] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_235 
+ bl[233] br[233] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_236 
+ bl[234] br[234] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_237 
+ bl[235] br[235] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_238 
+ bl[236] br[236] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_239 
+ bl[237] br[237] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_240 
+ bl[238] br[238] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_241 
+ bl[239] br[239] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_242 
+ bl[240] br[240] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_243 
+ bl[241] br[241] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_244 
+ bl[242] br[242] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_245 
+ bl[243] br[243] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_246 
+ bl[244] br[244] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_247 
+ bl[245] br[245] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_248 
+ bl[246] br[246] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_249 
+ bl[247] br[247] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_250 
+ bl[248] br[248] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_251 
+ bl[249] br[249] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_252 
+ bl[250] br[250] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_253 
+ bl[251] br[251] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_254 
+ bl[252] br[252] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_255 
+ bl[253] br[253] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_256 
+ bl[254] br[254] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_257 
+ bl[255] br[255] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_258 
+ vdd vdd vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_259 
+ vdd vdd vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_0 
+ vdd vdd vss vdd vpb vnb wl[126] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_128_1 
+ rbl rbr vss vdd vpb vnb wl[126] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_128_2 
+ bl[0] br[0] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_3 
+ bl[1] br[1] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_4 
+ bl[2] br[2] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_5 
+ bl[3] br[3] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_6 
+ bl[4] br[4] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_7 
+ bl[5] br[5] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_8 
+ bl[6] br[6] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_9 
+ bl[7] br[7] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_10 
+ bl[8] br[8] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_11 
+ bl[9] br[9] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_12 
+ bl[10] br[10] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_13 
+ bl[11] br[11] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_14 
+ bl[12] br[12] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_15 
+ bl[13] br[13] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_16 
+ bl[14] br[14] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_17 
+ bl[15] br[15] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_18 
+ bl[16] br[16] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_19 
+ bl[17] br[17] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_20 
+ bl[18] br[18] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_21 
+ bl[19] br[19] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_22 
+ bl[20] br[20] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_23 
+ bl[21] br[21] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_24 
+ bl[22] br[22] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_25 
+ bl[23] br[23] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_26 
+ bl[24] br[24] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_27 
+ bl[25] br[25] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_28 
+ bl[26] br[26] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_29 
+ bl[27] br[27] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_30 
+ bl[28] br[28] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_31 
+ bl[29] br[29] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_32 
+ bl[30] br[30] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_33 
+ bl[31] br[31] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_34 
+ bl[32] br[32] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_35 
+ bl[33] br[33] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_36 
+ bl[34] br[34] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_37 
+ bl[35] br[35] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_38 
+ bl[36] br[36] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_39 
+ bl[37] br[37] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_40 
+ bl[38] br[38] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_41 
+ bl[39] br[39] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_42 
+ bl[40] br[40] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_43 
+ bl[41] br[41] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_44 
+ bl[42] br[42] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_45 
+ bl[43] br[43] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_46 
+ bl[44] br[44] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_47 
+ bl[45] br[45] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_48 
+ bl[46] br[46] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_49 
+ bl[47] br[47] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_50 
+ bl[48] br[48] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_51 
+ bl[49] br[49] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_52 
+ bl[50] br[50] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_53 
+ bl[51] br[51] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_54 
+ bl[52] br[52] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_55 
+ bl[53] br[53] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_56 
+ bl[54] br[54] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_57 
+ bl[55] br[55] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_58 
+ bl[56] br[56] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_59 
+ bl[57] br[57] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_60 
+ bl[58] br[58] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_61 
+ bl[59] br[59] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_62 
+ bl[60] br[60] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_63 
+ bl[61] br[61] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_64 
+ bl[62] br[62] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_65 
+ bl[63] br[63] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_66 
+ bl[64] br[64] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_67 
+ bl[65] br[65] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_68 
+ bl[66] br[66] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_69 
+ bl[67] br[67] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_70 
+ bl[68] br[68] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_71 
+ bl[69] br[69] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_72 
+ bl[70] br[70] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_73 
+ bl[71] br[71] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_74 
+ bl[72] br[72] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_75 
+ bl[73] br[73] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_76 
+ bl[74] br[74] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_77 
+ bl[75] br[75] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_78 
+ bl[76] br[76] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_79 
+ bl[77] br[77] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_80 
+ bl[78] br[78] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_81 
+ bl[79] br[79] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_82 
+ bl[80] br[80] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_83 
+ bl[81] br[81] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_84 
+ bl[82] br[82] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_85 
+ bl[83] br[83] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_86 
+ bl[84] br[84] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_87 
+ bl[85] br[85] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_88 
+ bl[86] br[86] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_89 
+ bl[87] br[87] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_90 
+ bl[88] br[88] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_91 
+ bl[89] br[89] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_92 
+ bl[90] br[90] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_93 
+ bl[91] br[91] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_94 
+ bl[92] br[92] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_95 
+ bl[93] br[93] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_96 
+ bl[94] br[94] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_97 
+ bl[95] br[95] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_98 
+ bl[96] br[96] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_99 
+ bl[97] br[97] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_100 
+ bl[98] br[98] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_101 
+ bl[99] br[99] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_102 
+ bl[100] br[100] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_103 
+ bl[101] br[101] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_104 
+ bl[102] br[102] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_105 
+ bl[103] br[103] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_106 
+ bl[104] br[104] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_107 
+ bl[105] br[105] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_108 
+ bl[106] br[106] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_109 
+ bl[107] br[107] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_110 
+ bl[108] br[108] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_111 
+ bl[109] br[109] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_112 
+ bl[110] br[110] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_113 
+ bl[111] br[111] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_114 
+ bl[112] br[112] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_115 
+ bl[113] br[113] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_116 
+ bl[114] br[114] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_117 
+ bl[115] br[115] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_118 
+ bl[116] br[116] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_119 
+ bl[117] br[117] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_120 
+ bl[118] br[118] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_121 
+ bl[119] br[119] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_122 
+ bl[120] br[120] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_123 
+ bl[121] br[121] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_124 
+ bl[122] br[122] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_125 
+ bl[123] br[123] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_126 
+ bl[124] br[124] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_127 
+ bl[125] br[125] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_128 
+ bl[126] br[126] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_129 
+ bl[127] br[127] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_130 
+ bl[128] br[128] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_131 
+ bl[129] br[129] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_132 
+ bl[130] br[130] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_133 
+ bl[131] br[131] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_134 
+ bl[132] br[132] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_135 
+ bl[133] br[133] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_136 
+ bl[134] br[134] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_137 
+ bl[135] br[135] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_138 
+ bl[136] br[136] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_139 
+ bl[137] br[137] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_140 
+ bl[138] br[138] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_141 
+ bl[139] br[139] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_142 
+ bl[140] br[140] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_143 
+ bl[141] br[141] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_144 
+ bl[142] br[142] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_145 
+ bl[143] br[143] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_146 
+ bl[144] br[144] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_147 
+ bl[145] br[145] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_148 
+ bl[146] br[146] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_149 
+ bl[147] br[147] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_150 
+ bl[148] br[148] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_151 
+ bl[149] br[149] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_152 
+ bl[150] br[150] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_153 
+ bl[151] br[151] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_154 
+ bl[152] br[152] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_155 
+ bl[153] br[153] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_156 
+ bl[154] br[154] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_157 
+ bl[155] br[155] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_158 
+ bl[156] br[156] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_159 
+ bl[157] br[157] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_160 
+ bl[158] br[158] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_161 
+ bl[159] br[159] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_162 
+ bl[160] br[160] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_163 
+ bl[161] br[161] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_164 
+ bl[162] br[162] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_165 
+ bl[163] br[163] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_166 
+ bl[164] br[164] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_167 
+ bl[165] br[165] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_168 
+ bl[166] br[166] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_169 
+ bl[167] br[167] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_170 
+ bl[168] br[168] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_171 
+ bl[169] br[169] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_172 
+ bl[170] br[170] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_173 
+ bl[171] br[171] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_174 
+ bl[172] br[172] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_175 
+ bl[173] br[173] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_176 
+ bl[174] br[174] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_177 
+ bl[175] br[175] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_178 
+ bl[176] br[176] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_179 
+ bl[177] br[177] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_180 
+ bl[178] br[178] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_181 
+ bl[179] br[179] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_182 
+ bl[180] br[180] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_183 
+ bl[181] br[181] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_184 
+ bl[182] br[182] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_185 
+ bl[183] br[183] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_186 
+ bl[184] br[184] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_187 
+ bl[185] br[185] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_188 
+ bl[186] br[186] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_189 
+ bl[187] br[187] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_190 
+ bl[188] br[188] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_191 
+ bl[189] br[189] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_192 
+ bl[190] br[190] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_193 
+ bl[191] br[191] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_194 
+ bl[192] br[192] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_195 
+ bl[193] br[193] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_196 
+ bl[194] br[194] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_197 
+ bl[195] br[195] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_198 
+ bl[196] br[196] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_199 
+ bl[197] br[197] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_200 
+ bl[198] br[198] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_201 
+ bl[199] br[199] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_202 
+ bl[200] br[200] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_203 
+ bl[201] br[201] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_204 
+ bl[202] br[202] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_205 
+ bl[203] br[203] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_206 
+ bl[204] br[204] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_207 
+ bl[205] br[205] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_208 
+ bl[206] br[206] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_209 
+ bl[207] br[207] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_210 
+ bl[208] br[208] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_211 
+ bl[209] br[209] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_212 
+ bl[210] br[210] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_213 
+ bl[211] br[211] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_214 
+ bl[212] br[212] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_215 
+ bl[213] br[213] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_216 
+ bl[214] br[214] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_217 
+ bl[215] br[215] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_218 
+ bl[216] br[216] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_219 
+ bl[217] br[217] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_220 
+ bl[218] br[218] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_221 
+ bl[219] br[219] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_222 
+ bl[220] br[220] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_223 
+ bl[221] br[221] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_224 
+ bl[222] br[222] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_225 
+ bl[223] br[223] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_226 
+ bl[224] br[224] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_227 
+ bl[225] br[225] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_228 
+ bl[226] br[226] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_229 
+ bl[227] br[227] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_230 
+ bl[228] br[228] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_231 
+ bl[229] br[229] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_232 
+ bl[230] br[230] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_233 
+ bl[231] br[231] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_234 
+ bl[232] br[232] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_235 
+ bl[233] br[233] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_236 
+ bl[234] br[234] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_237 
+ bl[235] br[235] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_238 
+ bl[236] br[236] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_239 
+ bl[237] br[237] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_240 
+ bl[238] br[238] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_241 
+ bl[239] br[239] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_242 
+ bl[240] br[240] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_243 
+ bl[241] br[241] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_244 
+ bl[242] br[242] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_245 
+ bl[243] br[243] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_246 
+ bl[244] br[244] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_247 
+ bl[245] br[245] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_248 
+ bl[246] br[246] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_249 
+ bl[247] br[247] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_250 
+ bl[248] br[248] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_251 
+ bl[249] br[249] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_252 
+ bl[250] br[250] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_253 
+ bl[251] br[251] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_254 
+ bl[252] br[252] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_255 
+ bl[253] br[253] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_256 
+ bl[254] br[254] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_257 
+ bl[255] br[255] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_258 
+ vdd vdd vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_259 
+ vdd vdd vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_0 
+ vdd vdd vss vdd vpb vnb wl[127] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_129_1 
+ rbl rbr vss vdd vpb vnb wl[127] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_129_2 
+ bl[0] br[0] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_3 
+ bl[1] br[1] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_4 
+ bl[2] br[2] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_5 
+ bl[3] br[3] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_6 
+ bl[4] br[4] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_7 
+ bl[5] br[5] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_8 
+ bl[6] br[6] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_9 
+ bl[7] br[7] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_10 
+ bl[8] br[8] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_11 
+ bl[9] br[9] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_12 
+ bl[10] br[10] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_13 
+ bl[11] br[11] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_14 
+ bl[12] br[12] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_15 
+ bl[13] br[13] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_16 
+ bl[14] br[14] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_17 
+ bl[15] br[15] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_18 
+ bl[16] br[16] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_19 
+ bl[17] br[17] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_20 
+ bl[18] br[18] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_21 
+ bl[19] br[19] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_22 
+ bl[20] br[20] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_23 
+ bl[21] br[21] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_24 
+ bl[22] br[22] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_25 
+ bl[23] br[23] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_26 
+ bl[24] br[24] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_27 
+ bl[25] br[25] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_28 
+ bl[26] br[26] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_29 
+ bl[27] br[27] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_30 
+ bl[28] br[28] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_31 
+ bl[29] br[29] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_32 
+ bl[30] br[30] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_33 
+ bl[31] br[31] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_34 
+ bl[32] br[32] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_35 
+ bl[33] br[33] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_36 
+ bl[34] br[34] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_37 
+ bl[35] br[35] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_38 
+ bl[36] br[36] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_39 
+ bl[37] br[37] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_40 
+ bl[38] br[38] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_41 
+ bl[39] br[39] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_42 
+ bl[40] br[40] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_43 
+ bl[41] br[41] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_44 
+ bl[42] br[42] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_45 
+ bl[43] br[43] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_46 
+ bl[44] br[44] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_47 
+ bl[45] br[45] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_48 
+ bl[46] br[46] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_49 
+ bl[47] br[47] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_50 
+ bl[48] br[48] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_51 
+ bl[49] br[49] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_52 
+ bl[50] br[50] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_53 
+ bl[51] br[51] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_54 
+ bl[52] br[52] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_55 
+ bl[53] br[53] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_56 
+ bl[54] br[54] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_57 
+ bl[55] br[55] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_58 
+ bl[56] br[56] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_59 
+ bl[57] br[57] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_60 
+ bl[58] br[58] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_61 
+ bl[59] br[59] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_62 
+ bl[60] br[60] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_63 
+ bl[61] br[61] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_64 
+ bl[62] br[62] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_65 
+ bl[63] br[63] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_66 
+ bl[64] br[64] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_67 
+ bl[65] br[65] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_68 
+ bl[66] br[66] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_69 
+ bl[67] br[67] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_70 
+ bl[68] br[68] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_71 
+ bl[69] br[69] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_72 
+ bl[70] br[70] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_73 
+ bl[71] br[71] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_74 
+ bl[72] br[72] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_75 
+ bl[73] br[73] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_76 
+ bl[74] br[74] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_77 
+ bl[75] br[75] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_78 
+ bl[76] br[76] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_79 
+ bl[77] br[77] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_80 
+ bl[78] br[78] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_81 
+ bl[79] br[79] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_82 
+ bl[80] br[80] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_83 
+ bl[81] br[81] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_84 
+ bl[82] br[82] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_85 
+ bl[83] br[83] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_86 
+ bl[84] br[84] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_87 
+ bl[85] br[85] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_88 
+ bl[86] br[86] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_89 
+ bl[87] br[87] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_90 
+ bl[88] br[88] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_91 
+ bl[89] br[89] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_92 
+ bl[90] br[90] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_93 
+ bl[91] br[91] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_94 
+ bl[92] br[92] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_95 
+ bl[93] br[93] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_96 
+ bl[94] br[94] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_97 
+ bl[95] br[95] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_98 
+ bl[96] br[96] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_99 
+ bl[97] br[97] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_100 
+ bl[98] br[98] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_101 
+ bl[99] br[99] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_102 
+ bl[100] br[100] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_103 
+ bl[101] br[101] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_104 
+ bl[102] br[102] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_105 
+ bl[103] br[103] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_106 
+ bl[104] br[104] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_107 
+ bl[105] br[105] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_108 
+ bl[106] br[106] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_109 
+ bl[107] br[107] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_110 
+ bl[108] br[108] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_111 
+ bl[109] br[109] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_112 
+ bl[110] br[110] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_113 
+ bl[111] br[111] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_114 
+ bl[112] br[112] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_115 
+ bl[113] br[113] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_116 
+ bl[114] br[114] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_117 
+ bl[115] br[115] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_118 
+ bl[116] br[116] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_119 
+ bl[117] br[117] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_120 
+ bl[118] br[118] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_121 
+ bl[119] br[119] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_122 
+ bl[120] br[120] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_123 
+ bl[121] br[121] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_124 
+ bl[122] br[122] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_125 
+ bl[123] br[123] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_126 
+ bl[124] br[124] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_127 
+ bl[125] br[125] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_128 
+ bl[126] br[126] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_129 
+ bl[127] br[127] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_130 
+ bl[128] br[128] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_131 
+ bl[129] br[129] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_132 
+ bl[130] br[130] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_133 
+ bl[131] br[131] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_134 
+ bl[132] br[132] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_135 
+ bl[133] br[133] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_136 
+ bl[134] br[134] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_137 
+ bl[135] br[135] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_138 
+ bl[136] br[136] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_139 
+ bl[137] br[137] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_140 
+ bl[138] br[138] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_141 
+ bl[139] br[139] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_142 
+ bl[140] br[140] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_143 
+ bl[141] br[141] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_144 
+ bl[142] br[142] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_145 
+ bl[143] br[143] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_146 
+ bl[144] br[144] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_147 
+ bl[145] br[145] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_148 
+ bl[146] br[146] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_149 
+ bl[147] br[147] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_150 
+ bl[148] br[148] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_151 
+ bl[149] br[149] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_152 
+ bl[150] br[150] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_153 
+ bl[151] br[151] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_154 
+ bl[152] br[152] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_155 
+ bl[153] br[153] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_156 
+ bl[154] br[154] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_157 
+ bl[155] br[155] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_158 
+ bl[156] br[156] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_159 
+ bl[157] br[157] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_160 
+ bl[158] br[158] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_161 
+ bl[159] br[159] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_162 
+ bl[160] br[160] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_163 
+ bl[161] br[161] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_164 
+ bl[162] br[162] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_165 
+ bl[163] br[163] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_166 
+ bl[164] br[164] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_167 
+ bl[165] br[165] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_168 
+ bl[166] br[166] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_169 
+ bl[167] br[167] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_170 
+ bl[168] br[168] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_171 
+ bl[169] br[169] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_172 
+ bl[170] br[170] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_173 
+ bl[171] br[171] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_174 
+ bl[172] br[172] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_175 
+ bl[173] br[173] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_176 
+ bl[174] br[174] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_177 
+ bl[175] br[175] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_178 
+ bl[176] br[176] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_179 
+ bl[177] br[177] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_180 
+ bl[178] br[178] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_181 
+ bl[179] br[179] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_182 
+ bl[180] br[180] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_183 
+ bl[181] br[181] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_184 
+ bl[182] br[182] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_185 
+ bl[183] br[183] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_186 
+ bl[184] br[184] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_187 
+ bl[185] br[185] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_188 
+ bl[186] br[186] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_189 
+ bl[187] br[187] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_190 
+ bl[188] br[188] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_191 
+ bl[189] br[189] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_192 
+ bl[190] br[190] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_193 
+ bl[191] br[191] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_194 
+ bl[192] br[192] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_195 
+ bl[193] br[193] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_196 
+ bl[194] br[194] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_197 
+ bl[195] br[195] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_198 
+ bl[196] br[196] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_199 
+ bl[197] br[197] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_200 
+ bl[198] br[198] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_201 
+ bl[199] br[199] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_202 
+ bl[200] br[200] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_203 
+ bl[201] br[201] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_204 
+ bl[202] br[202] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_205 
+ bl[203] br[203] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_206 
+ bl[204] br[204] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_207 
+ bl[205] br[205] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_208 
+ bl[206] br[206] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_209 
+ bl[207] br[207] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_210 
+ bl[208] br[208] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_211 
+ bl[209] br[209] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_212 
+ bl[210] br[210] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_213 
+ bl[211] br[211] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_214 
+ bl[212] br[212] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_215 
+ bl[213] br[213] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_216 
+ bl[214] br[214] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_217 
+ bl[215] br[215] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_218 
+ bl[216] br[216] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_219 
+ bl[217] br[217] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_220 
+ bl[218] br[218] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_221 
+ bl[219] br[219] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_222 
+ bl[220] br[220] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_223 
+ bl[221] br[221] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_224 
+ bl[222] br[222] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_225 
+ bl[223] br[223] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_226 
+ bl[224] br[224] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_227 
+ bl[225] br[225] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_228 
+ bl[226] br[226] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_229 
+ bl[227] br[227] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_230 
+ bl[228] br[228] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_231 
+ bl[229] br[229] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_232 
+ bl[230] br[230] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_233 
+ bl[231] br[231] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_234 
+ bl[232] br[232] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_235 
+ bl[233] br[233] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_236 
+ bl[234] br[234] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_237 
+ bl[235] br[235] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_238 
+ bl[236] br[236] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_239 
+ bl[237] br[237] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_240 
+ bl[238] br[238] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_241 
+ bl[239] br[239] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_242 
+ bl[240] br[240] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_243 
+ bl[241] br[241] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_244 
+ bl[242] br[242] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_245 
+ bl[243] br[243] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_246 
+ bl[244] br[244] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_247 
+ bl[245] br[245] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_248 
+ bl[246] br[246] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_249 
+ bl[247] br[247] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_250 
+ bl[248] br[248] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_251 
+ bl[249] br[249] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_252 
+ bl[250] br[250] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_253 
+ bl[251] br[251] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_254 
+ bl[252] br[252] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_255 
+ bl[253] br[253] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_256 
+ bl[254] br[254] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_257 
+ bl[255] br[255] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_258 
+ vdd vdd vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_259 
+ vdd vdd vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_0 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_1 
+ rbl rbr vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_2 
+ bl[0] br[0] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_3 
+ bl[1] br[1] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_4 
+ bl[2] br[2] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_5 
+ bl[3] br[3] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_6 
+ bl[4] br[4] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_7 
+ bl[5] br[5] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_8 
+ bl[6] br[6] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_9 
+ bl[7] br[7] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_10 
+ bl[8] br[8] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_11 
+ bl[9] br[9] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_12 
+ bl[10] br[10] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_13 
+ bl[11] br[11] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_14 
+ bl[12] br[12] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_15 
+ bl[13] br[13] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_16 
+ bl[14] br[14] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_17 
+ bl[15] br[15] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_18 
+ bl[16] br[16] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_19 
+ bl[17] br[17] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_20 
+ bl[18] br[18] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_21 
+ bl[19] br[19] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_22 
+ bl[20] br[20] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_23 
+ bl[21] br[21] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_24 
+ bl[22] br[22] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_25 
+ bl[23] br[23] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_26 
+ bl[24] br[24] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_27 
+ bl[25] br[25] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_28 
+ bl[26] br[26] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_29 
+ bl[27] br[27] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_30 
+ bl[28] br[28] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_31 
+ bl[29] br[29] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_32 
+ bl[30] br[30] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_33 
+ bl[31] br[31] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_34 
+ bl[32] br[32] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_35 
+ bl[33] br[33] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_36 
+ bl[34] br[34] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_37 
+ bl[35] br[35] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_38 
+ bl[36] br[36] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_39 
+ bl[37] br[37] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_40 
+ bl[38] br[38] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_41 
+ bl[39] br[39] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_42 
+ bl[40] br[40] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_43 
+ bl[41] br[41] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_44 
+ bl[42] br[42] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_45 
+ bl[43] br[43] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_46 
+ bl[44] br[44] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_47 
+ bl[45] br[45] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_48 
+ bl[46] br[46] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_49 
+ bl[47] br[47] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_50 
+ bl[48] br[48] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_51 
+ bl[49] br[49] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_52 
+ bl[50] br[50] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_53 
+ bl[51] br[51] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_54 
+ bl[52] br[52] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_55 
+ bl[53] br[53] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_56 
+ bl[54] br[54] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_57 
+ bl[55] br[55] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_58 
+ bl[56] br[56] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_59 
+ bl[57] br[57] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_60 
+ bl[58] br[58] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_61 
+ bl[59] br[59] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_62 
+ bl[60] br[60] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_63 
+ bl[61] br[61] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_64 
+ bl[62] br[62] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_65 
+ bl[63] br[63] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_66 
+ bl[64] br[64] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_67 
+ bl[65] br[65] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_68 
+ bl[66] br[66] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_69 
+ bl[67] br[67] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_70 
+ bl[68] br[68] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_71 
+ bl[69] br[69] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_72 
+ bl[70] br[70] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_73 
+ bl[71] br[71] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_74 
+ bl[72] br[72] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_75 
+ bl[73] br[73] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_76 
+ bl[74] br[74] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_77 
+ bl[75] br[75] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_78 
+ bl[76] br[76] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_79 
+ bl[77] br[77] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_80 
+ bl[78] br[78] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_81 
+ bl[79] br[79] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_82 
+ bl[80] br[80] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_83 
+ bl[81] br[81] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_84 
+ bl[82] br[82] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_85 
+ bl[83] br[83] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_86 
+ bl[84] br[84] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_87 
+ bl[85] br[85] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_88 
+ bl[86] br[86] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_89 
+ bl[87] br[87] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_90 
+ bl[88] br[88] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_91 
+ bl[89] br[89] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_92 
+ bl[90] br[90] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_93 
+ bl[91] br[91] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_94 
+ bl[92] br[92] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_95 
+ bl[93] br[93] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_96 
+ bl[94] br[94] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_97 
+ bl[95] br[95] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_98 
+ bl[96] br[96] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_99 
+ bl[97] br[97] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_100 
+ bl[98] br[98] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_101 
+ bl[99] br[99] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_102 
+ bl[100] br[100] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_103 
+ bl[101] br[101] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_104 
+ bl[102] br[102] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_105 
+ bl[103] br[103] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_106 
+ bl[104] br[104] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_107 
+ bl[105] br[105] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_108 
+ bl[106] br[106] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_109 
+ bl[107] br[107] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_110 
+ bl[108] br[108] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_111 
+ bl[109] br[109] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_112 
+ bl[110] br[110] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_113 
+ bl[111] br[111] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_114 
+ bl[112] br[112] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_115 
+ bl[113] br[113] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_116 
+ bl[114] br[114] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_117 
+ bl[115] br[115] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_118 
+ bl[116] br[116] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_119 
+ bl[117] br[117] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_120 
+ bl[118] br[118] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_121 
+ bl[119] br[119] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_122 
+ bl[120] br[120] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_123 
+ bl[121] br[121] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_124 
+ bl[122] br[122] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_125 
+ bl[123] br[123] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_126 
+ bl[124] br[124] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_127 
+ bl[125] br[125] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_128 
+ bl[126] br[126] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_129 
+ bl[127] br[127] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_130 
+ bl[128] br[128] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_131 
+ bl[129] br[129] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_132 
+ bl[130] br[130] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_133 
+ bl[131] br[131] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_134 
+ bl[132] br[132] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_135 
+ bl[133] br[133] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_136 
+ bl[134] br[134] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_137 
+ bl[135] br[135] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_138 
+ bl[136] br[136] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_139 
+ bl[137] br[137] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_140 
+ bl[138] br[138] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_141 
+ bl[139] br[139] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_142 
+ bl[140] br[140] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_143 
+ bl[141] br[141] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_144 
+ bl[142] br[142] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_145 
+ bl[143] br[143] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_146 
+ bl[144] br[144] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_147 
+ bl[145] br[145] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_148 
+ bl[146] br[146] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_149 
+ bl[147] br[147] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_150 
+ bl[148] br[148] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_151 
+ bl[149] br[149] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_152 
+ bl[150] br[150] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_153 
+ bl[151] br[151] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_154 
+ bl[152] br[152] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_155 
+ bl[153] br[153] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_156 
+ bl[154] br[154] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_157 
+ bl[155] br[155] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_158 
+ bl[156] br[156] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_159 
+ bl[157] br[157] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_160 
+ bl[158] br[158] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_161 
+ bl[159] br[159] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_162 
+ bl[160] br[160] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_163 
+ bl[161] br[161] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_164 
+ bl[162] br[162] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_165 
+ bl[163] br[163] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_166 
+ bl[164] br[164] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_167 
+ bl[165] br[165] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_168 
+ bl[166] br[166] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_169 
+ bl[167] br[167] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_170 
+ bl[168] br[168] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_171 
+ bl[169] br[169] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_172 
+ bl[170] br[170] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_173 
+ bl[171] br[171] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_174 
+ bl[172] br[172] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_175 
+ bl[173] br[173] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_176 
+ bl[174] br[174] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_177 
+ bl[175] br[175] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_178 
+ bl[176] br[176] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_179 
+ bl[177] br[177] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_180 
+ bl[178] br[178] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_181 
+ bl[179] br[179] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_182 
+ bl[180] br[180] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_183 
+ bl[181] br[181] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_184 
+ bl[182] br[182] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_185 
+ bl[183] br[183] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_186 
+ bl[184] br[184] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_187 
+ bl[185] br[185] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_188 
+ bl[186] br[186] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_189 
+ bl[187] br[187] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_190 
+ bl[188] br[188] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_191 
+ bl[189] br[189] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_192 
+ bl[190] br[190] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_193 
+ bl[191] br[191] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_194 
+ bl[192] br[192] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_195 
+ bl[193] br[193] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_196 
+ bl[194] br[194] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_197 
+ bl[195] br[195] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_198 
+ bl[196] br[196] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_199 
+ bl[197] br[197] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_200 
+ bl[198] br[198] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_201 
+ bl[199] br[199] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_202 
+ bl[200] br[200] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_203 
+ bl[201] br[201] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_204 
+ bl[202] br[202] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_205 
+ bl[203] br[203] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_206 
+ bl[204] br[204] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_207 
+ bl[205] br[205] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_208 
+ bl[206] br[206] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_209 
+ bl[207] br[207] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_210 
+ bl[208] br[208] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_211 
+ bl[209] br[209] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_212 
+ bl[210] br[210] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_213 
+ bl[211] br[211] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_214 
+ bl[212] br[212] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_215 
+ bl[213] br[213] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_216 
+ bl[214] br[214] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_217 
+ bl[215] br[215] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_218 
+ bl[216] br[216] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_219 
+ bl[217] br[217] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_220 
+ bl[218] br[218] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_221 
+ bl[219] br[219] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_222 
+ bl[220] br[220] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_223 
+ bl[221] br[221] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_224 
+ bl[222] br[222] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_225 
+ bl[223] br[223] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_226 
+ bl[224] br[224] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_227 
+ bl[225] br[225] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_228 
+ bl[226] br[226] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_229 
+ bl[227] br[227] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_230 
+ bl[228] br[228] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_231 
+ bl[229] br[229] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_232 
+ bl[230] br[230] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_233 
+ bl[231] br[231] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_234 
+ bl[232] br[232] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_235 
+ bl[233] br[233] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_236 
+ bl[234] br[234] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_237 
+ bl[235] br[235] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_238 
+ bl[236] br[236] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_239 
+ bl[237] br[237] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_240 
+ bl[238] br[238] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_241 
+ bl[239] br[239] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_242 
+ bl[240] br[240] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_243 
+ bl[241] br[241] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_244 
+ bl[242] br[242] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_245 
+ bl[243] br[243] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_246 
+ bl[244] br[244] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_247 
+ bl[245] br[245] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_248 
+ bl[246] br[246] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_249 
+ bl[247] br[247] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_250 
+ bl[248] br[248] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_251 
+ bl[249] br[249] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_252 
+ bl[250] br[250] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_253 
+ bl[251] br[251] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_254 
+ bl[252] br[252] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_255 
+ bl[253] br[253] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_256 
+ bl[254] br[254] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_257 
+ bl[255] br[255] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_258 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_259 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_0 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_1 
+ rbl rbr vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_2 
+ bl[0] br[0] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_3 
+ bl[1] br[1] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_4 
+ bl[2] br[2] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_5 
+ bl[3] br[3] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_6 
+ bl[4] br[4] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_7 
+ bl[5] br[5] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_8 
+ bl[6] br[6] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_9 
+ bl[7] br[7] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_10 
+ bl[8] br[8] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_11 
+ bl[9] br[9] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_12 
+ bl[10] br[10] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_13 
+ bl[11] br[11] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_14 
+ bl[12] br[12] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_15 
+ bl[13] br[13] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_16 
+ bl[14] br[14] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_17 
+ bl[15] br[15] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_18 
+ bl[16] br[16] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_19 
+ bl[17] br[17] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_20 
+ bl[18] br[18] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_21 
+ bl[19] br[19] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_22 
+ bl[20] br[20] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_23 
+ bl[21] br[21] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_24 
+ bl[22] br[22] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_25 
+ bl[23] br[23] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_26 
+ bl[24] br[24] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_27 
+ bl[25] br[25] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_28 
+ bl[26] br[26] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_29 
+ bl[27] br[27] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_30 
+ bl[28] br[28] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_31 
+ bl[29] br[29] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_32 
+ bl[30] br[30] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_33 
+ bl[31] br[31] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_34 
+ bl[32] br[32] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_35 
+ bl[33] br[33] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_36 
+ bl[34] br[34] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_37 
+ bl[35] br[35] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_38 
+ bl[36] br[36] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_39 
+ bl[37] br[37] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_40 
+ bl[38] br[38] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_41 
+ bl[39] br[39] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_42 
+ bl[40] br[40] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_43 
+ bl[41] br[41] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_44 
+ bl[42] br[42] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_45 
+ bl[43] br[43] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_46 
+ bl[44] br[44] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_47 
+ bl[45] br[45] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_48 
+ bl[46] br[46] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_49 
+ bl[47] br[47] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_50 
+ bl[48] br[48] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_51 
+ bl[49] br[49] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_52 
+ bl[50] br[50] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_53 
+ bl[51] br[51] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_54 
+ bl[52] br[52] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_55 
+ bl[53] br[53] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_56 
+ bl[54] br[54] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_57 
+ bl[55] br[55] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_58 
+ bl[56] br[56] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_59 
+ bl[57] br[57] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_60 
+ bl[58] br[58] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_61 
+ bl[59] br[59] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_62 
+ bl[60] br[60] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_63 
+ bl[61] br[61] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_64 
+ bl[62] br[62] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_65 
+ bl[63] br[63] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_66 
+ bl[64] br[64] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_67 
+ bl[65] br[65] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_68 
+ bl[66] br[66] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_69 
+ bl[67] br[67] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_70 
+ bl[68] br[68] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_71 
+ bl[69] br[69] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_72 
+ bl[70] br[70] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_73 
+ bl[71] br[71] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_74 
+ bl[72] br[72] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_75 
+ bl[73] br[73] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_76 
+ bl[74] br[74] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_77 
+ bl[75] br[75] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_78 
+ bl[76] br[76] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_79 
+ bl[77] br[77] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_80 
+ bl[78] br[78] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_81 
+ bl[79] br[79] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_82 
+ bl[80] br[80] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_83 
+ bl[81] br[81] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_84 
+ bl[82] br[82] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_85 
+ bl[83] br[83] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_86 
+ bl[84] br[84] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_87 
+ bl[85] br[85] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_88 
+ bl[86] br[86] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_89 
+ bl[87] br[87] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_90 
+ bl[88] br[88] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_91 
+ bl[89] br[89] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_92 
+ bl[90] br[90] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_93 
+ bl[91] br[91] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_94 
+ bl[92] br[92] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_95 
+ bl[93] br[93] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_96 
+ bl[94] br[94] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_97 
+ bl[95] br[95] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_98 
+ bl[96] br[96] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_99 
+ bl[97] br[97] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_100 
+ bl[98] br[98] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_101 
+ bl[99] br[99] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_102 
+ bl[100] br[100] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_103 
+ bl[101] br[101] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_104 
+ bl[102] br[102] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_105 
+ bl[103] br[103] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_106 
+ bl[104] br[104] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_107 
+ bl[105] br[105] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_108 
+ bl[106] br[106] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_109 
+ bl[107] br[107] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_110 
+ bl[108] br[108] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_111 
+ bl[109] br[109] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_112 
+ bl[110] br[110] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_113 
+ bl[111] br[111] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_114 
+ bl[112] br[112] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_115 
+ bl[113] br[113] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_116 
+ bl[114] br[114] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_117 
+ bl[115] br[115] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_118 
+ bl[116] br[116] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_119 
+ bl[117] br[117] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_120 
+ bl[118] br[118] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_121 
+ bl[119] br[119] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_122 
+ bl[120] br[120] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_123 
+ bl[121] br[121] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_124 
+ bl[122] br[122] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_125 
+ bl[123] br[123] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_126 
+ bl[124] br[124] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_127 
+ bl[125] br[125] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_128 
+ bl[126] br[126] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_129 
+ bl[127] br[127] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_130 
+ bl[128] br[128] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_131 
+ bl[129] br[129] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_132 
+ bl[130] br[130] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_133 
+ bl[131] br[131] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_134 
+ bl[132] br[132] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_135 
+ bl[133] br[133] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_136 
+ bl[134] br[134] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_137 
+ bl[135] br[135] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_138 
+ bl[136] br[136] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_139 
+ bl[137] br[137] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_140 
+ bl[138] br[138] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_141 
+ bl[139] br[139] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_142 
+ bl[140] br[140] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_143 
+ bl[141] br[141] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_144 
+ bl[142] br[142] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_145 
+ bl[143] br[143] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_146 
+ bl[144] br[144] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_147 
+ bl[145] br[145] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_148 
+ bl[146] br[146] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_149 
+ bl[147] br[147] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_150 
+ bl[148] br[148] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_151 
+ bl[149] br[149] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_152 
+ bl[150] br[150] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_153 
+ bl[151] br[151] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_154 
+ bl[152] br[152] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_155 
+ bl[153] br[153] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_156 
+ bl[154] br[154] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_157 
+ bl[155] br[155] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_158 
+ bl[156] br[156] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_159 
+ bl[157] br[157] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_160 
+ bl[158] br[158] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_161 
+ bl[159] br[159] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_162 
+ bl[160] br[160] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_163 
+ bl[161] br[161] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_164 
+ bl[162] br[162] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_165 
+ bl[163] br[163] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_166 
+ bl[164] br[164] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_167 
+ bl[165] br[165] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_168 
+ bl[166] br[166] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_169 
+ bl[167] br[167] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_170 
+ bl[168] br[168] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_171 
+ bl[169] br[169] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_172 
+ bl[170] br[170] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_173 
+ bl[171] br[171] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_174 
+ bl[172] br[172] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_175 
+ bl[173] br[173] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_176 
+ bl[174] br[174] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_177 
+ bl[175] br[175] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_178 
+ bl[176] br[176] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_179 
+ bl[177] br[177] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_180 
+ bl[178] br[178] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_181 
+ bl[179] br[179] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_182 
+ bl[180] br[180] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_183 
+ bl[181] br[181] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_184 
+ bl[182] br[182] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_185 
+ bl[183] br[183] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_186 
+ bl[184] br[184] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_187 
+ bl[185] br[185] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_188 
+ bl[186] br[186] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_189 
+ bl[187] br[187] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_190 
+ bl[188] br[188] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_191 
+ bl[189] br[189] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_192 
+ bl[190] br[190] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_193 
+ bl[191] br[191] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_194 
+ bl[192] br[192] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_195 
+ bl[193] br[193] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_196 
+ bl[194] br[194] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_197 
+ bl[195] br[195] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_198 
+ bl[196] br[196] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_199 
+ bl[197] br[197] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_200 
+ bl[198] br[198] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_201 
+ bl[199] br[199] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_202 
+ bl[200] br[200] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_203 
+ bl[201] br[201] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_204 
+ bl[202] br[202] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_205 
+ bl[203] br[203] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_206 
+ bl[204] br[204] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_207 
+ bl[205] br[205] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_208 
+ bl[206] br[206] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_209 
+ bl[207] br[207] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_210 
+ bl[208] br[208] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_211 
+ bl[209] br[209] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_212 
+ bl[210] br[210] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_213 
+ bl[211] br[211] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_214 
+ bl[212] br[212] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_215 
+ bl[213] br[213] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_216 
+ bl[214] br[214] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_217 
+ bl[215] br[215] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_218 
+ bl[216] br[216] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_219 
+ bl[217] br[217] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_220 
+ bl[218] br[218] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_221 
+ bl[219] br[219] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_222 
+ bl[220] br[220] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_223 
+ bl[221] br[221] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_224 
+ bl[222] br[222] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_225 
+ bl[223] br[223] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_226 
+ bl[224] br[224] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_227 
+ bl[225] br[225] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_228 
+ bl[226] br[226] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_229 
+ bl[227] br[227] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_230 
+ bl[228] br[228] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_231 
+ bl[229] br[229] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_232 
+ bl[230] br[230] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_233 
+ bl[231] br[231] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_234 
+ bl[232] br[232] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_235 
+ bl[233] br[233] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_236 
+ bl[234] br[234] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_237 
+ bl[235] br[235] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_238 
+ bl[236] br[236] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_239 
+ bl[237] br[237] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_240 
+ bl[238] br[238] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_241 
+ bl[239] br[239] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_242 
+ bl[240] br[240] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_243 
+ bl[241] br[241] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_244 
+ bl[242] br[242] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_245 
+ bl[243] br[243] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_246 
+ bl[244] br[244] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_247 
+ bl[245] br[245] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_248 
+ bl[246] br[246] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_249 
+ bl[247] br[247] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_250 
+ bl[248] br[248] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_251 
+ bl[249] br[249] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_252 
+ bl[250] br[250] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_253 
+ bl[251] br[251] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_254 
+ bl[252] br[252] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_255 
+ bl[253] br[253] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_256 
+ bl[254] br[254] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_257 
+ bl[255] br[255] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_258 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_259 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xcolend_0_bot 
+ vdd vdd vss vdd vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_0_top 
+ vdd vdd vss vdd vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_1_bot 
+ rbr vdd vss rbl vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_1_top 
+ rbr vdd vss rbl vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_2_bot 
+ br[0] vdd vss bl[0] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_2_top 
+ br[0] vdd vss bl[0] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_3_bot 
+ br[1] vdd vss bl[1] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_3_top 
+ br[1] vdd vss bl[1] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_4_bot 
+ br[2] vdd vss bl[2] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_4_top 
+ br[2] vdd vss bl[2] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_5_bot 
+ br[3] vdd vss bl[3] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_5_top 
+ br[3] vdd vss bl[3] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_6_bot 
+ br[4] vdd vss bl[4] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_6_top 
+ br[4] vdd vss bl[4] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_7_bot 
+ br[5] vdd vss bl[5] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_7_top 
+ br[5] vdd vss bl[5] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_8_bot 
+ br[6] vdd vss bl[6] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_8_top 
+ br[6] vdd vss bl[6] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_9_bot 
+ br[7] vdd vss bl[7] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_9_top 
+ br[7] vdd vss bl[7] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_10_bot 
+ br[8] vdd vss bl[8] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_10_top 
+ br[8] vdd vss bl[8] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_11_bot 
+ br[9] vdd vss bl[9] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_11_top 
+ br[9] vdd vss bl[9] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_12_bot 
+ br[10] vdd vss bl[10] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_12_top 
+ br[10] vdd vss bl[10] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_13_bot 
+ br[11] vdd vss bl[11] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_13_top 
+ br[11] vdd vss bl[11] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_14_bot 
+ br[12] vdd vss bl[12] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_14_top 
+ br[12] vdd vss bl[12] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_15_bot 
+ br[13] vdd vss bl[13] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_15_top 
+ br[13] vdd vss bl[13] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_16_bot 
+ br[14] vdd vss bl[14] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_16_top 
+ br[14] vdd vss bl[14] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_17_bot 
+ br[15] vdd vss bl[15] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_17_top 
+ br[15] vdd vss bl[15] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_18_bot 
+ br[16] vdd vss bl[16] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_18_top 
+ br[16] vdd vss bl[16] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_19_bot 
+ br[17] vdd vss bl[17] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_19_top 
+ br[17] vdd vss bl[17] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_20_bot 
+ br[18] vdd vss bl[18] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_20_top 
+ br[18] vdd vss bl[18] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_21_bot 
+ br[19] vdd vss bl[19] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_21_top 
+ br[19] vdd vss bl[19] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_22_bot 
+ br[20] vdd vss bl[20] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_22_top 
+ br[20] vdd vss bl[20] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_23_bot 
+ br[21] vdd vss bl[21] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_23_top 
+ br[21] vdd vss bl[21] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_24_bot 
+ br[22] vdd vss bl[22] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_24_top 
+ br[22] vdd vss bl[22] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_25_bot 
+ br[23] vdd vss bl[23] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_25_top 
+ br[23] vdd vss bl[23] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_26_bot 
+ br[24] vdd vss bl[24] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_26_top 
+ br[24] vdd vss bl[24] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_27_bot 
+ br[25] vdd vss bl[25] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_27_top 
+ br[25] vdd vss bl[25] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_28_bot 
+ br[26] vdd vss bl[26] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_28_top 
+ br[26] vdd vss bl[26] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_29_bot 
+ br[27] vdd vss bl[27] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_29_top 
+ br[27] vdd vss bl[27] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_30_bot 
+ br[28] vdd vss bl[28] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_30_top 
+ br[28] vdd vss bl[28] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_31_bot 
+ br[29] vdd vss bl[29] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_31_top 
+ br[29] vdd vss bl[29] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_32_bot 
+ br[30] vdd vss bl[30] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_32_top 
+ br[30] vdd vss bl[30] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_33_bot 
+ br[31] vdd vss bl[31] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_33_top 
+ br[31] vdd vss bl[31] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_34_bot 
+ br[32] vdd vss bl[32] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_34_top 
+ br[32] vdd vss bl[32] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_35_bot 
+ br[33] vdd vss bl[33] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_35_top 
+ br[33] vdd vss bl[33] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_36_bot 
+ br[34] vdd vss bl[34] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_36_top 
+ br[34] vdd vss bl[34] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_37_bot 
+ br[35] vdd vss bl[35] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_37_top 
+ br[35] vdd vss bl[35] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_38_bot 
+ br[36] vdd vss bl[36] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_38_top 
+ br[36] vdd vss bl[36] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_39_bot 
+ br[37] vdd vss bl[37] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_39_top 
+ br[37] vdd vss bl[37] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_40_bot 
+ br[38] vdd vss bl[38] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_40_top 
+ br[38] vdd vss bl[38] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_41_bot 
+ br[39] vdd vss bl[39] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_41_top 
+ br[39] vdd vss bl[39] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_42_bot 
+ br[40] vdd vss bl[40] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_42_top 
+ br[40] vdd vss bl[40] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_43_bot 
+ br[41] vdd vss bl[41] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_43_top 
+ br[41] vdd vss bl[41] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_44_bot 
+ br[42] vdd vss bl[42] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_44_top 
+ br[42] vdd vss bl[42] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_45_bot 
+ br[43] vdd vss bl[43] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_45_top 
+ br[43] vdd vss bl[43] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_46_bot 
+ br[44] vdd vss bl[44] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_46_top 
+ br[44] vdd vss bl[44] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_47_bot 
+ br[45] vdd vss bl[45] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_47_top 
+ br[45] vdd vss bl[45] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_48_bot 
+ br[46] vdd vss bl[46] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_48_top 
+ br[46] vdd vss bl[46] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_49_bot 
+ br[47] vdd vss bl[47] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_49_top 
+ br[47] vdd vss bl[47] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_50_bot 
+ br[48] vdd vss bl[48] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_50_top 
+ br[48] vdd vss bl[48] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_51_bot 
+ br[49] vdd vss bl[49] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_51_top 
+ br[49] vdd vss bl[49] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_52_bot 
+ br[50] vdd vss bl[50] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_52_top 
+ br[50] vdd vss bl[50] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_53_bot 
+ br[51] vdd vss bl[51] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_53_top 
+ br[51] vdd vss bl[51] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_54_bot 
+ br[52] vdd vss bl[52] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_54_top 
+ br[52] vdd vss bl[52] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_55_bot 
+ br[53] vdd vss bl[53] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_55_top 
+ br[53] vdd vss bl[53] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_56_bot 
+ br[54] vdd vss bl[54] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_56_top 
+ br[54] vdd vss bl[54] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_57_bot 
+ br[55] vdd vss bl[55] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_57_top 
+ br[55] vdd vss bl[55] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_58_bot 
+ br[56] vdd vss bl[56] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_58_top 
+ br[56] vdd vss bl[56] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_59_bot 
+ br[57] vdd vss bl[57] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_59_top 
+ br[57] vdd vss bl[57] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_60_bot 
+ br[58] vdd vss bl[58] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_60_top 
+ br[58] vdd vss bl[58] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_61_bot 
+ br[59] vdd vss bl[59] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_61_top 
+ br[59] vdd vss bl[59] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_62_bot 
+ br[60] vdd vss bl[60] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_62_top 
+ br[60] vdd vss bl[60] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_63_bot 
+ br[61] vdd vss bl[61] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_63_top 
+ br[61] vdd vss bl[61] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_64_bot 
+ br[62] vdd vss bl[62] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_64_top 
+ br[62] vdd vss bl[62] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_65_bot 
+ br[63] vdd vss bl[63] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_65_top 
+ br[63] vdd vss bl[63] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_66_bot 
+ br[64] vdd vss bl[64] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_66_top 
+ br[64] vdd vss bl[64] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_67_bot 
+ br[65] vdd vss bl[65] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_67_top 
+ br[65] vdd vss bl[65] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_68_bot 
+ br[66] vdd vss bl[66] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_68_top 
+ br[66] vdd vss bl[66] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_69_bot 
+ br[67] vdd vss bl[67] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_69_top 
+ br[67] vdd vss bl[67] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_70_bot 
+ br[68] vdd vss bl[68] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_70_top 
+ br[68] vdd vss bl[68] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_71_bot 
+ br[69] vdd vss bl[69] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_71_top 
+ br[69] vdd vss bl[69] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_72_bot 
+ br[70] vdd vss bl[70] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_72_top 
+ br[70] vdd vss bl[70] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_73_bot 
+ br[71] vdd vss bl[71] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_73_top 
+ br[71] vdd vss bl[71] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_74_bot 
+ br[72] vdd vss bl[72] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_74_top 
+ br[72] vdd vss bl[72] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_75_bot 
+ br[73] vdd vss bl[73] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_75_top 
+ br[73] vdd vss bl[73] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_76_bot 
+ br[74] vdd vss bl[74] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_76_top 
+ br[74] vdd vss bl[74] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_77_bot 
+ br[75] vdd vss bl[75] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_77_top 
+ br[75] vdd vss bl[75] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_78_bot 
+ br[76] vdd vss bl[76] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_78_top 
+ br[76] vdd vss bl[76] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_79_bot 
+ br[77] vdd vss bl[77] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_79_top 
+ br[77] vdd vss bl[77] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_80_bot 
+ br[78] vdd vss bl[78] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_80_top 
+ br[78] vdd vss bl[78] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_81_bot 
+ br[79] vdd vss bl[79] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_81_top 
+ br[79] vdd vss bl[79] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_82_bot 
+ br[80] vdd vss bl[80] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_82_top 
+ br[80] vdd vss bl[80] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_83_bot 
+ br[81] vdd vss bl[81] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_83_top 
+ br[81] vdd vss bl[81] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_84_bot 
+ br[82] vdd vss bl[82] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_84_top 
+ br[82] vdd vss bl[82] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_85_bot 
+ br[83] vdd vss bl[83] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_85_top 
+ br[83] vdd vss bl[83] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_86_bot 
+ br[84] vdd vss bl[84] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_86_top 
+ br[84] vdd vss bl[84] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_87_bot 
+ br[85] vdd vss bl[85] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_87_top 
+ br[85] vdd vss bl[85] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_88_bot 
+ br[86] vdd vss bl[86] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_88_top 
+ br[86] vdd vss bl[86] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_89_bot 
+ br[87] vdd vss bl[87] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_89_top 
+ br[87] vdd vss bl[87] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_90_bot 
+ br[88] vdd vss bl[88] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_90_top 
+ br[88] vdd vss bl[88] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_91_bot 
+ br[89] vdd vss bl[89] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_91_top 
+ br[89] vdd vss bl[89] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_92_bot 
+ br[90] vdd vss bl[90] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_92_top 
+ br[90] vdd vss bl[90] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_93_bot 
+ br[91] vdd vss bl[91] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_93_top 
+ br[91] vdd vss bl[91] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_94_bot 
+ br[92] vdd vss bl[92] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_94_top 
+ br[92] vdd vss bl[92] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_95_bot 
+ br[93] vdd vss bl[93] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_95_top 
+ br[93] vdd vss bl[93] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_96_bot 
+ br[94] vdd vss bl[94] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_96_top 
+ br[94] vdd vss bl[94] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_97_bot 
+ br[95] vdd vss bl[95] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_97_top 
+ br[95] vdd vss bl[95] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_98_bot 
+ br[96] vdd vss bl[96] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_98_top 
+ br[96] vdd vss bl[96] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_99_bot 
+ br[97] vdd vss bl[97] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_99_top 
+ br[97] vdd vss bl[97] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_100_bot 
+ br[98] vdd vss bl[98] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_100_top 
+ br[98] vdd vss bl[98] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_101_bot 
+ br[99] vdd vss bl[99] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_101_top 
+ br[99] vdd vss bl[99] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_102_bot 
+ br[100] vdd vss bl[100] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_102_top 
+ br[100] vdd vss bl[100] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_103_bot 
+ br[101] vdd vss bl[101] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_103_top 
+ br[101] vdd vss bl[101] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_104_bot 
+ br[102] vdd vss bl[102] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_104_top 
+ br[102] vdd vss bl[102] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_105_bot 
+ br[103] vdd vss bl[103] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_105_top 
+ br[103] vdd vss bl[103] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_106_bot 
+ br[104] vdd vss bl[104] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_106_top 
+ br[104] vdd vss bl[104] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_107_bot 
+ br[105] vdd vss bl[105] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_107_top 
+ br[105] vdd vss bl[105] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_108_bot 
+ br[106] vdd vss bl[106] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_108_top 
+ br[106] vdd vss bl[106] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_109_bot 
+ br[107] vdd vss bl[107] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_109_top 
+ br[107] vdd vss bl[107] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_110_bot 
+ br[108] vdd vss bl[108] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_110_top 
+ br[108] vdd vss bl[108] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_111_bot 
+ br[109] vdd vss bl[109] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_111_top 
+ br[109] vdd vss bl[109] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_112_bot 
+ br[110] vdd vss bl[110] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_112_top 
+ br[110] vdd vss bl[110] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_113_bot 
+ br[111] vdd vss bl[111] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_113_top 
+ br[111] vdd vss bl[111] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_114_bot 
+ br[112] vdd vss bl[112] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_114_top 
+ br[112] vdd vss bl[112] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_115_bot 
+ br[113] vdd vss bl[113] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_115_top 
+ br[113] vdd vss bl[113] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_116_bot 
+ br[114] vdd vss bl[114] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_116_top 
+ br[114] vdd vss bl[114] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_117_bot 
+ br[115] vdd vss bl[115] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_117_top 
+ br[115] vdd vss bl[115] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_118_bot 
+ br[116] vdd vss bl[116] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_118_top 
+ br[116] vdd vss bl[116] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_119_bot 
+ br[117] vdd vss bl[117] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_119_top 
+ br[117] vdd vss bl[117] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_120_bot 
+ br[118] vdd vss bl[118] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_120_top 
+ br[118] vdd vss bl[118] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_121_bot 
+ br[119] vdd vss bl[119] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_121_top 
+ br[119] vdd vss bl[119] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_122_bot 
+ br[120] vdd vss bl[120] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_122_top 
+ br[120] vdd vss bl[120] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_123_bot 
+ br[121] vdd vss bl[121] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_123_top 
+ br[121] vdd vss bl[121] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_124_bot 
+ br[122] vdd vss bl[122] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_124_top 
+ br[122] vdd vss bl[122] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_125_bot 
+ br[123] vdd vss bl[123] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_125_top 
+ br[123] vdd vss bl[123] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_126_bot 
+ br[124] vdd vss bl[124] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_126_top 
+ br[124] vdd vss bl[124] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_127_bot 
+ br[125] vdd vss bl[125] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_127_top 
+ br[125] vdd vss bl[125] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_128_bot 
+ br[126] vdd vss bl[126] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_128_top 
+ br[126] vdd vss bl[126] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_129_bot 
+ br[127] vdd vss bl[127] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_129_top 
+ br[127] vdd vss bl[127] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_130_bot 
+ br[128] vdd vss bl[128] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_130_top 
+ br[128] vdd vss bl[128] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_131_bot 
+ br[129] vdd vss bl[129] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_131_top 
+ br[129] vdd vss bl[129] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_132_bot 
+ br[130] vdd vss bl[130] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_132_top 
+ br[130] vdd vss bl[130] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_133_bot 
+ br[131] vdd vss bl[131] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_133_top 
+ br[131] vdd vss bl[131] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_134_bot 
+ br[132] vdd vss bl[132] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_134_top 
+ br[132] vdd vss bl[132] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_135_bot 
+ br[133] vdd vss bl[133] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_135_top 
+ br[133] vdd vss bl[133] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_136_bot 
+ br[134] vdd vss bl[134] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_136_top 
+ br[134] vdd vss bl[134] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_137_bot 
+ br[135] vdd vss bl[135] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_137_top 
+ br[135] vdd vss bl[135] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_138_bot 
+ br[136] vdd vss bl[136] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_138_top 
+ br[136] vdd vss bl[136] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_139_bot 
+ br[137] vdd vss bl[137] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_139_top 
+ br[137] vdd vss bl[137] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_140_bot 
+ br[138] vdd vss bl[138] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_140_top 
+ br[138] vdd vss bl[138] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_141_bot 
+ br[139] vdd vss bl[139] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_141_top 
+ br[139] vdd vss bl[139] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_142_bot 
+ br[140] vdd vss bl[140] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_142_top 
+ br[140] vdd vss bl[140] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_143_bot 
+ br[141] vdd vss bl[141] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_143_top 
+ br[141] vdd vss bl[141] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_144_bot 
+ br[142] vdd vss bl[142] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_144_top 
+ br[142] vdd vss bl[142] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_145_bot 
+ br[143] vdd vss bl[143] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_145_top 
+ br[143] vdd vss bl[143] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_146_bot 
+ br[144] vdd vss bl[144] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_146_top 
+ br[144] vdd vss bl[144] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_147_bot 
+ br[145] vdd vss bl[145] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_147_top 
+ br[145] vdd vss bl[145] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_148_bot 
+ br[146] vdd vss bl[146] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_148_top 
+ br[146] vdd vss bl[146] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_149_bot 
+ br[147] vdd vss bl[147] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_149_top 
+ br[147] vdd vss bl[147] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_150_bot 
+ br[148] vdd vss bl[148] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_150_top 
+ br[148] vdd vss bl[148] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_151_bot 
+ br[149] vdd vss bl[149] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_151_top 
+ br[149] vdd vss bl[149] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_152_bot 
+ br[150] vdd vss bl[150] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_152_top 
+ br[150] vdd vss bl[150] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_153_bot 
+ br[151] vdd vss bl[151] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_153_top 
+ br[151] vdd vss bl[151] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_154_bot 
+ br[152] vdd vss bl[152] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_154_top 
+ br[152] vdd vss bl[152] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_155_bot 
+ br[153] vdd vss bl[153] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_155_top 
+ br[153] vdd vss bl[153] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_156_bot 
+ br[154] vdd vss bl[154] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_156_top 
+ br[154] vdd vss bl[154] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_157_bot 
+ br[155] vdd vss bl[155] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_157_top 
+ br[155] vdd vss bl[155] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_158_bot 
+ br[156] vdd vss bl[156] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_158_top 
+ br[156] vdd vss bl[156] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_159_bot 
+ br[157] vdd vss bl[157] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_159_top 
+ br[157] vdd vss bl[157] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_160_bot 
+ br[158] vdd vss bl[158] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_160_top 
+ br[158] vdd vss bl[158] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_161_bot 
+ br[159] vdd vss bl[159] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_161_top 
+ br[159] vdd vss bl[159] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_162_bot 
+ br[160] vdd vss bl[160] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_162_top 
+ br[160] vdd vss bl[160] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_163_bot 
+ br[161] vdd vss bl[161] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_163_top 
+ br[161] vdd vss bl[161] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_164_bot 
+ br[162] vdd vss bl[162] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_164_top 
+ br[162] vdd vss bl[162] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_165_bot 
+ br[163] vdd vss bl[163] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_165_top 
+ br[163] vdd vss bl[163] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_166_bot 
+ br[164] vdd vss bl[164] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_166_top 
+ br[164] vdd vss bl[164] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_167_bot 
+ br[165] vdd vss bl[165] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_167_top 
+ br[165] vdd vss bl[165] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_168_bot 
+ br[166] vdd vss bl[166] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_168_top 
+ br[166] vdd vss bl[166] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_169_bot 
+ br[167] vdd vss bl[167] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_169_top 
+ br[167] vdd vss bl[167] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_170_bot 
+ br[168] vdd vss bl[168] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_170_top 
+ br[168] vdd vss bl[168] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_171_bot 
+ br[169] vdd vss bl[169] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_171_top 
+ br[169] vdd vss bl[169] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_172_bot 
+ br[170] vdd vss bl[170] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_172_top 
+ br[170] vdd vss bl[170] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_173_bot 
+ br[171] vdd vss bl[171] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_173_top 
+ br[171] vdd vss bl[171] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_174_bot 
+ br[172] vdd vss bl[172] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_174_top 
+ br[172] vdd vss bl[172] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_175_bot 
+ br[173] vdd vss bl[173] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_175_top 
+ br[173] vdd vss bl[173] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_176_bot 
+ br[174] vdd vss bl[174] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_176_top 
+ br[174] vdd vss bl[174] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_177_bot 
+ br[175] vdd vss bl[175] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_177_top 
+ br[175] vdd vss bl[175] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_178_bot 
+ br[176] vdd vss bl[176] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_178_top 
+ br[176] vdd vss bl[176] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_179_bot 
+ br[177] vdd vss bl[177] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_179_top 
+ br[177] vdd vss bl[177] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_180_bot 
+ br[178] vdd vss bl[178] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_180_top 
+ br[178] vdd vss bl[178] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_181_bot 
+ br[179] vdd vss bl[179] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_181_top 
+ br[179] vdd vss bl[179] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_182_bot 
+ br[180] vdd vss bl[180] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_182_top 
+ br[180] vdd vss bl[180] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_183_bot 
+ br[181] vdd vss bl[181] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_183_top 
+ br[181] vdd vss bl[181] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_184_bot 
+ br[182] vdd vss bl[182] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_184_top 
+ br[182] vdd vss bl[182] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_185_bot 
+ br[183] vdd vss bl[183] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_185_top 
+ br[183] vdd vss bl[183] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_186_bot 
+ br[184] vdd vss bl[184] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_186_top 
+ br[184] vdd vss bl[184] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_187_bot 
+ br[185] vdd vss bl[185] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_187_top 
+ br[185] vdd vss bl[185] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_188_bot 
+ br[186] vdd vss bl[186] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_188_top 
+ br[186] vdd vss bl[186] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_189_bot 
+ br[187] vdd vss bl[187] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_189_top 
+ br[187] vdd vss bl[187] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_190_bot 
+ br[188] vdd vss bl[188] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_190_top 
+ br[188] vdd vss bl[188] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_191_bot 
+ br[189] vdd vss bl[189] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_191_top 
+ br[189] vdd vss bl[189] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_192_bot 
+ br[190] vdd vss bl[190] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_192_top 
+ br[190] vdd vss bl[190] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_193_bot 
+ br[191] vdd vss bl[191] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_193_top 
+ br[191] vdd vss bl[191] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_194_bot 
+ br[192] vdd vss bl[192] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_194_top 
+ br[192] vdd vss bl[192] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_195_bot 
+ br[193] vdd vss bl[193] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_195_top 
+ br[193] vdd vss bl[193] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_196_bot 
+ br[194] vdd vss bl[194] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_196_top 
+ br[194] vdd vss bl[194] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_197_bot 
+ br[195] vdd vss bl[195] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_197_top 
+ br[195] vdd vss bl[195] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_198_bot 
+ br[196] vdd vss bl[196] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_198_top 
+ br[196] vdd vss bl[196] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_199_bot 
+ br[197] vdd vss bl[197] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_199_top 
+ br[197] vdd vss bl[197] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_200_bot 
+ br[198] vdd vss bl[198] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_200_top 
+ br[198] vdd vss bl[198] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_201_bot 
+ br[199] vdd vss bl[199] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_201_top 
+ br[199] vdd vss bl[199] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_202_bot 
+ br[200] vdd vss bl[200] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_202_top 
+ br[200] vdd vss bl[200] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_203_bot 
+ br[201] vdd vss bl[201] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_203_top 
+ br[201] vdd vss bl[201] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_204_bot 
+ br[202] vdd vss bl[202] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_204_top 
+ br[202] vdd vss bl[202] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_205_bot 
+ br[203] vdd vss bl[203] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_205_top 
+ br[203] vdd vss bl[203] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_206_bot 
+ br[204] vdd vss bl[204] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_206_top 
+ br[204] vdd vss bl[204] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_207_bot 
+ br[205] vdd vss bl[205] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_207_top 
+ br[205] vdd vss bl[205] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_208_bot 
+ br[206] vdd vss bl[206] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_208_top 
+ br[206] vdd vss bl[206] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_209_bot 
+ br[207] vdd vss bl[207] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_209_top 
+ br[207] vdd vss bl[207] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_210_bot 
+ br[208] vdd vss bl[208] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_210_top 
+ br[208] vdd vss bl[208] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_211_bot 
+ br[209] vdd vss bl[209] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_211_top 
+ br[209] vdd vss bl[209] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_212_bot 
+ br[210] vdd vss bl[210] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_212_top 
+ br[210] vdd vss bl[210] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_213_bot 
+ br[211] vdd vss bl[211] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_213_top 
+ br[211] vdd vss bl[211] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_214_bot 
+ br[212] vdd vss bl[212] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_214_top 
+ br[212] vdd vss bl[212] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_215_bot 
+ br[213] vdd vss bl[213] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_215_top 
+ br[213] vdd vss bl[213] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_216_bot 
+ br[214] vdd vss bl[214] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_216_top 
+ br[214] vdd vss bl[214] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_217_bot 
+ br[215] vdd vss bl[215] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_217_top 
+ br[215] vdd vss bl[215] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_218_bot 
+ br[216] vdd vss bl[216] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_218_top 
+ br[216] vdd vss bl[216] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_219_bot 
+ br[217] vdd vss bl[217] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_219_top 
+ br[217] vdd vss bl[217] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_220_bot 
+ br[218] vdd vss bl[218] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_220_top 
+ br[218] vdd vss bl[218] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_221_bot 
+ br[219] vdd vss bl[219] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_221_top 
+ br[219] vdd vss bl[219] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_222_bot 
+ br[220] vdd vss bl[220] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_222_top 
+ br[220] vdd vss bl[220] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_223_bot 
+ br[221] vdd vss bl[221] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_223_top 
+ br[221] vdd vss bl[221] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_224_bot 
+ br[222] vdd vss bl[222] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_224_top 
+ br[222] vdd vss bl[222] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_225_bot 
+ br[223] vdd vss bl[223] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_225_top 
+ br[223] vdd vss bl[223] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_226_bot 
+ br[224] vdd vss bl[224] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_226_top 
+ br[224] vdd vss bl[224] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_227_bot 
+ br[225] vdd vss bl[225] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_227_top 
+ br[225] vdd vss bl[225] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_228_bot 
+ br[226] vdd vss bl[226] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_228_top 
+ br[226] vdd vss bl[226] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_229_bot 
+ br[227] vdd vss bl[227] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_229_top 
+ br[227] vdd vss bl[227] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_230_bot 
+ br[228] vdd vss bl[228] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_230_top 
+ br[228] vdd vss bl[228] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_231_bot 
+ br[229] vdd vss bl[229] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_231_top 
+ br[229] vdd vss bl[229] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_232_bot 
+ br[230] vdd vss bl[230] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_232_top 
+ br[230] vdd vss bl[230] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_233_bot 
+ br[231] vdd vss bl[231] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_233_top 
+ br[231] vdd vss bl[231] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_234_bot 
+ br[232] vdd vss bl[232] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_234_top 
+ br[232] vdd vss bl[232] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_235_bot 
+ br[233] vdd vss bl[233] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_235_top 
+ br[233] vdd vss bl[233] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_236_bot 
+ br[234] vdd vss bl[234] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_236_top 
+ br[234] vdd vss bl[234] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_237_bot 
+ br[235] vdd vss bl[235] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_237_top 
+ br[235] vdd vss bl[235] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_238_bot 
+ br[236] vdd vss bl[236] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_238_top 
+ br[236] vdd vss bl[236] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_239_bot 
+ br[237] vdd vss bl[237] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_239_top 
+ br[237] vdd vss bl[237] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_240_bot 
+ br[238] vdd vss bl[238] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_240_top 
+ br[238] vdd vss bl[238] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_241_bot 
+ br[239] vdd vss bl[239] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_241_top 
+ br[239] vdd vss bl[239] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_242_bot 
+ br[240] vdd vss bl[240] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_242_top 
+ br[240] vdd vss bl[240] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_243_bot 
+ br[241] vdd vss bl[241] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_243_top 
+ br[241] vdd vss bl[241] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_244_bot 
+ br[242] vdd vss bl[242] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_244_top 
+ br[242] vdd vss bl[242] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_245_bot 
+ br[243] vdd vss bl[243] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_245_top 
+ br[243] vdd vss bl[243] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_246_bot 
+ br[244] vdd vss bl[244] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_246_top 
+ br[244] vdd vss bl[244] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_247_bot 
+ br[245] vdd vss bl[245] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_247_top 
+ br[245] vdd vss bl[245] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_248_bot 
+ br[246] vdd vss bl[246] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_248_top 
+ br[246] vdd vss bl[246] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_249_bot 
+ br[247] vdd vss bl[247] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_249_top 
+ br[247] vdd vss bl[247] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_250_bot 
+ br[248] vdd vss bl[248] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_250_top 
+ br[248] vdd vss bl[248] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_251_bot 
+ br[249] vdd vss bl[249] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_251_top 
+ br[249] vdd vss bl[249] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_252_bot 
+ br[250] vdd vss bl[250] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_252_top 
+ br[250] vdd vss bl[250] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_253_bot 
+ br[251] vdd vss bl[251] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_253_top 
+ br[251] vdd vss bl[251] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_254_bot 
+ br[252] vdd vss bl[252] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_254_top 
+ br[252] vdd vss bl[252] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_255_bot 
+ br[253] vdd vss bl[253] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_255_top 
+ br[253] vdd vss bl[253] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_256_bot 
+ br[254] vdd vss bl[254] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_256_top 
+ br[254] vdd vss bl[254] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_257_bot 
+ br[255] vdd vss bl[255] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_257_top 
+ br[255] vdd vss bl[255] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_258_bot 
+ vdd vdd vss vdd vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_258_top 
+ vdd vdd vss vdd vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_259_bot 
+ vdd vdd vss vdd vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_259_top 
+ vdd vdd vss vdd vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

.ENDS

.SUBCKT precharge 
+ vdd bl br en_b 

xbl_pull_up 
+ bl en_b vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='1.0' l='0.15' 

xbr_pull_up 
+ br en_b vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='1.0' l='0.15' 

xequalizer 
+ bl en_b br vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='1.0' l='0.15' 

.ENDS

.SUBCKT precharge_array 
+ vdd en_b bl[256] bl[255] bl[254] bl[253] bl[252] bl[251] bl[250] bl[249] bl[248] bl[247] bl[246] bl[245] bl[244] bl[243] bl[242] bl[241] bl[240] bl[239] bl[238] bl[237] bl[236] bl[235] bl[234] bl[233] bl[232] bl[231] bl[230] bl[229] bl[228] bl[227] bl[226] bl[225] bl[224] bl[223] bl[222] bl[221] bl[220] bl[219] bl[218] bl[217] bl[216] bl[215] bl[214] bl[213] bl[212] bl[211] bl[210] bl[209] bl[208] bl[207] bl[206] bl[205] bl[204] bl[203] bl[202] bl[201] bl[200] bl[199] bl[198] bl[197] bl[196] bl[195] bl[194] bl[193] bl[192] bl[191] bl[190] bl[189] bl[188] bl[187] bl[186] bl[185] bl[184] bl[183] bl[182] bl[181] bl[180] bl[179] bl[178] bl[177] bl[176] bl[175] bl[174] bl[173] bl[172] bl[171] bl[170] bl[169] bl[168] bl[167] bl[166] bl[165] bl[164] bl[163] bl[162] bl[161] bl[160] bl[159] bl[158] bl[157] bl[156] bl[155] bl[154] bl[153] bl[152] bl[151] bl[150] bl[149] bl[148] bl[147] bl[146] bl[145] bl[144] bl[143] bl[142] bl[141] bl[140] bl[139] bl[138] bl[137] bl[136] bl[135] bl[134] bl[133] bl[132] bl[131] bl[130] bl[129] bl[128] bl[127] bl[126] bl[125] bl[124] bl[123] bl[122] bl[121] bl[120] bl[119] bl[118] bl[117] bl[116] bl[115] bl[114] bl[113] bl[112] bl[111] bl[110] bl[109] bl[108] bl[107] bl[106] bl[105] bl[104] bl[103] bl[102] bl[101] bl[100] bl[99] bl[98] bl[97] bl[96] bl[95] bl[94] bl[93] bl[92] bl[91] bl[90] bl[89] bl[88] bl[87] bl[86] bl[85] bl[84] bl[83] bl[82] bl[81] bl[80] bl[79] bl[78] bl[77] bl[76] bl[75] bl[74] bl[73] bl[72] bl[71] bl[70] bl[69] bl[68] bl[67] bl[66] bl[65] bl[64] bl[63] bl[62] bl[61] bl[60] bl[59] bl[58] bl[57] bl[56] bl[55] bl[54] bl[53] bl[52] bl[51] bl[50] bl[49] bl[48] bl[47] bl[46] bl[45] bl[44] bl[43] bl[42] bl[41] bl[40] bl[39] bl[38] bl[37] bl[36] bl[35] bl[34] bl[33] bl[32] bl[31] bl[30] bl[29] bl[28] bl[27] bl[26] bl[25] bl[24] bl[23] bl[22] bl[21] bl[20] bl[19] bl[18] bl[17] bl[16] bl[15] bl[14] bl[13] bl[12] bl[11] bl[10] bl[9] bl[8] bl[7] bl[6] bl[5] bl[4] bl[3] bl[2] bl[1] bl[0] br[256] br[255] br[254] br[253] br[252] br[251] br[250] br[249] br[248] br[247] br[246] br[245] br[244] br[243] br[242] br[241] br[240] br[239] br[238] br[237] br[236] br[235] br[234] br[233] br[232] br[231] br[230] br[229] br[228] br[227] br[226] br[225] br[224] br[223] br[222] br[221] br[220] br[219] br[218] br[217] br[216] br[215] br[214] br[213] br[212] br[211] br[210] br[209] br[208] br[207] br[206] br[205] br[204] br[203] br[202] br[201] br[200] br[199] br[198] br[197] br[196] br[195] br[194] br[193] br[192] br[191] br[190] br[189] br[188] br[187] br[186] br[185] br[184] br[183] br[182] br[181] br[180] br[179] br[178] br[177] br[176] br[175] br[174] br[173] br[172] br[171] br[170] br[169] br[168] br[167] br[166] br[165] br[164] br[163] br[162] br[161] br[160] br[159] br[158] br[157] br[156] br[155] br[154] br[153] br[152] br[151] br[150] br[149] br[148] br[147] br[146] br[145] br[144] br[143] br[142] br[141] br[140] br[139] br[138] br[137] br[136] br[135] br[134] br[133] br[132] br[131] br[130] br[129] br[128] br[127] br[126] br[125] br[124] br[123] br[122] br[121] br[120] br[119] br[118] br[117] br[116] br[115] br[114] br[113] br[112] br[111] br[110] br[109] br[108] br[107] br[106] br[105] br[104] br[103] br[102] br[101] br[100] br[99] br[98] br[97] br[96] br[95] br[94] br[93] br[92] br[91] br[90] br[89] br[88] br[87] br[86] br[85] br[84] br[83] br[82] br[81] br[80] br[79] br[78] br[77] br[76] br[75] br[74] br[73] br[72] br[71] br[70] br[69] br[68] br[67] br[66] br[65] br[64] br[63] br[62] br[61] br[60] br[59] br[58] br[57] br[56] br[55] br[54] br[53] br[52] br[51] br[50] br[49] br[48] br[47] br[46] br[45] br[44] br[43] br[42] br[41] br[40] br[39] br[38] br[37] br[36] br[35] br[34] br[33] br[32] br[31] br[30] br[29] br[28] br[27] br[26] br[25] br[24] br[23] br[22] br[21] br[20] br[19] br[18] br[17] br[16] br[15] br[14] br[13] br[12] br[11] br[10] br[9] br[8] br[7] br[6] br[5] br[4] br[3] br[2] br[1] br[0] 

xprecharge_0 
+ vdd bl[0] br[0] en_b 
+ precharge 
* No parameters

xprecharge_1 
+ vdd bl[1] br[1] en_b 
+ precharge 
* No parameters

xprecharge_2 
+ vdd bl[2] br[2] en_b 
+ precharge 
* No parameters

xprecharge_3 
+ vdd bl[3] br[3] en_b 
+ precharge 
* No parameters

xprecharge_4 
+ vdd bl[4] br[4] en_b 
+ precharge 
* No parameters

xprecharge_5 
+ vdd bl[5] br[5] en_b 
+ precharge 
* No parameters

xprecharge_6 
+ vdd bl[6] br[6] en_b 
+ precharge 
* No parameters

xprecharge_7 
+ vdd bl[7] br[7] en_b 
+ precharge 
* No parameters

xprecharge_8 
+ vdd bl[8] br[8] en_b 
+ precharge 
* No parameters

xprecharge_9 
+ vdd bl[9] br[9] en_b 
+ precharge 
* No parameters

xprecharge_10 
+ vdd bl[10] br[10] en_b 
+ precharge 
* No parameters

xprecharge_11 
+ vdd bl[11] br[11] en_b 
+ precharge 
* No parameters

xprecharge_12 
+ vdd bl[12] br[12] en_b 
+ precharge 
* No parameters

xprecharge_13 
+ vdd bl[13] br[13] en_b 
+ precharge 
* No parameters

xprecharge_14 
+ vdd bl[14] br[14] en_b 
+ precharge 
* No parameters

xprecharge_15 
+ vdd bl[15] br[15] en_b 
+ precharge 
* No parameters

xprecharge_16 
+ vdd bl[16] br[16] en_b 
+ precharge 
* No parameters

xprecharge_17 
+ vdd bl[17] br[17] en_b 
+ precharge 
* No parameters

xprecharge_18 
+ vdd bl[18] br[18] en_b 
+ precharge 
* No parameters

xprecharge_19 
+ vdd bl[19] br[19] en_b 
+ precharge 
* No parameters

xprecharge_20 
+ vdd bl[20] br[20] en_b 
+ precharge 
* No parameters

xprecharge_21 
+ vdd bl[21] br[21] en_b 
+ precharge 
* No parameters

xprecharge_22 
+ vdd bl[22] br[22] en_b 
+ precharge 
* No parameters

xprecharge_23 
+ vdd bl[23] br[23] en_b 
+ precharge 
* No parameters

xprecharge_24 
+ vdd bl[24] br[24] en_b 
+ precharge 
* No parameters

xprecharge_25 
+ vdd bl[25] br[25] en_b 
+ precharge 
* No parameters

xprecharge_26 
+ vdd bl[26] br[26] en_b 
+ precharge 
* No parameters

xprecharge_27 
+ vdd bl[27] br[27] en_b 
+ precharge 
* No parameters

xprecharge_28 
+ vdd bl[28] br[28] en_b 
+ precharge 
* No parameters

xprecharge_29 
+ vdd bl[29] br[29] en_b 
+ precharge 
* No parameters

xprecharge_30 
+ vdd bl[30] br[30] en_b 
+ precharge 
* No parameters

xprecharge_31 
+ vdd bl[31] br[31] en_b 
+ precharge 
* No parameters

xprecharge_32 
+ vdd bl[32] br[32] en_b 
+ precharge 
* No parameters

xprecharge_33 
+ vdd bl[33] br[33] en_b 
+ precharge 
* No parameters

xprecharge_34 
+ vdd bl[34] br[34] en_b 
+ precharge 
* No parameters

xprecharge_35 
+ vdd bl[35] br[35] en_b 
+ precharge 
* No parameters

xprecharge_36 
+ vdd bl[36] br[36] en_b 
+ precharge 
* No parameters

xprecharge_37 
+ vdd bl[37] br[37] en_b 
+ precharge 
* No parameters

xprecharge_38 
+ vdd bl[38] br[38] en_b 
+ precharge 
* No parameters

xprecharge_39 
+ vdd bl[39] br[39] en_b 
+ precharge 
* No parameters

xprecharge_40 
+ vdd bl[40] br[40] en_b 
+ precharge 
* No parameters

xprecharge_41 
+ vdd bl[41] br[41] en_b 
+ precharge 
* No parameters

xprecharge_42 
+ vdd bl[42] br[42] en_b 
+ precharge 
* No parameters

xprecharge_43 
+ vdd bl[43] br[43] en_b 
+ precharge 
* No parameters

xprecharge_44 
+ vdd bl[44] br[44] en_b 
+ precharge 
* No parameters

xprecharge_45 
+ vdd bl[45] br[45] en_b 
+ precharge 
* No parameters

xprecharge_46 
+ vdd bl[46] br[46] en_b 
+ precharge 
* No parameters

xprecharge_47 
+ vdd bl[47] br[47] en_b 
+ precharge 
* No parameters

xprecharge_48 
+ vdd bl[48] br[48] en_b 
+ precharge 
* No parameters

xprecharge_49 
+ vdd bl[49] br[49] en_b 
+ precharge 
* No parameters

xprecharge_50 
+ vdd bl[50] br[50] en_b 
+ precharge 
* No parameters

xprecharge_51 
+ vdd bl[51] br[51] en_b 
+ precharge 
* No parameters

xprecharge_52 
+ vdd bl[52] br[52] en_b 
+ precharge 
* No parameters

xprecharge_53 
+ vdd bl[53] br[53] en_b 
+ precharge 
* No parameters

xprecharge_54 
+ vdd bl[54] br[54] en_b 
+ precharge 
* No parameters

xprecharge_55 
+ vdd bl[55] br[55] en_b 
+ precharge 
* No parameters

xprecharge_56 
+ vdd bl[56] br[56] en_b 
+ precharge 
* No parameters

xprecharge_57 
+ vdd bl[57] br[57] en_b 
+ precharge 
* No parameters

xprecharge_58 
+ vdd bl[58] br[58] en_b 
+ precharge 
* No parameters

xprecharge_59 
+ vdd bl[59] br[59] en_b 
+ precharge 
* No parameters

xprecharge_60 
+ vdd bl[60] br[60] en_b 
+ precharge 
* No parameters

xprecharge_61 
+ vdd bl[61] br[61] en_b 
+ precharge 
* No parameters

xprecharge_62 
+ vdd bl[62] br[62] en_b 
+ precharge 
* No parameters

xprecharge_63 
+ vdd bl[63] br[63] en_b 
+ precharge 
* No parameters

xprecharge_64 
+ vdd bl[64] br[64] en_b 
+ precharge 
* No parameters

xprecharge_65 
+ vdd bl[65] br[65] en_b 
+ precharge 
* No parameters

xprecharge_66 
+ vdd bl[66] br[66] en_b 
+ precharge 
* No parameters

xprecharge_67 
+ vdd bl[67] br[67] en_b 
+ precharge 
* No parameters

xprecharge_68 
+ vdd bl[68] br[68] en_b 
+ precharge 
* No parameters

xprecharge_69 
+ vdd bl[69] br[69] en_b 
+ precharge 
* No parameters

xprecharge_70 
+ vdd bl[70] br[70] en_b 
+ precharge 
* No parameters

xprecharge_71 
+ vdd bl[71] br[71] en_b 
+ precharge 
* No parameters

xprecharge_72 
+ vdd bl[72] br[72] en_b 
+ precharge 
* No parameters

xprecharge_73 
+ vdd bl[73] br[73] en_b 
+ precharge 
* No parameters

xprecharge_74 
+ vdd bl[74] br[74] en_b 
+ precharge 
* No parameters

xprecharge_75 
+ vdd bl[75] br[75] en_b 
+ precharge 
* No parameters

xprecharge_76 
+ vdd bl[76] br[76] en_b 
+ precharge 
* No parameters

xprecharge_77 
+ vdd bl[77] br[77] en_b 
+ precharge 
* No parameters

xprecharge_78 
+ vdd bl[78] br[78] en_b 
+ precharge 
* No parameters

xprecharge_79 
+ vdd bl[79] br[79] en_b 
+ precharge 
* No parameters

xprecharge_80 
+ vdd bl[80] br[80] en_b 
+ precharge 
* No parameters

xprecharge_81 
+ vdd bl[81] br[81] en_b 
+ precharge 
* No parameters

xprecharge_82 
+ vdd bl[82] br[82] en_b 
+ precharge 
* No parameters

xprecharge_83 
+ vdd bl[83] br[83] en_b 
+ precharge 
* No parameters

xprecharge_84 
+ vdd bl[84] br[84] en_b 
+ precharge 
* No parameters

xprecharge_85 
+ vdd bl[85] br[85] en_b 
+ precharge 
* No parameters

xprecharge_86 
+ vdd bl[86] br[86] en_b 
+ precharge 
* No parameters

xprecharge_87 
+ vdd bl[87] br[87] en_b 
+ precharge 
* No parameters

xprecharge_88 
+ vdd bl[88] br[88] en_b 
+ precharge 
* No parameters

xprecharge_89 
+ vdd bl[89] br[89] en_b 
+ precharge 
* No parameters

xprecharge_90 
+ vdd bl[90] br[90] en_b 
+ precharge 
* No parameters

xprecharge_91 
+ vdd bl[91] br[91] en_b 
+ precharge 
* No parameters

xprecharge_92 
+ vdd bl[92] br[92] en_b 
+ precharge 
* No parameters

xprecharge_93 
+ vdd bl[93] br[93] en_b 
+ precharge 
* No parameters

xprecharge_94 
+ vdd bl[94] br[94] en_b 
+ precharge 
* No parameters

xprecharge_95 
+ vdd bl[95] br[95] en_b 
+ precharge 
* No parameters

xprecharge_96 
+ vdd bl[96] br[96] en_b 
+ precharge 
* No parameters

xprecharge_97 
+ vdd bl[97] br[97] en_b 
+ precharge 
* No parameters

xprecharge_98 
+ vdd bl[98] br[98] en_b 
+ precharge 
* No parameters

xprecharge_99 
+ vdd bl[99] br[99] en_b 
+ precharge 
* No parameters

xprecharge_100 
+ vdd bl[100] br[100] en_b 
+ precharge 
* No parameters

xprecharge_101 
+ vdd bl[101] br[101] en_b 
+ precharge 
* No parameters

xprecharge_102 
+ vdd bl[102] br[102] en_b 
+ precharge 
* No parameters

xprecharge_103 
+ vdd bl[103] br[103] en_b 
+ precharge 
* No parameters

xprecharge_104 
+ vdd bl[104] br[104] en_b 
+ precharge 
* No parameters

xprecharge_105 
+ vdd bl[105] br[105] en_b 
+ precharge 
* No parameters

xprecharge_106 
+ vdd bl[106] br[106] en_b 
+ precharge 
* No parameters

xprecharge_107 
+ vdd bl[107] br[107] en_b 
+ precharge 
* No parameters

xprecharge_108 
+ vdd bl[108] br[108] en_b 
+ precharge 
* No parameters

xprecharge_109 
+ vdd bl[109] br[109] en_b 
+ precharge 
* No parameters

xprecharge_110 
+ vdd bl[110] br[110] en_b 
+ precharge 
* No parameters

xprecharge_111 
+ vdd bl[111] br[111] en_b 
+ precharge 
* No parameters

xprecharge_112 
+ vdd bl[112] br[112] en_b 
+ precharge 
* No parameters

xprecharge_113 
+ vdd bl[113] br[113] en_b 
+ precharge 
* No parameters

xprecharge_114 
+ vdd bl[114] br[114] en_b 
+ precharge 
* No parameters

xprecharge_115 
+ vdd bl[115] br[115] en_b 
+ precharge 
* No parameters

xprecharge_116 
+ vdd bl[116] br[116] en_b 
+ precharge 
* No parameters

xprecharge_117 
+ vdd bl[117] br[117] en_b 
+ precharge 
* No parameters

xprecharge_118 
+ vdd bl[118] br[118] en_b 
+ precharge 
* No parameters

xprecharge_119 
+ vdd bl[119] br[119] en_b 
+ precharge 
* No parameters

xprecharge_120 
+ vdd bl[120] br[120] en_b 
+ precharge 
* No parameters

xprecharge_121 
+ vdd bl[121] br[121] en_b 
+ precharge 
* No parameters

xprecharge_122 
+ vdd bl[122] br[122] en_b 
+ precharge 
* No parameters

xprecharge_123 
+ vdd bl[123] br[123] en_b 
+ precharge 
* No parameters

xprecharge_124 
+ vdd bl[124] br[124] en_b 
+ precharge 
* No parameters

xprecharge_125 
+ vdd bl[125] br[125] en_b 
+ precharge 
* No parameters

xprecharge_126 
+ vdd bl[126] br[126] en_b 
+ precharge 
* No parameters

xprecharge_127 
+ vdd bl[127] br[127] en_b 
+ precharge 
* No parameters

xprecharge_128 
+ vdd bl[128] br[128] en_b 
+ precharge 
* No parameters

xprecharge_129 
+ vdd bl[129] br[129] en_b 
+ precharge 
* No parameters

xprecharge_130 
+ vdd bl[130] br[130] en_b 
+ precharge 
* No parameters

xprecharge_131 
+ vdd bl[131] br[131] en_b 
+ precharge 
* No parameters

xprecharge_132 
+ vdd bl[132] br[132] en_b 
+ precharge 
* No parameters

xprecharge_133 
+ vdd bl[133] br[133] en_b 
+ precharge 
* No parameters

xprecharge_134 
+ vdd bl[134] br[134] en_b 
+ precharge 
* No parameters

xprecharge_135 
+ vdd bl[135] br[135] en_b 
+ precharge 
* No parameters

xprecharge_136 
+ vdd bl[136] br[136] en_b 
+ precharge 
* No parameters

xprecharge_137 
+ vdd bl[137] br[137] en_b 
+ precharge 
* No parameters

xprecharge_138 
+ vdd bl[138] br[138] en_b 
+ precharge 
* No parameters

xprecharge_139 
+ vdd bl[139] br[139] en_b 
+ precharge 
* No parameters

xprecharge_140 
+ vdd bl[140] br[140] en_b 
+ precharge 
* No parameters

xprecharge_141 
+ vdd bl[141] br[141] en_b 
+ precharge 
* No parameters

xprecharge_142 
+ vdd bl[142] br[142] en_b 
+ precharge 
* No parameters

xprecharge_143 
+ vdd bl[143] br[143] en_b 
+ precharge 
* No parameters

xprecharge_144 
+ vdd bl[144] br[144] en_b 
+ precharge 
* No parameters

xprecharge_145 
+ vdd bl[145] br[145] en_b 
+ precharge 
* No parameters

xprecharge_146 
+ vdd bl[146] br[146] en_b 
+ precharge 
* No parameters

xprecharge_147 
+ vdd bl[147] br[147] en_b 
+ precharge 
* No parameters

xprecharge_148 
+ vdd bl[148] br[148] en_b 
+ precharge 
* No parameters

xprecharge_149 
+ vdd bl[149] br[149] en_b 
+ precharge 
* No parameters

xprecharge_150 
+ vdd bl[150] br[150] en_b 
+ precharge 
* No parameters

xprecharge_151 
+ vdd bl[151] br[151] en_b 
+ precharge 
* No parameters

xprecharge_152 
+ vdd bl[152] br[152] en_b 
+ precharge 
* No parameters

xprecharge_153 
+ vdd bl[153] br[153] en_b 
+ precharge 
* No parameters

xprecharge_154 
+ vdd bl[154] br[154] en_b 
+ precharge 
* No parameters

xprecharge_155 
+ vdd bl[155] br[155] en_b 
+ precharge 
* No parameters

xprecharge_156 
+ vdd bl[156] br[156] en_b 
+ precharge 
* No parameters

xprecharge_157 
+ vdd bl[157] br[157] en_b 
+ precharge 
* No parameters

xprecharge_158 
+ vdd bl[158] br[158] en_b 
+ precharge 
* No parameters

xprecharge_159 
+ vdd bl[159] br[159] en_b 
+ precharge 
* No parameters

xprecharge_160 
+ vdd bl[160] br[160] en_b 
+ precharge 
* No parameters

xprecharge_161 
+ vdd bl[161] br[161] en_b 
+ precharge 
* No parameters

xprecharge_162 
+ vdd bl[162] br[162] en_b 
+ precharge 
* No parameters

xprecharge_163 
+ vdd bl[163] br[163] en_b 
+ precharge 
* No parameters

xprecharge_164 
+ vdd bl[164] br[164] en_b 
+ precharge 
* No parameters

xprecharge_165 
+ vdd bl[165] br[165] en_b 
+ precharge 
* No parameters

xprecharge_166 
+ vdd bl[166] br[166] en_b 
+ precharge 
* No parameters

xprecharge_167 
+ vdd bl[167] br[167] en_b 
+ precharge 
* No parameters

xprecharge_168 
+ vdd bl[168] br[168] en_b 
+ precharge 
* No parameters

xprecharge_169 
+ vdd bl[169] br[169] en_b 
+ precharge 
* No parameters

xprecharge_170 
+ vdd bl[170] br[170] en_b 
+ precharge 
* No parameters

xprecharge_171 
+ vdd bl[171] br[171] en_b 
+ precharge 
* No parameters

xprecharge_172 
+ vdd bl[172] br[172] en_b 
+ precharge 
* No parameters

xprecharge_173 
+ vdd bl[173] br[173] en_b 
+ precharge 
* No parameters

xprecharge_174 
+ vdd bl[174] br[174] en_b 
+ precharge 
* No parameters

xprecharge_175 
+ vdd bl[175] br[175] en_b 
+ precharge 
* No parameters

xprecharge_176 
+ vdd bl[176] br[176] en_b 
+ precharge 
* No parameters

xprecharge_177 
+ vdd bl[177] br[177] en_b 
+ precharge 
* No parameters

xprecharge_178 
+ vdd bl[178] br[178] en_b 
+ precharge 
* No parameters

xprecharge_179 
+ vdd bl[179] br[179] en_b 
+ precharge 
* No parameters

xprecharge_180 
+ vdd bl[180] br[180] en_b 
+ precharge 
* No parameters

xprecharge_181 
+ vdd bl[181] br[181] en_b 
+ precharge 
* No parameters

xprecharge_182 
+ vdd bl[182] br[182] en_b 
+ precharge 
* No parameters

xprecharge_183 
+ vdd bl[183] br[183] en_b 
+ precharge 
* No parameters

xprecharge_184 
+ vdd bl[184] br[184] en_b 
+ precharge 
* No parameters

xprecharge_185 
+ vdd bl[185] br[185] en_b 
+ precharge 
* No parameters

xprecharge_186 
+ vdd bl[186] br[186] en_b 
+ precharge 
* No parameters

xprecharge_187 
+ vdd bl[187] br[187] en_b 
+ precharge 
* No parameters

xprecharge_188 
+ vdd bl[188] br[188] en_b 
+ precharge 
* No parameters

xprecharge_189 
+ vdd bl[189] br[189] en_b 
+ precharge 
* No parameters

xprecharge_190 
+ vdd bl[190] br[190] en_b 
+ precharge 
* No parameters

xprecharge_191 
+ vdd bl[191] br[191] en_b 
+ precharge 
* No parameters

xprecharge_192 
+ vdd bl[192] br[192] en_b 
+ precharge 
* No parameters

xprecharge_193 
+ vdd bl[193] br[193] en_b 
+ precharge 
* No parameters

xprecharge_194 
+ vdd bl[194] br[194] en_b 
+ precharge 
* No parameters

xprecharge_195 
+ vdd bl[195] br[195] en_b 
+ precharge 
* No parameters

xprecharge_196 
+ vdd bl[196] br[196] en_b 
+ precharge 
* No parameters

xprecharge_197 
+ vdd bl[197] br[197] en_b 
+ precharge 
* No parameters

xprecharge_198 
+ vdd bl[198] br[198] en_b 
+ precharge 
* No parameters

xprecharge_199 
+ vdd bl[199] br[199] en_b 
+ precharge 
* No parameters

xprecharge_200 
+ vdd bl[200] br[200] en_b 
+ precharge 
* No parameters

xprecharge_201 
+ vdd bl[201] br[201] en_b 
+ precharge 
* No parameters

xprecharge_202 
+ vdd bl[202] br[202] en_b 
+ precharge 
* No parameters

xprecharge_203 
+ vdd bl[203] br[203] en_b 
+ precharge 
* No parameters

xprecharge_204 
+ vdd bl[204] br[204] en_b 
+ precharge 
* No parameters

xprecharge_205 
+ vdd bl[205] br[205] en_b 
+ precharge 
* No parameters

xprecharge_206 
+ vdd bl[206] br[206] en_b 
+ precharge 
* No parameters

xprecharge_207 
+ vdd bl[207] br[207] en_b 
+ precharge 
* No parameters

xprecharge_208 
+ vdd bl[208] br[208] en_b 
+ precharge 
* No parameters

xprecharge_209 
+ vdd bl[209] br[209] en_b 
+ precharge 
* No parameters

xprecharge_210 
+ vdd bl[210] br[210] en_b 
+ precharge 
* No parameters

xprecharge_211 
+ vdd bl[211] br[211] en_b 
+ precharge 
* No parameters

xprecharge_212 
+ vdd bl[212] br[212] en_b 
+ precharge 
* No parameters

xprecharge_213 
+ vdd bl[213] br[213] en_b 
+ precharge 
* No parameters

xprecharge_214 
+ vdd bl[214] br[214] en_b 
+ precharge 
* No parameters

xprecharge_215 
+ vdd bl[215] br[215] en_b 
+ precharge 
* No parameters

xprecharge_216 
+ vdd bl[216] br[216] en_b 
+ precharge 
* No parameters

xprecharge_217 
+ vdd bl[217] br[217] en_b 
+ precharge 
* No parameters

xprecharge_218 
+ vdd bl[218] br[218] en_b 
+ precharge 
* No parameters

xprecharge_219 
+ vdd bl[219] br[219] en_b 
+ precharge 
* No parameters

xprecharge_220 
+ vdd bl[220] br[220] en_b 
+ precharge 
* No parameters

xprecharge_221 
+ vdd bl[221] br[221] en_b 
+ precharge 
* No parameters

xprecharge_222 
+ vdd bl[222] br[222] en_b 
+ precharge 
* No parameters

xprecharge_223 
+ vdd bl[223] br[223] en_b 
+ precharge 
* No parameters

xprecharge_224 
+ vdd bl[224] br[224] en_b 
+ precharge 
* No parameters

xprecharge_225 
+ vdd bl[225] br[225] en_b 
+ precharge 
* No parameters

xprecharge_226 
+ vdd bl[226] br[226] en_b 
+ precharge 
* No parameters

xprecharge_227 
+ vdd bl[227] br[227] en_b 
+ precharge 
* No parameters

xprecharge_228 
+ vdd bl[228] br[228] en_b 
+ precharge 
* No parameters

xprecharge_229 
+ vdd bl[229] br[229] en_b 
+ precharge 
* No parameters

xprecharge_230 
+ vdd bl[230] br[230] en_b 
+ precharge 
* No parameters

xprecharge_231 
+ vdd bl[231] br[231] en_b 
+ precharge 
* No parameters

xprecharge_232 
+ vdd bl[232] br[232] en_b 
+ precharge 
* No parameters

xprecharge_233 
+ vdd bl[233] br[233] en_b 
+ precharge 
* No parameters

xprecharge_234 
+ vdd bl[234] br[234] en_b 
+ precharge 
* No parameters

xprecharge_235 
+ vdd bl[235] br[235] en_b 
+ precharge 
* No parameters

xprecharge_236 
+ vdd bl[236] br[236] en_b 
+ precharge 
* No parameters

xprecharge_237 
+ vdd bl[237] br[237] en_b 
+ precharge 
* No parameters

xprecharge_238 
+ vdd bl[238] br[238] en_b 
+ precharge 
* No parameters

xprecharge_239 
+ vdd bl[239] br[239] en_b 
+ precharge 
* No parameters

xprecharge_240 
+ vdd bl[240] br[240] en_b 
+ precharge 
* No parameters

xprecharge_241 
+ vdd bl[241] br[241] en_b 
+ precharge 
* No parameters

xprecharge_242 
+ vdd bl[242] br[242] en_b 
+ precharge 
* No parameters

xprecharge_243 
+ vdd bl[243] br[243] en_b 
+ precharge 
* No parameters

xprecharge_244 
+ vdd bl[244] br[244] en_b 
+ precharge 
* No parameters

xprecharge_245 
+ vdd bl[245] br[245] en_b 
+ precharge 
* No parameters

xprecharge_246 
+ vdd bl[246] br[246] en_b 
+ precharge 
* No parameters

xprecharge_247 
+ vdd bl[247] br[247] en_b 
+ precharge 
* No parameters

xprecharge_248 
+ vdd bl[248] br[248] en_b 
+ precharge 
* No parameters

xprecharge_249 
+ vdd bl[249] br[249] en_b 
+ precharge 
* No parameters

xprecharge_250 
+ vdd bl[250] br[250] en_b 
+ precharge 
* No parameters

xprecharge_251 
+ vdd bl[251] br[251] en_b 
+ precharge 
* No parameters

xprecharge_252 
+ vdd bl[252] br[252] en_b 
+ precharge 
* No parameters

xprecharge_253 
+ vdd bl[253] br[253] en_b 
+ precharge 
* No parameters

xprecharge_254 
+ vdd bl[254] br[254] en_b 
+ precharge 
* No parameters

xprecharge_255 
+ vdd bl[255] br[255] en_b 
+ precharge 
* No parameters

xprecharge_256 
+ vdd bl[256] br[256] en_b 
+ precharge 
* No parameters

.ENDS

.SUBCKT read_mux 
+ sel_b bl br bl_out br_out vdd 

xMBL 
+ bl_out sel_b bl vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='1.2' l='0.15' 

xMBR 
+ br_out sel_b br vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='1.2' l='0.15' 

.ENDS

.SUBCKT read_mux_array 
+ sel_b[7] sel_b[6] sel_b[5] sel_b[4] sel_b[3] sel_b[2] sel_b[1] sel_b[0] bl[255] bl[254] bl[253] bl[252] bl[251] bl[250] bl[249] bl[248] bl[247] bl[246] bl[245] bl[244] bl[243] bl[242] bl[241] bl[240] bl[239] bl[238] bl[237] bl[236] bl[235] bl[234] bl[233] bl[232] bl[231] bl[230] bl[229] bl[228] bl[227] bl[226] bl[225] bl[224] bl[223] bl[222] bl[221] bl[220] bl[219] bl[218] bl[217] bl[216] bl[215] bl[214] bl[213] bl[212] bl[211] bl[210] bl[209] bl[208] bl[207] bl[206] bl[205] bl[204] bl[203] bl[202] bl[201] bl[200] bl[199] bl[198] bl[197] bl[196] bl[195] bl[194] bl[193] bl[192] bl[191] bl[190] bl[189] bl[188] bl[187] bl[186] bl[185] bl[184] bl[183] bl[182] bl[181] bl[180] bl[179] bl[178] bl[177] bl[176] bl[175] bl[174] bl[173] bl[172] bl[171] bl[170] bl[169] bl[168] bl[167] bl[166] bl[165] bl[164] bl[163] bl[162] bl[161] bl[160] bl[159] bl[158] bl[157] bl[156] bl[155] bl[154] bl[153] bl[152] bl[151] bl[150] bl[149] bl[148] bl[147] bl[146] bl[145] bl[144] bl[143] bl[142] bl[141] bl[140] bl[139] bl[138] bl[137] bl[136] bl[135] bl[134] bl[133] bl[132] bl[131] bl[130] bl[129] bl[128] bl[127] bl[126] bl[125] bl[124] bl[123] bl[122] bl[121] bl[120] bl[119] bl[118] bl[117] bl[116] bl[115] bl[114] bl[113] bl[112] bl[111] bl[110] bl[109] bl[108] bl[107] bl[106] bl[105] bl[104] bl[103] bl[102] bl[101] bl[100] bl[99] bl[98] bl[97] bl[96] bl[95] bl[94] bl[93] bl[92] bl[91] bl[90] bl[89] bl[88] bl[87] bl[86] bl[85] bl[84] bl[83] bl[82] bl[81] bl[80] bl[79] bl[78] bl[77] bl[76] bl[75] bl[74] bl[73] bl[72] bl[71] bl[70] bl[69] bl[68] bl[67] bl[66] bl[65] bl[64] bl[63] bl[62] bl[61] bl[60] bl[59] bl[58] bl[57] bl[56] bl[55] bl[54] bl[53] bl[52] bl[51] bl[50] bl[49] bl[48] bl[47] bl[46] bl[45] bl[44] bl[43] bl[42] bl[41] bl[40] bl[39] bl[38] bl[37] bl[36] bl[35] bl[34] bl[33] bl[32] bl[31] bl[30] bl[29] bl[28] bl[27] bl[26] bl[25] bl[24] bl[23] bl[22] bl[21] bl[20] bl[19] bl[18] bl[17] bl[16] bl[15] bl[14] bl[13] bl[12] bl[11] bl[10] bl[9] bl[8] bl[7] bl[6] bl[5] bl[4] bl[3] bl[2] bl[1] bl[0] br[255] br[254] br[253] br[252] br[251] br[250] br[249] br[248] br[247] br[246] br[245] br[244] br[243] br[242] br[241] br[240] br[239] br[238] br[237] br[236] br[235] br[234] br[233] br[232] br[231] br[230] br[229] br[228] br[227] br[226] br[225] br[224] br[223] br[222] br[221] br[220] br[219] br[218] br[217] br[216] br[215] br[214] br[213] br[212] br[211] br[210] br[209] br[208] br[207] br[206] br[205] br[204] br[203] br[202] br[201] br[200] br[199] br[198] br[197] br[196] br[195] br[194] br[193] br[192] br[191] br[190] br[189] br[188] br[187] br[186] br[185] br[184] br[183] br[182] br[181] br[180] br[179] br[178] br[177] br[176] br[175] br[174] br[173] br[172] br[171] br[170] br[169] br[168] br[167] br[166] br[165] br[164] br[163] br[162] br[161] br[160] br[159] br[158] br[157] br[156] br[155] br[154] br[153] br[152] br[151] br[150] br[149] br[148] br[147] br[146] br[145] br[144] br[143] br[142] br[141] br[140] br[139] br[138] br[137] br[136] br[135] br[134] br[133] br[132] br[131] br[130] br[129] br[128] br[127] br[126] br[125] br[124] br[123] br[122] br[121] br[120] br[119] br[118] br[117] br[116] br[115] br[114] br[113] br[112] br[111] br[110] br[109] br[108] br[107] br[106] br[105] br[104] br[103] br[102] br[101] br[100] br[99] br[98] br[97] br[96] br[95] br[94] br[93] br[92] br[91] br[90] br[89] br[88] br[87] br[86] br[85] br[84] br[83] br[82] br[81] br[80] br[79] br[78] br[77] br[76] br[75] br[74] br[73] br[72] br[71] br[70] br[69] br[68] br[67] br[66] br[65] br[64] br[63] br[62] br[61] br[60] br[59] br[58] br[57] br[56] br[55] br[54] br[53] br[52] br[51] br[50] br[49] br[48] br[47] br[46] br[45] br[44] br[43] br[42] br[41] br[40] br[39] br[38] br[37] br[36] br[35] br[34] br[33] br[32] br[31] br[30] br[29] br[28] br[27] br[26] br[25] br[24] br[23] br[22] br[21] br[20] br[19] br[18] br[17] br[16] br[15] br[14] br[13] br[12] br[11] br[10] br[9] br[8] br[7] br[6] br[5] br[4] br[3] br[2] br[1] br[0] bl_out[31] bl_out[30] bl_out[29] bl_out[28] bl_out[27] bl_out[26] bl_out[25] bl_out[24] bl_out[23] bl_out[22] bl_out[21] bl_out[20] bl_out[19] bl_out[18] bl_out[17] bl_out[16] bl_out[15] bl_out[14] bl_out[13] bl_out[12] bl_out[11] bl_out[10] bl_out[9] bl_out[8] bl_out[7] bl_out[6] bl_out[5] bl_out[4] bl_out[3] bl_out[2] bl_out[1] bl_out[0] br_out[31] br_out[30] br_out[29] br_out[28] br_out[27] br_out[26] br_out[25] br_out[24] br_out[23] br_out[22] br_out[21] br_out[20] br_out[19] br_out[18] br_out[17] br_out[16] br_out[15] br_out[14] br_out[13] br_out[12] br_out[11] br_out[10] br_out[9] br_out[8] br_out[7] br_out[6] br_out[5] br_out[4] br_out[3] br_out[2] br_out[1] br_out[0] vdd 

xmux_0 
+ sel_b[0] bl[0] br[0] bl_out[0] br_out[0] vdd 
+ read_mux 
* No parameters

xmux_1 
+ sel_b[1] bl[1] br[1] bl_out[0] br_out[0] vdd 
+ read_mux 
* No parameters

xmux_2 
+ sel_b[2] bl[2] br[2] bl_out[0] br_out[0] vdd 
+ read_mux 
* No parameters

xmux_3 
+ sel_b[3] bl[3] br[3] bl_out[0] br_out[0] vdd 
+ read_mux 
* No parameters

xmux_4 
+ sel_b[4] bl[4] br[4] bl_out[0] br_out[0] vdd 
+ read_mux 
* No parameters

xmux_5 
+ sel_b[5] bl[5] br[5] bl_out[0] br_out[0] vdd 
+ read_mux 
* No parameters

xmux_6 
+ sel_b[6] bl[6] br[6] bl_out[0] br_out[0] vdd 
+ read_mux 
* No parameters

xmux_7 
+ sel_b[7] bl[7] br[7] bl_out[0] br_out[0] vdd 
+ read_mux 
* No parameters

xmux_8 
+ sel_b[0] bl[8] br[8] bl_out[1] br_out[1] vdd 
+ read_mux 
* No parameters

xmux_9 
+ sel_b[1] bl[9] br[9] bl_out[1] br_out[1] vdd 
+ read_mux 
* No parameters

xmux_10 
+ sel_b[2] bl[10] br[10] bl_out[1] br_out[1] vdd 
+ read_mux 
* No parameters

xmux_11 
+ sel_b[3] bl[11] br[11] bl_out[1] br_out[1] vdd 
+ read_mux 
* No parameters

xmux_12 
+ sel_b[4] bl[12] br[12] bl_out[1] br_out[1] vdd 
+ read_mux 
* No parameters

xmux_13 
+ sel_b[5] bl[13] br[13] bl_out[1] br_out[1] vdd 
+ read_mux 
* No parameters

xmux_14 
+ sel_b[6] bl[14] br[14] bl_out[1] br_out[1] vdd 
+ read_mux 
* No parameters

xmux_15 
+ sel_b[7] bl[15] br[15] bl_out[1] br_out[1] vdd 
+ read_mux 
* No parameters

xmux_16 
+ sel_b[0] bl[16] br[16] bl_out[2] br_out[2] vdd 
+ read_mux 
* No parameters

xmux_17 
+ sel_b[1] bl[17] br[17] bl_out[2] br_out[2] vdd 
+ read_mux 
* No parameters

xmux_18 
+ sel_b[2] bl[18] br[18] bl_out[2] br_out[2] vdd 
+ read_mux 
* No parameters

xmux_19 
+ sel_b[3] bl[19] br[19] bl_out[2] br_out[2] vdd 
+ read_mux 
* No parameters

xmux_20 
+ sel_b[4] bl[20] br[20] bl_out[2] br_out[2] vdd 
+ read_mux 
* No parameters

xmux_21 
+ sel_b[5] bl[21] br[21] bl_out[2] br_out[2] vdd 
+ read_mux 
* No parameters

xmux_22 
+ sel_b[6] bl[22] br[22] bl_out[2] br_out[2] vdd 
+ read_mux 
* No parameters

xmux_23 
+ sel_b[7] bl[23] br[23] bl_out[2] br_out[2] vdd 
+ read_mux 
* No parameters

xmux_24 
+ sel_b[0] bl[24] br[24] bl_out[3] br_out[3] vdd 
+ read_mux 
* No parameters

xmux_25 
+ sel_b[1] bl[25] br[25] bl_out[3] br_out[3] vdd 
+ read_mux 
* No parameters

xmux_26 
+ sel_b[2] bl[26] br[26] bl_out[3] br_out[3] vdd 
+ read_mux 
* No parameters

xmux_27 
+ sel_b[3] bl[27] br[27] bl_out[3] br_out[3] vdd 
+ read_mux 
* No parameters

xmux_28 
+ sel_b[4] bl[28] br[28] bl_out[3] br_out[3] vdd 
+ read_mux 
* No parameters

xmux_29 
+ sel_b[5] bl[29] br[29] bl_out[3] br_out[3] vdd 
+ read_mux 
* No parameters

xmux_30 
+ sel_b[6] bl[30] br[30] bl_out[3] br_out[3] vdd 
+ read_mux 
* No parameters

xmux_31 
+ sel_b[7] bl[31] br[31] bl_out[3] br_out[3] vdd 
+ read_mux 
* No parameters

xmux_32 
+ sel_b[0] bl[32] br[32] bl_out[4] br_out[4] vdd 
+ read_mux 
* No parameters

xmux_33 
+ sel_b[1] bl[33] br[33] bl_out[4] br_out[4] vdd 
+ read_mux 
* No parameters

xmux_34 
+ sel_b[2] bl[34] br[34] bl_out[4] br_out[4] vdd 
+ read_mux 
* No parameters

xmux_35 
+ sel_b[3] bl[35] br[35] bl_out[4] br_out[4] vdd 
+ read_mux 
* No parameters

xmux_36 
+ sel_b[4] bl[36] br[36] bl_out[4] br_out[4] vdd 
+ read_mux 
* No parameters

xmux_37 
+ sel_b[5] bl[37] br[37] bl_out[4] br_out[4] vdd 
+ read_mux 
* No parameters

xmux_38 
+ sel_b[6] bl[38] br[38] bl_out[4] br_out[4] vdd 
+ read_mux 
* No parameters

xmux_39 
+ sel_b[7] bl[39] br[39] bl_out[4] br_out[4] vdd 
+ read_mux 
* No parameters

xmux_40 
+ sel_b[0] bl[40] br[40] bl_out[5] br_out[5] vdd 
+ read_mux 
* No parameters

xmux_41 
+ sel_b[1] bl[41] br[41] bl_out[5] br_out[5] vdd 
+ read_mux 
* No parameters

xmux_42 
+ sel_b[2] bl[42] br[42] bl_out[5] br_out[5] vdd 
+ read_mux 
* No parameters

xmux_43 
+ sel_b[3] bl[43] br[43] bl_out[5] br_out[5] vdd 
+ read_mux 
* No parameters

xmux_44 
+ sel_b[4] bl[44] br[44] bl_out[5] br_out[5] vdd 
+ read_mux 
* No parameters

xmux_45 
+ sel_b[5] bl[45] br[45] bl_out[5] br_out[5] vdd 
+ read_mux 
* No parameters

xmux_46 
+ sel_b[6] bl[46] br[46] bl_out[5] br_out[5] vdd 
+ read_mux 
* No parameters

xmux_47 
+ sel_b[7] bl[47] br[47] bl_out[5] br_out[5] vdd 
+ read_mux 
* No parameters

xmux_48 
+ sel_b[0] bl[48] br[48] bl_out[6] br_out[6] vdd 
+ read_mux 
* No parameters

xmux_49 
+ sel_b[1] bl[49] br[49] bl_out[6] br_out[6] vdd 
+ read_mux 
* No parameters

xmux_50 
+ sel_b[2] bl[50] br[50] bl_out[6] br_out[6] vdd 
+ read_mux 
* No parameters

xmux_51 
+ sel_b[3] bl[51] br[51] bl_out[6] br_out[6] vdd 
+ read_mux 
* No parameters

xmux_52 
+ sel_b[4] bl[52] br[52] bl_out[6] br_out[6] vdd 
+ read_mux 
* No parameters

xmux_53 
+ sel_b[5] bl[53] br[53] bl_out[6] br_out[6] vdd 
+ read_mux 
* No parameters

xmux_54 
+ sel_b[6] bl[54] br[54] bl_out[6] br_out[6] vdd 
+ read_mux 
* No parameters

xmux_55 
+ sel_b[7] bl[55] br[55] bl_out[6] br_out[6] vdd 
+ read_mux 
* No parameters

xmux_56 
+ sel_b[0] bl[56] br[56] bl_out[7] br_out[7] vdd 
+ read_mux 
* No parameters

xmux_57 
+ sel_b[1] bl[57] br[57] bl_out[7] br_out[7] vdd 
+ read_mux 
* No parameters

xmux_58 
+ sel_b[2] bl[58] br[58] bl_out[7] br_out[7] vdd 
+ read_mux 
* No parameters

xmux_59 
+ sel_b[3] bl[59] br[59] bl_out[7] br_out[7] vdd 
+ read_mux 
* No parameters

xmux_60 
+ sel_b[4] bl[60] br[60] bl_out[7] br_out[7] vdd 
+ read_mux 
* No parameters

xmux_61 
+ sel_b[5] bl[61] br[61] bl_out[7] br_out[7] vdd 
+ read_mux 
* No parameters

xmux_62 
+ sel_b[6] bl[62] br[62] bl_out[7] br_out[7] vdd 
+ read_mux 
* No parameters

xmux_63 
+ sel_b[7] bl[63] br[63] bl_out[7] br_out[7] vdd 
+ read_mux 
* No parameters

xmux_64 
+ sel_b[0] bl[64] br[64] bl_out[8] br_out[8] vdd 
+ read_mux 
* No parameters

xmux_65 
+ sel_b[1] bl[65] br[65] bl_out[8] br_out[8] vdd 
+ read_mux 
* No parameters

xmux_66 
+ sel_b[2] bl[66] br[66] bl_out[8] br_out[8] vdd 
+ read_mux 
* No parameters

xmux_67 
+ sel_b[3] bl[67] br[67] bl_out[8] br_out[8] vdd 
+ read_mux 
* No parameters

xmux_68 
+ sel_b[4] bl[68] br[68] bl_out[8] br_out[8] vdd 
+ read_mux 
* No parameters

xmux_69 
+ sel_b[5] bl[69] br[69] bl_out[8] br_out[8] vdd 
+ read_mux 
* No parameters

xmux_70 
+ sel_b[6] bl[70] br[70] bl_out[8] br_out[8] vdd 
+ read_mux 
* No parameters

xmux_71 
+ sel_b[7] bl[71] br[71] bl_out[8] br_out[8] vdd 
+ read_mux 
* No parameters

xmux_72 
+ sel_b[0] bl[72] br[72] bl_out[9] br_out[9] vdd 
+ read_mux 
* No parameters

xmux_73 
+ sel_b[1] bl[73] br[73] bl_out[9] br_out[9] vdd 
+ read_mux 
* No parameters

xmux_74 
+ sel_b[2] bl[74] br[74] bl_out[9] br_out[9] vdd 
+ read_mux 
* No parameters

xmux_75 
+ sel_b[3] bl[75] br[75] bl_out[9] br_out[9] vdd 
+ read_mux 
* No parameters

xmux_76 
+ sel_b[4] bl[76] br[76] bl_out[9] br_out[9] vdd 
+ read_mux 
* No parameters

xmux_77 
+ sel_b[5] bl[77] br[77] bl_out[9] br_out[9] vdd 
+ read_mux 
* No parameters

xmux_78 
+ sel_b[6] bl[78] br[78] bl_out[9] br_out[9] vdd 
+ read_mux 
* No parameters

xmux_79 
+ sel_b[7] bl[79] br[79] bl_out[9] br_out[9] vdd 
+ read_mux 
* No parameters

xmux_80 
+ sel_b[0] bl[80] br[80] bl_out[10] br_out[10] vdd 
+ read_mux 
* No parameters

xmux_81 
+ sel_b[1] bl[81] br[81] bl_out[10] br_out[10] vdd 
+ read_mux 
* No parameters

xmux_82 
+ sel_b[2] bl[82] br[82] bl_out[10] br_out[10] vdd 
+ read_mux 
* No parameters

xmux_83 
+ sel_b[3] bl[83] br[83] bl_out[10] br_out[10] vdd 
+ read_mux 
* No parameters

xmux_84 
+ sel_b[4] bl[84] br[84] bl_out[10] br_out[10] vdd 
+ read_mux 
* No parameters

xmux_85 
+ sel_b[5] bl[85] br[85] bl_out[10] br_out[10] vdd 
+ read_mux 
* No parameters

xmux_86 
+ sel_b[6] bl[86] br[86] bl_out[10] br_out[10] vdd 
+ read_mux 
* No parameters

xmux_87 
+ sel_b[7] bl[87] br[87] bl_out[10] br_out[10] vdd 
+ read_mux 
* No parameters

xmux_88 
+ sel_b[0] bl[88] br[88] bl_out[11] br_out[11] vdd 
+ read_mux 
* No parameters

xmux_89 
+ sel_b[1] bl[89] br[89] bl_out[11] br_out[11] vdd 
+ read_mux 
* No parameters

xmux_90 
+ sel_b[2] bl[90] br[90] bl_out[11] br_out[11] vdd 
+ read_mux 
* No parameters

xmux_91 
+ sel_b[3] bl[91] br[91] bl_out[11] br_out[11] vdd 
+ read_mux 
* No parameters

xmux_92 
+ sel_b[4] bl[92] br[92] bl_out[11] br_out[11] vdd 
+ read_mux 
* No parameters

xmux_93 
+ sel_b[5] bl[93] br[93] bl_out[11] br_out[11] vdd 
+ read_mux 
* No parameters

xmux_94 
+ sel_b[6] bl[94] br[94] bl_out[11] br_out[11] vdd 
+ read_mux 
* No parameters

xmux_95 
+ sel_b[7] bl[95] br[95] bl_out[11] br_out[11] vdd 
+ read_mux 
* No parameters

xmux_96 
+ sel_b[0] bl[96] br[96] bl_out[12] br_out[12] vdd 
+ read_mux 
* No parameters

xmux_97 
+ sel_b[1] bl[97] br[97] bl_out[12] br_out[12] vdd 
+ read_mux 
* No parameters

xmux_98 
+ sel_b[2] bl[98] br[98] bl_out[12] br_out[12] vdd 
+ read_mux 
* No parameters

xmux_99 
+ sel_b[3] bl[99] br[99] bl_out[12] br_out[12] vdd 
+ read_mux 
* No parameters

xmux_100 
+ sel_b[4] bl[100] br[100] bl_out[12] br_out[12] vdd 
+ read_mux 
* No parameters

xmux_101 
+ sel_b[5] bl[101] br[101] bl_out[12] br_out[12] vdd 
+ read_mux 
* No parameters

xmux_102 
+ sel_b[6] bl[102] br[102] bl_out[12] br_out[12] vdd 
+ read_mux 
* No parameters

xmux_103 
+ sel_b[7] bl[103] br[103] bl_out[12] br_out[12] vdd 
+ read_mux 
* No parameters

xmux_104 
+ sel_b[0] bl[104] br[104] bl_out[13] br_out[13] vdd 
+ read_mux 
* No parameters

xmux_105 
+ sel_b[1] bl[105] br[105] bl_out[13] br_out[13] vdd 
+ read_mux 
* No parameters

xmux_106 
+ sel_b[2] bl[106] br[106] bl_out[13] br_out[13] vdd 
+ read_mux 
* No parameters

xmux_107 
+ sel_b[3] bl[107] br[107] bl_out[13] br_out[13] vdd 
+ read_mux 
* No parameters

xmux_108 
+ sel_b[4] bl[108] br[108] bl_out[13] br_out[13] vdd 
+ read_mux 
* No parameters

xmux_109 
+ sel_b[5] bl[109] br[109] bl_out[13] br_out[13] vdd 
+ read_mux 
* No parameters

xmux_110 
+ sel_b[6] bl[110] br[110] bl_out[13] br_out[13] vdd 
+ read_mux 
* No parameters

xmux_111 
+ sel_b[7] bl[111] br[111] bl_out[13] br_out[13] vdd 
+ read_mux 
* No parameters

xmux_112 
+ sel_b[0] bl[112] br[112] bl_out[14] br_out[14] vdd 
+ read_mux 
* No parameters

xmux_113 
+ sel_b[1] bl[113] br[113] bl_out[14] br_out[14] vdd 
+ read_mux 
* No parameters

xmux_114 
+ sel_b[2] bl[114] br[114] bl_out[14] br_out[14] vdd 
+ read_mux 
* No parameters

xmux_115 
+ sel_b[3] bl[115] br[115] bl_out[14] br_out[14] vdd 
+ read_mux 
* No parameters

xmux_116 
+ sel_b[4] bl[116] br[116] bl_out[14] br_out[14] vdd 
+ read_mux 
* No parameters

xmux_117 
+ sel_b[5] bl[117] br[117] bl_out[14] br_out[14] vdd 
+ read_mux 
* No parameters

xmux_118 
+ sel_b[6] bl[118] br[118] bl_out[14] br_out[14] vdd 
+ read_mux 
* No parameters

xmux_119 
+ sel_b[7] bl[119] br[119] bl_out[14] br_out[14] vdd 
+ read_mux 
* No parameters

xmux_120 
+ sel_b[0] bl[120] br[120] bl_out[15] br_out[15] vdd 
+ read_mux 
* No parameters

xmux_121 
+ sel_b[1] bl[121] br[121] bl_out[15] br_out[15] vdd 
+ read_mux 
* No parameters

xmux_122 
+ sel_b[2] bl[122] br[122] bl_out[15] br_out[15] vdd 
+ read_mux 
* No parameters

xmux_123 
+ sel_b[3] bl[123] br[123] bl_out[15] br_out[15] vdd 
+ read_mux 
* No parameters

xmux_124 
+ sel_b[4] bl[124] br[124] bl_out[15] br_out[15] vdd 
+ read_mux 
* No parameters

xmux_125 
+ sel_b[5] bl[125] br[125] bl_out[15] br_out[15] vdd 
+ read_mux 
* No parameters

xmux_126 
+ sel_b[6] bl[126] br[126] bl_out[15] br_out[15] vdd 
+ read_mux 
* No parameters

xmux_127 
+ sel_b[7] bl[127] br[127] bl_out[15] br_out[15] vdd 
+ read_mux 
* No parameters

xmux_128 
+ sel_b[0] bl[128] br[128] bl_out[16] br_out[16] vdd 
+ read_mux 
* No parameters

xmux_129 
+ sel_b[1] bl[129] br[129] bl_out[16] br_out[16] vdd 
+ read_mux 
* No parameters

xmux_130 
+ sel_b[2] bl[130] br[130] bl_out[16] br_out[16] vdd 
+ read_mux 
* No parameters

xmux_131 
+ sel_b[3] bl[131] br[131] bl_out[16] br_out[16] vdd 
+ read_mux 
* No parameters

xmux_132 
+ sel_b[4] bl[132] br[132] bl_out[16] br_out[16] vdd 
+ read_mux 
* No parameters

xmux_133 
+ sel_b[5] bl[133] br[133] bl_out[16] br_out[16] vdd 
+ read_mux 
* No parameters

xmux_134 
+ sel_b[6] bl[134] br[134] bl_out[16] br_out[16] vdd 
+ read_mux 
* No parameters

xmux_135 
+ sel_b[7] bl[135] br[135] bl_out[16] br_out[16] vdd 
+ read_mux 
* No parameters

xmux_136 
+ sel_b[0] bl[136] br[136] bl_out[17] br_out[17] vdd 
+ read_mux 
* No parameters

xmux_137 
+ sel_b[1] bl[137] br[137] bl_out[17] br_out[17] vdd 
+ read_mux 
* No parameters

xmux_138 
+ sel_b[2] bl[138] br[138] bl_out[17] br_out[17] vdd 
+ read_mux 
* No parameters

xmux_139 
+ sel_b[3] bl[139] br[139] bl_out[17] br_out[17] vdd 
+ read_mux 
* No parameters

xmux_140 
+ sel_b[4] bl[140] br[140] bl_out[17] br_out[17] vdd 
+ read_mux 
* No parameters

xmux_141 
+ sel_b[5] bl[141] br[141] bl_out[17] br_out[17] vdd 
+ read_mux 
* No parameters

xmux_142 
+ sel_b[6] bl[142] br[142] bl_out[17] br_out[17] vdd 
+ read_mux 
* No parameters

xmux_143 
+ sel_b[7] bl[143] br[143] bl_out[17] br_out[17] vdd 
+ read_mux 
* No parameters

xmux_144 
+ sel_b[0] bl[144] br[144] bl_out[18] br_out[18] vdd 
+ read_mux 
* No parameters

xmux_145 
+ sel_b[1] bl[145] br[145] bl_out[18] br_out[18] vdd 
+ read_mux 
* No parameters

xmux_146 
+ sel_b[2] bl[146] br[146] bl_out[18] br_out[18] vdd 
+ read_mux 
* No parameters

xmux_147 
+ sel_b[3] bl[147] br[147] bl_out[18] br_out[18] vdd 
+ read_mux 
* No parameters

xmux_148 
+ sel_b[4] bl[148] br[148] bl_out[18] br_out[18] vdd 
+ read_mux 
* No parameters

xmux_149 
+ sel_b[5] bl[149] br[149] bl_out[18] br_out[18] vdd 
+ read_mux 
* No parameters

xmux_150 
+ sel_b[6] bl[150] br[150] bl_out[18] br_out[18] vdd 
+ read_mux 
* No parameters

xmux_151 
+ sel_b[7] bl[151] br[151] bl_out[18] br_out[18] vdd 
+ read_mux 
* No parameters

xmux_152 
+ sel_b[0] bl[152] br[152] bl_out[19] br_out[19] vdd 
+ read_mux 
* No parameters

xmux_153 
+ sel_b[1] bl[153] br[153] bl_out[19] br_out[19] vdd 
+ read_mux 
* No parameters

xmux_154 
+ sel_b[2] bl[154] br[154] bl_out[19] br_out[19] vdd 
+ read_mux 
* No parameters

xmux_155 
+ sel_b[3] bl[155] br[155] bl_out[19] br_out[19] vdd 
+ read_mux 
* No parameters

xmux_156 
+ sel_b[4] bl[156] br[156] bl_out[19] br_out[19] vdd 
+ read_mux 
* No parameters

xmux_157 
+ sel_b[5] bl[157] br[157] bl_out[19] br_out[19] vdd 
+ read_mux 
* No parameters

xmux_158 
+ sel_b[6] bl[158] br[158] bl_out[19] br_out[19] vdd 
+ read_mux 
* No parameters

xmux_159 
+ sel_b[7] bl[159] br[159] bl_out[19] br_out[19] vdd 
+ read_mux 
* No parameters

xmux_160 
+ sel_b[0] bl[160] br[160] bl_out[20] br_out[20] vdd 
+ read_mux 
* No parameters

xmux_161 
+ sel_b[1] bl[161] br[161] bl_out[20] br_out[20] vdd 
+ read_mux 
* No parameters

xmux_162 
+ sel_b[2] bl[162] br[162] bl_out[20] br_out[20] vdd 
+ read_mux 
* No parameters

xmux_163 
+ sel_b[3] bl[163] br[163] bl_out[20] br_out[20] vdd 
+ read_mux 
* No parameters

xmux_164 
+ sel_b[4] bl[164] br[164] bl_out[20] br_out[20] vdd 
+ read_mux 
* No parameters

xmux_165 
+ sel_b[5] bl[165] br[165] bl_out[20] br_out[20] vdd 
+ read_mux 
* No parameters

xmux_166 
+ sel_b[6] bl[166] br[166] bl_out[20] br_out[20] vdd 
+ read_mux 
* No parameters

xmux_167 
+ sel_b[7] bl[167] br[167] bl_out[20] br_out[20] vdd 
+ read_mux 
* No parameters

xmux_168 
+ sel_b[0] bl[168] br[168] bl_out[21] br_out[21] vdd 
+ read_mux 
* No parameters

xmux_169 
+ sel_b[1] bl[169] br[169] bl_out[21] br_out[21] vdd 
+ read_mux 
* No parameters

xmux_170 
+ sel_b[2] bl[170] br[170] bl_out[21] br_out[21] vdd 
+ read_mux 
* No parameters

xmux_171 
+ sel_b[3] bl[171] br[171] bl_out[21] br_out[21] vdd 
+ read_mux 
* No parameters

xmux_172 
+ sel_b[4] bl[172] br[172] bl_out[21] br_out[21] vdd 
+ read_mux 
* No parameters

xmux_173 
+ sel_b[5] bl[173] br[173] bl_out[21] br_out[21] vdd 
+ read_mux 
* No parameters

xmux_174 
+ sel_b[6] bl[174] br[174] bl_out[21] br_out[21] vdd 
+ read_mux 
* No parameters

xmux_175 
+ sel_b[7] bl[175] br[175] bl_out[21] br_out[21] vdd 
+ read_mux 
* No parameters

xmux_176 
+ sel_b[0] bl[176] br[176] bl_out[22] br_out[22] vdd 
+ read_mux 
* No parameters

xmux_177 
+ sel_b[1] bl[177] br[177] bl_out[22] br_out[22] vdd 
+ read_mux 
* No parameters

xmux_178 
+ sel_b[2] bl[178] br[178] bl_out[22] br_out[22] vdd 
+ read_mux 
* No parameters

xmux_179 
+ sel_b[3] bl[179] br[179] bl_out[22] br_out[22] vdd 
+ read_mux 
* No parameters

xmux_180 
+ sel_b[4] bl[180] br[180] bl_out[22] br_out[22] vdd 
+ read_mux 
* No parameters

xmux_181 
+ sel_b[5] bl[181] br[181] bl_out[22] br_out[22] vdd 
+ read_mux 
* No parameters

xmux_182 
+ sel_b[6] bl[182] br[182] bl_out[22] br_out[22] vdd 
+ read_mux 
* No parameters

xmux_183 
+ sel_b[7] bl[183] br[183] bl_out[22] br_out[22] vdd 
+ read_mux 
* No parameters

xmux_184 
+ sel_b[0] bl[184] br[184] bl_out[23] br_out[23] vdd 
+ read_mux 
* No parameters

xmux_185 
+ sel_b[1] bl[185] br[185] bl_out[23] br_out[23] vdd 
+ read_mux 
* No parameters

xmux_186 
+ sel_b[2] bl[186] br[186] bl_out[23] br_out[23] vdd 
+ read_mux 
* No parameters

xmux_187 
+ sel_b[3] bl[187] br[187] bl_out[23] br_out[23] vdd 
+ read_mux 
* No parameters

xmux_188 
+ sel_b[4] bl[188] br[188] bl_out[23] br_out[23] vdd 
+ read_mux 
* No parameters

xmux_189 
+ sel_b[5] bl[189] br[189] bl_out[23] br_out[23] vdd 
+ read_mux 
* No parameters

xmux_190 
+ sel_b[6] bl[190] br[190] bl_out[23] br_out[23] vdd 
+ read_mux 
* No parameters

xmux_191 
+ sel_b[7] bl[191] br[191] bl_out[23] br_out[23] vdd 
+ read_mux 
* No parameters

xmux_192 
+ sel_b[0] bl[192] br[192] bl_out[24] br_out[24] vdd 
+ read_mux 
* No parameters

xmux_193 
+ sel_b[1] bl[193] br[193] bl_out[24] br_out[24] vdd 
+ read_mux 
* No parameters

xmux_194 
+ sel_b[2] bl[194] br[194] bl_out[24] br_out[24] vdd 
+ read_mux 
* No parameters

xmux_195 
+ sel_b[3] bl[195] br[195] bl_out[24] br_out[24] vdd 
+ read_mux 
* No parameters

xmux_196 
+ sel_b[4] bl[196] br[196] bl_out[24] br_out[24] vdd 
+ read_mux 
* No parameters

xmux_197 
+ sel_b[5] bl[197] br[197] bl_out[24] br_out[24] vdd 
+ read_mux 
* No parameters

xmux_198 
+ sel_b[6] bl[198] br[198] bl_out[24] br_out[24] vdd 
+ read_mux 
* No parameters

xmux_199 
+ sel_b[7] bl[199] br[199] bl_out[24] br_out[24] vdd 
+ read_mux 
* No parameters

xmux_200 
+ sel_b[0] bl[200] br[200] bl_out[25] br_out[25] vdd 
+ read_mux 
* No parameters

xmux_201 
+ sel_b[1] bl[201] br[201] bl_out[25] br_out[25] vdd 
+ read_mux 
* No parameters

xmux_202 
+ sel_b[2] bl[202] br[202] bl_out[25] br_out[25] vdd 
+ read_mux 
* No parameters

xmux_203 
+ sel_b[3] bl[203] br[203] bl_out[25] br_out[25] vdd 
+ read_mux 
* No parameters

xmux_204 
+ sel_b[4] bl[204] br[204] bl_out[25] br_out[25] vdd 
+ read_mux 
* No parameters

xmux_205 
+ sel_b[5] bl[205] br[205] bl_out[25] br_out[25] vdd 
+ read_mux 
* No parameters

xmux_206 
+ sel_b[6] bl[206] br[206] bl_out[25] br_out[25] vdd 
+ read_mux 
* No parameters

xmux_207 
+ sel_b[7] bl[207] br[207] bl_out[25] br_out[25] vdd 
+ read_mux 
* No parameters

xmux_208 
+ sel_b[0] bl[208] br[208] bl_out[26] br_out[26] vdd 
+ read_mux 
* No parameters

xmux_209 
+ sel_b[1] bl[209] br[209] bl_out[26] br_out[26] vdd 
+ read_mux 
* No parameters

xmux_210 
+ sel_b[2] bl[210] br[210] bl_out[26] br_out[26] vdd 
+ read_mux 
* No parameters

xmux_211 
+ sel_b[3] bl[211] br[211] bl_out[26] br_out[26] vdd 
+ read_mux 
* No parameters

xmux_212 
+ sel_b[4] bl[212] br[212] bl_out[26] br_out[26] vdd 
+ read_mux 
* No parameters

xmux_213 
+ sel_b[5] bl[213] br[213] bl_out[26] br_out[26] vdd 
+ read_mux 
* No parameters

xmux_214 
+ sel_b[6] bl[214] br[214] bl_out[26] br_out[26] vdd 
+ read_mux 
* No parameters

xmux_215 
+ sel_b[7] bl[215] br[215] bl_out[26] br_out[26] vdd 
+ read_mux 
* No parameters

xmux_216 
+ sel_b[0] bl[216] br[216] bl_out[27] br_out[27] vdd 
+ read_mux 
* No parameters

xmux_217 
+ sel_b[1] bl[217] br[217] bl_out[27] br_out[27] vdd 
+ read_mux 
* No parameters

xmux_218 
+ sel_b[2] bl[218] br[218] bl_out[27] br_out[27] vdd 
+ read_mux 
* No parameters

xmux_219 
+ sel_b[3] bl[219] br[219] bl_out[27] br_out[27] vdd 
+ read_mux 
* No parameters

xmux_220 
+ sel_b[4] bl[220] br[220] bl_out[27] br_out[27] vdd 
+ read_mux 
* No parameters

xmux_221 
+ sel_b[5] bl[221] br[221] bl_out[27] br_out[27] vdd 
+ read_mux 
* No parameters

xmux_222 
+ sel_b[6] bl[222] br[222] bl_out[27] br_out[27] vdd 
+ read_mux 
* No parameters

xmux_223 
+ sel_b[7] bl[223] br[223] bl_out[27] br_out[27] vdd 
+ read_mux 
* No parameters

xmux_224 
+ sel_b[0] bl[224] br[224] bl_out[28] br_out[28] vdd 
+ read_mux 
* No parameters

xmux_225 
+ sel_b[1] bl[225] br[225] bl_out[28] br_out[28] vdd 
+ read_mux 
* No parameters

xmux_226 
+ sel_b[2] bl[226] br[226] bl_out[28] br_out[28] vdd 
+ read_mux 
* No parameters

xmux_227 
+ sel_b[3] bl[227] br[227] bl_out[28] br_out[28] vdd 
+ read_mux 
* No parameters

xmux_228 
+ sel_b[4] bl[228] br[228] bl_out[28] br_out[28] vdd 
+ read_mux 
* No parameters

xmux_229 
+ sel_b[5] bl[229] br[229] bl_out[28] br_out[28] vdd 
+ read_mux 
* No parameters

xmux_230 
+ sel_b[6] bl[230] br[230] bl_out[28] br_out[28] vdd 
+ read_mux 
* No parameters

xmux_231 
+ sel_b[7] bl[231] br[231] bl_out[28] br_out[28] vdd 
+ read_mux 
* No parameters

xmux_232 
+ sel_b[0] bl[232] br[232] bl_out[29] br_out[29] vdd 
+ read_mux 
* No parameters

xmux_233 
+ sel_b[1] bl[233] br[233] bl_out[29] br_out[29] vdd 
+ read_mux 
* No parameters

xmux_234 
+ sel_b[2] bl[234] br[234] bl_out[29] br_out[29] vdd 
+ read_mux 
* No parameters

xmux_235 
+ sel_b[3] bl[235] br[235] bl_out[29] br_out[29] vdd 
+ read_mux 
* No parameters

xmux_236 
+ sel_b[4] bl[236] br[236] bl_out[29] br_out[29] vdd 
+ read_mux 
* No parameters

xmux_237 
+ sel_b[5] bl[237] br[237] bl_out[29] br_out[29] vdd 
+ read_mux 
* No parameters

xmux_238 
+ sel_b[6] bl[238] br[238] bl_out[29] br_out[29] vdd 
+ read_mux 
* No parameters

xmux_239 
+ sel_b[7] bl[239] br[239] bl_out[29] br_out[29] vdd 
+ read_mux 
* No parameters

xmux_240 
+ sel_b[0] bl[240] br[240] bl_out[30] br_out[30] vdd 
+ read_mux 
* No parameters

xmux_241 
+ sel_b[1] bl[241] br[241] bl_out[30] br_out[30] vdd 
+ read_mux 
* No parameters

xmux_242 
+ sel_b[2] bl[242] br[242] bl_out[30] br_out[30] vdd 
+ read_mux 
* No parameters

xmux_243 
+ sel_b[3] bl[243] br[243] bl_out[30] br_out[30] vdd 
+ read_mux 
* No parameters

xmux_244 
+ sel_b[4] bl[244] br[244] bl_out[30] br_out[30] vdd 
+ read_mux 
* No parameters

xmux_245 
+ sel_b[5] bl[245] br[245] bl_out[30] br_out[30] vdd 
+ read_mux 
* No parameters

xmux_246 
+ sel_b[6] bl[246] br[246] bl_out[30] br_out[30] vdd 
+ read_mux 
* No parameters

xmux_247 
+ sel_b[7] bl[247] br[247] bl_out[30] br_out[30] vdd 
+ read_mux 
* No parameters

xmux_248 
+ sel_b[0] bl[248] br[248] bl_out[31] br_out[31] vdd 
+ read_mux 
* No parameters

xmux_249 
+ sel_b[1] bl[249] br[249] bl_out[31] br_out[31] vdd 
+ read_mux 
* No parameters

xmux_250 
+ sel_b[2] bl[250] br[250] bl_out[31] br_out[31] vdd 
+ read_mux 
* No parameters

xmux_251 
+ sel_b[3] bl[251] br[251] bl_out[31] br_out[31] vdd 
+ read_mux 
* No parameters

xmux_252 
+ sel_b[4] bl[252] br[252] bl_out[31] br_out[31] vdd 
+ read_mux 
* No parameters

xmux_253 
+ sel_b[5] bl[253] br[253] bl_out[31] br_out[31] vdd 
+ read_mux 
* No parameters

xmux_254 
+ sel_b[6] bl[254] br[254] bl_out[31] br_out[31] vdd 
+ read_mux 
* No parameters

xmux_255 
+ sel_b[7] bl[255] br[255] bl_out[31] br_out[31] vdd 
+ read_mux 
* No parameters

.ENDS

.SUBCKT write_mux 
+ we wmask data data_b bl br vss 

xMMUXBR 
+ br data x vss 
+ sky130_fd_pr__nfet_01v8 
+ w='2.0' l='0.15' 

xMMUXBL 
+ bl data_b x vss 
+ sky130_fd_pr__nfet_01v8 
+ w='2.0' l='0.15' 

xMWMASK 
+ x wmask y vss 
+ sky130_fd_pr__nfet_01v8 
+ w='2.0' l='0.15' 

xMPD 
+ y we vss vss 
+ sky130_fd_pr__nfet_01v8 
+ w='2.0' l='0.15' 

.ENDS

.SUBCKT write_mux_array 
+ we[7] we[6] we[5] we[4] we[3] we[2] we[1] we[0] wmask[3] wmask[2] wmask[1] wmask[0] data[31] data[30] data[29] data[28] data[27] data[26] data[25] data[24] data[23] data[22] data[21] data[20] data[19] data[18] data[17] data[16] data[15] data[14] data[13] data[12] data[11] data[10] data[9] data[8] data[7] data[6] data[5] data[4] data[3] data[2] data[1] data[0] data_b[31] data_b[30] data_b[29] data_b[28] data_b[27] data_b[26] data_b[25] data_b[24] data_b[23] data_b[22] data_b[21] data_b[20] data_b[19] data_b[18] data_b[17] data_b[16] data_b[15] data_b[14] data_b[13] data_b[12] data_b[11] data_b[10] data_b[9] data_b[8] data_b[7] data_b[6] data_b[5] data_b[4] data_b[3] data_b[2] data_b[1] data_b[0] bl[255] bl[254] bl[253] bl[252] bl[251] bl[250] bl[249] bl[248] bl[247] bl[246] bl[245] bl[244] bl[243] bl[242] bl[241] bl[240] bl[239] bl[238] bl[237] bl[236] bl[235] bl[234] bl[233] bl[232] bl[231] bl[230] bl[229] bl[228] bl[227] bl[226] bl[225] bl[224] bl[223] bl[222] bl[221] bl[220] bl[219] bl[218] bl[217] bl[216] bl[215] bl[214] bl[213] bl[212] bl[211] bl[210] bl[209] bl[208] bl[207] bl[206] bl[205] bl[204] bl[203] bl[202] bl[201] bl[200] bl[199] bl[198] bl[197] bl[196] bl[195] bl[194] bl[193] bl[192] bl[191] bl[190] bl[189] bl[188] bl[187] bl[186] bl[185] bl[184] bl[183] bl[182] bl[181] bl[180] bl[179] bl[178] bl[177] bl[176] bl[175] bl[174] bl[173] bl[172] bl[171] bl[170] bl[169] bl[168] bl[167] bl[166] bl[165] bl[164] bl[163] bl[162] bl[161] bl[160] bl[159] bl[158] bl[157] bl[156] bl[155] bl[154] bl[153] bl[152] bl[151] bl[150] bl[149] bl[148] bl[147] bl[146] bl[145] bl[144] bl[143] bl[142] bl[141] bl[140] bl[139] bl[138] bl[137] bl[136] bl[135] bl[134] bl[133] bl[132] bl[131] bl[130] bl[129] bl[128] bl[127] bl[126] bl[125] bl[124] bl[123] bl[122] bl[121] bl[120] bl[119] bl[118] bl[117] bl[116] bl[115] bl[114] bl[113] bl[112] bl[111] bl[110] bl[109] bl[108] bl[107] bl[106] bl[105] bl[104] bl[103] bl[102] bl[101] bl[100] bl[99] bl[98] bl[97] bl[96] bl[95] bl[94] bl[93] bl[92] bl[91] bl[90] bl[89] bl[88] bl[87] bl[86] bl[85] bl[84] bl[83] bl[82] bl[81] bl[80] bl[79] bl[78] bl[77] bl[76] bl[75] bl[74] bl[73] bl[72] bl[71] bl[70] bl[69] bl[68] bl[67] bl[66] bl[65] bl[64] bl[63] bl[62] bl[61] bl[60] bl[59] bl[58] bl[57] bl[56] bl[55] bl[54] bl[53] bl[52] bl[51] bl[50] bl[49] bl[48] bl[47] bl[46] bl[45] bl[44] bl[43] bl[42] bl[41] bl[40] bl[39] bl[38] bl[37] bl[36] bl[35] bl[34] bl[33] bl[32] bl[31] bl[30] bl[29] bl[28] bl[27] bl[26] bl[25] bl[24] bl[23] bl[22] bl[21] bl[20] bl[19] bl[18] bl[17] bl[16] bl[15] bl[14] bl[13] bl[12] bl[11] bl[10] bl[9] bl[8] bl[7] bl[6] bl[5] bl[4] bl[3] bl[2] bl[1] bl[0] br[255] br[254] br[253] br[252] br[251] br[250] br[249] br[248] br[247] br[246] br[245] br[244] br[243] br[242] br[241] br[240] br[239] br[238] br[237] br[236] br[235] br[234] br[233] br[232] br[231] br[230] br[229] br[228] br[227] br[226] br[225] br[224] br[223] br[222] br[221] br[220] br[219] br[218] br[217] br[216] br[215] br[214] br[213] br[212] br[211] br[210] br[209] br[208] br[207] br[206] br[205] br[204] br[203] br[202] br[201] br[200] br[199] br[198] br[197] br[196] br[195] br[194] br[193] br[192] br[191] br[190] br[189] br[188] br[187] br[186] br[185] br[184] br[183] br[182] br[181] br[180] br[179] br[178] br[177] br[176] br[175] br[174] br[173] br[172] br[171] br[170] br[169] br[168] br[167] br[166] br[165] br[164] br[163] br[162] br[161] br[160] br[159] br[158] br[157] br[156] br[155] br[154] br[153] br[152] br[151] br[150] br[149] br[148] br[147] br[146] br[145] br[144] br[143] br[142] br[141] br[140] br[139] br[138] br[137] br[136] br[135] br[134] br[133] br[132] br[131] br[130] br[129] br[128] br[127] br[126] br[125] br[124] br[123] br[122] br[121] br[120] br[119] br[118] br[117] br[116] br[115] br[114] br[113] br[112] br[111] br[110] br[109] br[108] br[107] br[106] br[105] br[104] br[103] br[102] br[101] br[100] br[99] br[98] br[97] br[96] br[95] br[94] br[93] br[92] br[91] br[90] br[89] br[88] br[87] br[86] br[85] br[84] br[83] br[82] br[81] br[80] br[79] br[78] br[77] br[76] br[75] br[74] br[73] br[72] br[71] br[70] br[69] br[68] br[67] br[66] br[65] br[64] br[63] br[62] br[61] br[60] br[59] br[58] br[57] br[56] br[55] br[54] br[53] br[52] br[51] br[50] br[49] br[48] br[47] br[46] br[45] br[44] br[43] br[42] br[41] br[40] br[39] br[38] br[37] br[36] br[35] br[34] br[33] br[32] br[31] br[30] br[29] br[28] br[27] br[26] br[25] br[24] br[23] br[22] br[21] br[20] br[19] br[18] br[17] br[16] br[15] br[14] br[13] br[12] br[11] br[10] br[9] br[8] br[7] br[6] br[5] br[4] br[3] br[2] br[1] br[0] vss 

xmux_0 
+ we[0] wmask[0] data[0] data_b[0] bl[0] br[0] vss 
+ write_mux 
* No parameters

xmux_1 
+ we[1] wmask[0] data[0] data_b[0] bl[1] br[1] vss 
+ write_mux 
* No parameters

xmux_2 
+ we[2] wmask[0] data[0] data_b[0] bl[2] br[2] vss 
+ write_mux 
* No parameters

xmux_3 
+ we[3] wmask[0] data[0] data_b[0] bl[3] br[3] vss 
+ write_mux 
* No parameters

xmux_4 
+ we[4] wmask[0] data[0] data_b[0] bl[4] br[4] vss 
+ write_mux 
* No parameters

xmux_5 
+ we[5] wmask[0] data[0] data_b[0] bl[5] br[5] vss 
+ write_mux 
* No parameters

xmux_6 
+ we[6] wmask[0] data[0] data_b[0] bl[6] br[6] vss 
+ write_mux 
* No parameters

xmux_7 
+ we[7] wmask[0] data[0] data_b[0] bl[7] br[7] vss 
+ write_mux 
* No parameters

xmux_8 
+ we[0] wmask[0] data[1] data_b[1] bl[8] br[8] vss 
+ write_mux 
* No parameters

xmux_9 
+ we[1] wmask[0] data[1] data_b[1] bl[9] br[9] vss 
+ write_mux 
* No parameters

xmux_10 
+ we[2] wmask[0] data[1] data_b[1] bl[10] br[10] vss 
+ write_mux 
* No parameters

xmux_11 
+ we[3] wmask[0] data[1] data_b[1] bl[11] br[11] vss 
+ write_mux 
* No parameters

xmux_12 
+ we[4] wmask[0] data[1] data_b[1] bl[12] br[12] vss 
+ write_mux 
* No parameters

xmux_13 
+ we[5] wmask[0] data[1] data_b[1] bl[13] br[13] vss 
+ write_mux 
* No parameters

xmux_14 
+ we[6] wmask[0] data[1] data_b[1] bl[14] br[14] vss 
+ write_mux 
* No parameters

xmux_15 
+ we[7] wmask[0] data[1] data_b[1] bl[15] br[15] vss 
+ write_mux 
* No parameters

xmux_16 
+ we[0] wmask[0] data[2] data_b[2] bl[16] br[16] vss 
+ write_mux 
* No parameters

xmux_17 
+ we[1] wmask[0] data[2] data_b[2] bl[17] br[17] vss 
+ write_mux 
* No parameters

xmux_18 
+ we[2] wmask[0] data[2] data_b[2] bl[18] br[18] vss 
+ write_mux 
* No parameters

xmux_19 
+ we[3] wmask[0] data[2] data_b[2] bl[19] br[19] vss 
+ write_mux 
* No parameters

xmux_20 
+ we[4] wmask[0] data[2] data_b[2] bl[20] br[20] vss 
+ write_mux 
* No parameters

xmux_21 
+ we[5] wmask[0] data[2] data_b[2] bl[21] br[21] vss 
+ write_mux 
* No parameters

xmux_22 
+ we[6] wmask[0] data[2] data_b[2] bl[22] br[22] vss 
+ write_mux 
* No parameters

xmux_23 
+ we[7] wmask[0] data[2] data_b[2] bl[23] br[23] vss 
+ write_mux 
* No parameters

xmux_24 
+ we[0] wmask[0] data[3] data_b[3] bl[24] br[24] vss 
+ write_mux 
* No parameters

xmux_25 
+ we[1] wmask[0] data[3] data_b[3] bl[25] br[25] vss 
+ write_mux 
* No parameters

xmux_26 
+ we[2] wmask[0] data[3] data_b[3] bl[26] br[26] vss 
+ write_mux 
* No parameters

xmux_27 
+ we[3] wmask[0] data[3] data_b[3] bl[27] br[27] vss 
+ write_mux 
* No parameters

xmux_28 
+ we[4] wmask[0] data[3] data_b[3] bl[28] br[28] vss 
+ write_mux 
* No parameters

xmux_29 
+ we[5] wmask[0] data[3] data_b[3] bl[29] br[29] vss 
+ write_mux 
* No parameters

xmux_30 
+ we[6] wmask[0] data[3] data_b[3] bl[30] br[30] vss 
+ write_mux 
* No parameters

xmux_31 
+ we[7] wmask[0] data[3] data_b[3] bl[31] br[31] vss 
+ write_mux 
* No parameters

xmux_32 
+ we[0] wmask[0] data[4] data_b[4] bl[32] br[32] vss 
+ write_mux 
* No parameters

xmux_33 
+ we[1] wmask[0] data[4] data_b[4] bl[33] br[33] vss 
+ write_mux 
* No parameters

xmux_34 
+ we[2] wmask[0] data[4] data_b[4] bl[34] br[34] vss 
+ write_mux 
* No parameters

xmux_35 
+ we[3] wmask[0] data[4] data_b[4] bl[35] br[35] vss 
+ write_mux 
* No parameters

xmux_36 
+ we[4] wmask[0] data[4] data_b[4] bl[36] br[36] vss 
+ write_mux 
* No parameters

xmux_37 
+ we[5] wmask[0] data[4] data_b[4] bl[37] br[37] vss 
+ write_mux 
* No parameters

xmux_38 
+ we[6] wmask[0] data[4] data_b[4] bl[38] br[38] vss 
+ write_mux 
* No parameters

xmux_39 
+ we[7] wmask[0] data[4] data_b[4] bl[39] br[39] vss 
+ write_mux 
* No parameters

xmux_40 
+ we[0] wmask[0] data[5] data_b[5] bl[40] br[40] vss 
+ write_mux 
* No parameters

xmux_41 
+ we[1] wmask[0] data[5] data_b[5] bl[41] br[41] vss 
+ write_mux 
* No parameters

xmux_42 
+ we[2] wmask[0] data[5] data_b[5] bl[42] br[42] vss 
+ write_mux 
* No parameters

xmux_43 
+ we[3] wmask[0] data[5] data_b[5] bl[43] br[43] vss 
+ write_mux 
* No parameters

xmux_44 
+ we[4] wmask[0] data[5] data_b[5] bl[44] br[44] vss 
+ write_mux 
* No parameters

xmux_45 
+ we[5] wmask[0] data[5] data_b[5] bl[45] br[45] vss 
+ write_mux 
* No parameters

xmux_46 
+ we[6] wmask[0] data[5] data_b[5] bl[46] br[46] vss 
+ write_mux 
* No parameters

xmux_47 
+ we[7] wmask[0] data[5] data_b[5] bl[47] br[47] vss 
+ write_mux 
* No parameters

xmux_48 
+ we[0] wmask[0] data[6] data_b[6] bl[48] br[48] vss 
+ write_mux 
* No parameters

xmux_49 
+ we[1] wmask[0] data[6] data_b[6] bl[49] br[49] vss 
+ write_mux 
* No parameters

xmux_50 
+ we[2] wmask[0] data[6] data_b[6] bl[50] br[50] vss 
+ write_mux 
* No parameters

xmux_51 
+ we[3] wmask[0] data[6] data_b[6] bl[51] br[51] vss 
+ write_mux 
* No parameters

xmux_52 
+ we[4] wmask[0] data[6] data_b[6] bl[52] br[52] vss 
+ write_mux 
* No parameters

xmux_53 
+ we[5] wmask[0] data[6] data_b[6] bl[53] br[53] vss 
+ write_mux 
* No parameters

xmux_54 
+ we[6] wmask[0] data[6] data_b[6] bl[54] br[54] vss 
+ write_mux 
* No parameters

xmux_55 
+ we[7] wmask[0] data[6] data_b[6] bl[55] br[55] vss 
+ write_mux 
* No parameters

xmux_56 
+ we[0] wmask[0] data[7] data_b[7] bl[56] br[56] vss 
+ write_mux 
* No parameters

xmux_57 
+ we[1] wmask[0] data[7] data_b[7] bl[57] br[57] vss 
+ write_mux 
* No parameters

xmux_58 
+ we[2] wmask[0] data[7] data_b[7] bl[58] br[58] vss 
+ write_mux 
* No parameters

xmux_59 
+ we[3] wmask[0] data[7] data_b[7] bl[59] br[59] vss 
+ write_mux 
* No parameters

xmux_60 
+ we[4] wmask[0] data[7] data_b[7] bl[60] br[60] vss 
+ write_mux 
* No parameters

xmux_61 
+ we[5] wmask[0] data[7] data_b[7] bl[61] br[61] vss 
+ write_mux 
* No parameters

xmux_62 
+ we[6] wmask[0] data[7] data_b[7] bl[62] br[62] vss 
+ write_mux 
* No parameters

xmux_63 
+ we[7] wmask[0] data[7] data_b[7] bl[63] br[63] vss 
+ write_mux 
* No parameters

xmux_64 
+ we[0] wmask[1] data[8] data_b[8] bl[64] br[64] vss 
+ write_mux 
* No parameters

xmux_65 
+ we[1] wmask[1] data[8] data_b[8] bl[65] br[65] vss 
+ write_mux 
* No parameters

xmux_66 
+ we[2] wmask[1] data[8] data_b[8] bl[66] br[66] vss 
+ write_mux 
* No parameters

xmux_67 
+ we[3] wmask[1] data[8] data_b[8] bl[67] br[67] vss 
+ write_mux 
* No parameters

xmux_68 
+ we[4] wmask[1] data[8] data_b[8] bl[68] br[68] vss 
+ write_mux 
* No parameters

xmux_69 
+ we[5] wmask[1] data[8] data_b[8] bl[69] br[69] vss 
+ write_mux 
* No parameters

xmux_70 
+ we[6] wmask[1] data[8] data_b[8] bl[70] br[70] vss 
+ write_mux 
* No parameters

xmux_71 
+ we[7] wmask[1] data[8] data_b[8] bl[71] br[71] vss 
+ write_mux 
* No parameters

xmux_72 
+ we[0] wmask[1] data[9] data_b[9] bl[72] br[72] vss 
+ write_mux 
* No parameters

xmux_73 
+ we[1] wmask[1] data[9] data_b[9] bl[73] br[73] vss 
+ write_mux 
* No parameters

xmux_74 
+ we[2] wmask[1] data[9] data_b[9] bl[74] br[74] vss 
+ write_mux 
* No parameters

xmux_75 
+ we[3] wmask[1] data[9] data_b[9] bl[75] br[75] vss 
+ write_mux 
* No parameters

xmux_76 
+ we[4] wmask[1] data[9] data_b[9] bl[76] br[76] vss 
+ write_mux 
* No parameters

xmux_77 
+ we[5] wmask[1] data[9] data_b[9] bl[77] br[77] vss 
+ write_mux 
* No parameters

xmux_78 
+ we[6] wmask[1] data[9] data_b[9] bl[78] br[78] vss 
+ write_mux 
* No parameters

xmux_79 
+ we[7] wmask[1] data[9] data_b[9] bl[79] br[79] vss 
+ write_mux 
* No parameters

xmux_80 
+ we[0] wmask[1] data[10] data_b[10] bl[80] br[80] vss 
+ write_mux 
* No parameters

xmux_81 
+ we[1] wmask[1] data[10] data_b[10] bl[81] br[81] vss 
+ write_mux 
* No parameters

xmux_82 
+ we[2] wmask[1] data[10] data_b[10] bl[82] br[82] vss 
+ write_mux 
* No parameters

xmux_83 
+ we[3] wmask[1] data[10] data_b[10] bl[83] br[83] vss 
+ write_mux 
* No parameters

xmux_84 
+ we[4] wmask[1] data[10] data_b[10] bl[84] br[84] vss 
+ write_mux 
* No parameters

xmux_85 
+ we[5] wmask[1] data[10] data_b[10] bl[85] br[85] vss 
+ write_mux 
* No parameters

xmux_86 
+ we[6] wmask[1] data[10] data_b[10] bl[86] br[86] vss 
+ write_mux 
* No parameters

xmux_87 
+ we[7] wmask[1] data[10] data_b[10] bl[87] br[87] vss 
+ write_mux 
* No parameters

xmux_88 
+ we[0] wmask[1] data[11] data_b[11] bl[88] br[88] vss 
+ write_mux 
* No parameters

xmux_89 
+ we[1] wmask[1] data[11] data_b[11] bl[89] br[89] vss 
+ write_mux 
* No parameters

xmux_90 
+ we[2] wmask[1] data[11] data_b[11] bl[90] br[90] vss 
+ write_mux 
* No parameters

xmux_91 
+ we[3] wmask[1] data[11] data_b[11] bl[91] br[91] vss 
+ write_mux 
* No parameters

xmux_92 
+ we[4] wmask[1] data[11] data_b[11] bl[92] br[92] vss 
+ write_mux 
* No parameters

xmux_93 
+ we[5] wmask[1] data[11] data_b[11] bl[93] br[93] vss 
+ write_mux 
* No parameters

xmux_94 
+ we[6] wmask[1] data[11] data_b[11] bl[94] br[94] vss 
+ write_mux 
* No parameters

xmux_95 
+ we[7] wmask[1] data[11] data_b[11] bl[95] br[95] vss 
+ write_mux 
* No parameters

xmux_96 
+ we[0] wmask[1] data[12] data_b[12] bl[96] br[96] vss 
+ write_mux 
* No parameters

xmux_97 
+ we[1] wmask[1] data[12] data_b[12] bl[97] br[97] vss 
+ write_mux 
* No parameters

xmux_98 
+ we[2] wmask[1] data[12] data_b[12] bl[98] br[98] vss 
+ write_mux 
* No parameters

xmux_99 
+ we[3] wmask[1] data[12] data_b[12] bl[99] br[99] vss 
+ write_mux 
* No parameters

xmux_100 
+ we[4] wmask[1] data[12] data_b[12] bl[100] br[100] vss 
+ write_mux 
* No parameters

xmux_101 
+ we[5] wmask[1] data[12] data_b[12] bl[101] br[101] vss 
+ write_mux 
* No parameters

xmux_102 
+ we[6] wmask[1] data[12] data_b[12] bl[102] br[102] vss 
+ write_mux 
* No parameters

xmux_103 
+ we[7] wmask[1] data[12] data_b[12] bl[103] br[103] vss 
+ write_mux 
* No parameters

xmux_104 
+ we[0] wmask[1] data[13] data_b[13] bl[104] br[104] vss 
+ write_mux 
* No parameters

xmux_105 
+ we[1] wmask[1] data[13] data_b[13] bl[105] br[105] vss 
+ write_mux 
* No parameters

xmux_106 
+ we[2] wmask[1] data[13] data_b[13] bl[106] br[106] vss 
+ write_mux 
* No parameters

xmux_107 
+ we[3] wmask[1] data[13] data_b[13] bl[107] br[107] vss 
+ write_mux 
* No parameters

xmux_108 
+ we[4] wmask[1] data[13] data_b[13] bl[108] br[108] vss 
+ write_mux 
* No parameters

xmux_109 
+ we[5] wmask[1] data[13] data_b[13] bl[109] br[109] vss 
+ write_mux 
* No parameters

xmux_110 
+ we[6] wmask[1] data[13] data_b[13] bl[110] br[110] vss 
+ write_mux 
* No parameters

xmux_111 
+ we[7] wmask[1] data[13] data_b[13] bl[111] br[111] vss 
+ write_mux 
* No parameters

xmux_112 
+ we[0] wmask[1] data[14] data_b[14] bl[112] br[112] vss 
+ write_mux 
* No parameters

xmux_113 
+ we[1] wmask[1] data[14] data_b[14] bl[113] br[113] vss 
+ write_mux 
* No parameters

xmux_114 
+ we[2] wmask[1] data[14] data_b[14] bl[114] br[114] vss 
+ write_mux 
* No parameters

xmux_115 
+ we[3] wmask[1] data[14] data_b[14] bl[115] br[115] vss 
+ write_mux 
* No parameters

xmux_116 
+ we[4] wmask[1] data[14] data_b[14] bl[116] br[116] vss 
+ write_mux 
* No parameters

xmux_117 
+ we[5] wmask[1] data[14] data_b[14] bl[117] br[117] vss 
+ write_mux 
* No parameters

xmux_118 
+ we[6] wmask[1] data[14] data_b[14] bl[118] br[118] vss 
+ write_mux 
* No parameters

xmux_119 
+ we[7] wmask[1] data[14] data_b[14] bl[119] br[119] vss 
+ write_mux 
* No parameters

xmux_120 
+ we[0] wmask[1] data[15] data_b[15] bl[120] br[120] vss 
+ write_mux 
* No parameters

xmux_121 
+ we[1] wmask[1] data[15] data_b[15] bl[121] br[121] vss 
+ write_mux 
* No parameters

xmux_122 
+ we[2] wmask[1] data[15] data_b[15] bl[122] br[122] vss 
+ write_mux 
* No parameters

xmux_123 
+ we[3] wmask[1] data[15] data_b[15] bl[123] br[123] vss 
+ write_mux 
* No parameters

xmux_124 
+ we[4] wmask[1] data[15] data_b[15] bl[124] br[124] vss 
+ write_mux 
* No parameters

xmux_125 
+ we[5] wmask[1] data[15] data_b[15] bl[125] br[125] vss 
+ write_mux 
* No parameters

xmux_126 
+ we[6] wmask[1] data[15] data_b[15] bl[126] br[126] vss 
+ write_mux 
* No parameters

xmux_127 
+ we[7] wmask[1] data[15] data_b[15] bl[127] br[127] vss 
+ write_mux 
* No parameters

xmux_128 
+ we[0] wmask[2] data[16] data_b[16] bl[128] br[128] vss 
+ write_mux 
* No parameters

xmux_129 
+ we[1] wmask[2] data[16] data_b[16] bl[129] br[129] vss 
+ write_mux 
* No parameters

xmux_130 
+ we[2] wmask[2] data[16] data_b[16] bl[130] br[130] vss 
+ write_mux 
* No parameters

xmux_131 
+ we[3] wmask[2] data[16] data_b[16] bl[131] br[131] vss 
+ write_mux 
* No parameters

xmux_132 
+ we[4] wmask[2] data[16] data_b[16] bl[132] br[132] vss 
+ write_mux 
* No parameters

xmux_133 
+ we[5] wmask[2] data[16] data_b[16] bl[133] br[133] vss 
+ write_mux 
* No parameters

xmux_134 
+ we[6] wmask[2] data[16] data_b[16] bl[134] br[134] vss 
+ write_mux 
* No parameters

xmux_135 
+ we[7] wmask[2] data[16] data_b[16] bl[135] br[135] vss 
+ write_mux 
* No parameters

xmux_136 
+ we[0] wmask[2] data[17] data_b[17] bl[136] br[136] vss 
+ write_mux 
* No parameters

xmux_137 
+ we[1] wmask[2] data[17] data_b[17] bl[137] br[137] vss 
+ write_mux 
* No parameters

xmux_138 
+ we[2] wmask[2] data[17] data_b[17] bl[138] br[138] vss 
+ write_mux 
* No parameters

xmux_139 
+ we[3] wmask[2] data[17] data_b[17] bl[139] br[139] vss 
+ write_mux 
* No parameters

xmux_140 
+ we[4] wmask[2] data[17] data_b[17] bl[140] br[140] vss 
+ write_mux 
* No parameters

xmux_141 
+ we[5] wmask[2] data[17] data_b[17] bl[141] br[141] vss 
+ write_mux 
* No parameters

xmux_142 
+ we[6] wmask[2] data[17] data_b[17] bl[142] br[142] vss 
+ write_mux 
* No parameters

xmux_143 
+ we[7] wmask[2] data[17] data_b[17] bl[143] br[143] vss 
+ write_mux 
* No parameters

xmux_144 
+ we[0] wmask[2] data[18] data_b[18] bl[144] br[144] vss 
+ write_mux 
* No parameters

xmux_145 
+ we[1] wmask[2] data[18] data_b[18] bl[145] br[145] vss 
+ write_mux 
* No parameters

xmux_146 
+ we[2] wmask[2] data[18] data_b[18] bl[146] br[146] vss 
+ write_mux 
* No parameters

xmux_147 
+ we[3] wmask[2] data[18] data_b[18] bl[147] br[147] vss 
+ write_mux 
* No parameters

xmux_148 
+ we[4] wmask[2] data[18] data_b[18] bl[148] br[148] vss 
+ write_mux 
* No parameters

xmux_149 
+ we[5] wmask[2] data[18] data_b[18] bl[149] br[149] vss 
+ write_mux 
* No parameters

xmux_150 
+ we[6] wmask[2] data[18] data_b[18] bl[150] br[150] vss 
+ write_mux 
* No parameters

xmux_151 
+ we[7] wmask[2] data[18] data_b[18] bl[151] br[151] vss 
+ write_mux 
* No parameters

xmux_152 
+ we[0] wmask[2] data[19] data_b[19] bl[152] br[152] vss 
+ write_mux 
* No parameters

xmux_153 
+ we[1] wmask[2] data[19] data_b[19] bl[153] br[153] vss 
+ write_mux 
* No parameters

xmux_154 
+ we[2] wmask[2] data[19] data_b[19] bl[154] br[154] vss 
+ write_mux 
* No parameters

xmux_155 
+ we[3] wmask[2] data[19] data_b[19] bl[155] br[155] vss 
+ write_mux 
* No parameters

xmux_156 
+ we[4] wmask[2] data[19] data_b[19] bl[156] br[156] vss 
+ write_mux 
* No parameters

xmux_157 
+ we[5] wmask[2] data[19] data_b[19] bl[157] br[157] vss 
+ write_mux 
* No parameters

xmux_158 
+ we[6] wmask[2] data[19] data_b[19] bl[158] br[158] vss 
+ write_mux 
* No parameters

xmux_159 
+ we[7] wmask[2] data[19] data_b[19] bl[159] br[159] vss 
+ write_mux 
* No parameters

xmux_160 
+ we[0] wmask[2] data[20] data_b[20] bl[160] br[160] vss 
+ write_mux 
* No parameters

xmux_161 
+ we[1] wmask[2] data[20] data_b[20] bl[161] br[161] vss 
+ write_mux 
* No parameters

xmux_162 
+ we[2] wmask[2] data[20] data_b[20] bl[162] br[162] vss 
+ write_mux 
* No parameters

xmux_163 
+ we[3] wmask[2] data[20] data_b[20] bl[163] br[163] vss 
+ write_mux 
* No parameters

xmux_164 
+ we[4] wmask[2] data[20] data_b[20] bl[164] br[164] vss 
+ write_mux 
* No parameters

xmux_165 
+ we[5] wmask[2] data[20] data_b[20] bl[165] br[165] vss 
+ write_mux 
* No parameters

xmux_166 
+ we[6] wmask[2] data[20] data_b[20] bl[166] br[166] vss 
+ write_mux 
* No parameters

xmux_167 
+ we[7] wmask[2] data[20] data_b[20] bl[167] br[167] vss 
+ write_mux 
* No parameters

xmux_168 
+ we[0] wmask[2] data[21] data_b[21] bl[168] br[168] vss 
+ write_mux 
* No parameters

xmux_169 
+ we[1] wmask[2] data[21] data_b[21] bl[169] br[169] vss 
+ write_mux 
* No parameters

xmux_170 
+ we[2] wmask[2] data[21] data_b[21] bl[170] br[170] vss 
+ write_mux 
* No parameters

xmux_171 
+ we[3] wmask[2] data[21] data_b[21] bl[171] br[171] vss 
+ write_mux 
* No parameters

xmux_172 
+ we[4] wmask[2] data[21] data_b[21] bl[172] br[172] vss 
+ write_mux 
* No parameters

xmux_173 
+ we[5] wmask[2] data[21] data_b[21] bl[173] br[173] vss 
+ write_mux 
* No parameters

xmux_174 
+ we[6] wmask[2] data[21] data_b[21] bl[174] br[174] vss 
+ write_mux 
* No parameters

xmux_175 
+ we[7] wmask[2] data[21] data_b[21] bl[175] br[175] vss 
+ write_mux 
* No parameters

xmux_176 
+ we[0] wmask[2] data[22] data_b[22] bl[176] br[176] vss 
+ write_mux 
* No parameters

xmux_177 
+ we[1] wmask[2] data[22] data_b[22] bl[177] br[177] vss 
+ write_mux 
* No parameters

xmux_178 
+ we[2] wmask[2] data[22] data_b[22] bl[178] br[178] vss 
+ write_mux 
* No parameters

xmux_179 
+ we[3] wmask[2] data[22] data_b[22] bl[179] br[179] vss 
+ write_mux 
* No parameters

xmux_180 
+ we[4] wmask[2] data[22] data_b[22] bl[180] br[180] vss 
+ write_mux 
* No parameters

xmux_181 
+ we[5] wmask[2] data[22] data_b[22] bl[181] br[181] vss 
+ write_mux 
* No parameters

xmux_182 
+ we[6] wmask[2] data[22] data_b[22] bl[182] br[182] vss 
+ write_mux 
* No parameters

xmux_183 
+ we[7] wmask[2] data[22] data_b[22] bl[183] br[183] vss 
+ write_mux 
* No parameters

xmux_184 
+ we[0] wmask[2] data[23] data_b[23] bl[184] br[184] vss 
+ write_mux 
* No parameters

xmux_185 
+ we[1] wmask[2] data[23] data_b[23] bl[185] br[185] vss 
+ write_mux 
* No parameters

xmux_186 
+ we[2] wmask[2] data[23] data_b[23] bl[186] br[186] vss 
+ write_mux 
* No parameters

xmux_187 
+ we[3] wmask[2] data[23] data_b[23] bl[187] br[187] vss 
+ write_mux 
* No parameters

xmux_188 
+ we[4] wmask[2] data[23] data_b[23] bl[188] br[188] vss 
+ write_mux 
* No parameters

xmux_189 
+ we[5] wmask[2] data[23] data_b[23] bl[189] br[189] vss 
+ write_mux 
* No parameters

xmux_190 
+ we[6] wmask[2] data[23] data_b[23] bl[190] br[190] vss 
+ write_mux 
* No parameters

xmux_191 
+ we[7] wmask[2] data[23] data_b[23] bl[191] br[191] vss 
+ write_mux 
* No parameters

xmux_192 
+ we[0] wmask[3] data[24] data_b[24] bl[192] br[192] vss 
+ write_mux 
* No parameters

xmux_193 
+ we[1] wmask[3] data[24] data_b[24] bl[193] br[193] vss 
+ write_mux 
* No parameters

xmux_194 
+ we[2] wmask[3] data[24] data_b[24] bl[194] br[194] vss 
+ write_mux 
* No parameters

xmux_195 
+ we[3] wmask[3] data[24] data_b[24] bl[195] br[195] vss 
+ write_mux 
* No parameters

xmux_196 
+ we[4] wmask[3] data[24] data_b[24] bl[196] br[196] vss 
+ write_mux 
* No parameters

xmux_197 
+ we[5] wmask[3] data[24] data_b[24] bl[197] br[197] vss 
+ write_mux 
* No parameters

xmux_198 
+ we[6] wmask[3] data[24] data_b[24] bl[198] br[198] vss 
+ write_mux 
* No parameters

xmux_199 
+ we[7] wmask[3] data[24] data_b[24] bl[199] br[199] vss 
+ write_mux 
* No parameters

xmux_200 
+ we[0] wmask[3] data[25] data_b[25] bl[200] br[200] vss 
+ write_mux 
* No parameters

xmux_201 
+ we[1] wmask[3] data[25] data_b[25] bl[201] br[201] vss 
+ write_mux 
* No parameters

xmux_202 
+ we[2] wmask[3] data[25] data_b[25] bl[202] br[202] vss 
+ write_mux 
* No parameters

xmux_203 
+ we[3] wmask[3] data[25] data_b[25] bl[203] br[203] vss 
+ write_mux 
* No parameters

xmux_204 
+ we[4] wmask[3] data[25] data_b[25] bl[204] br[204] vss 
+ write_mux 
* No parameters

xmux_205 
+ we[5] wmask[3] data[25] data_b[25] bl[205] br[205] vss 
+ write_mux 
* No parameters

xmux_206 
+ we[6] wmask[3] data[25] data_b[25] bl[206] br[206] vss 
+ write_mux 
* No parameters

xmux_207 
+ we[7] wmask[3] data[25] data_b[25] bl[207] br[207] vss 
+ write_mux 
* No parameters

xmux_208 
+ we[0] wmask[3] data[26] data_b[26] bl[208] br[208] vss 
+ write_mux 
* No parameters

xmux_209 
+ we[1] wmask[3] data[26] data_b[26] bl[209] br[209] vss 
+ write_mux 
* No parameters

xmux_210 
+ we[2] wmask[3] data[26] data_b[26] bl[210] br[210] vss 
+ write_mux 
* No parameters

xmux_211 
+ we[3] wmask[3] data[26] data_b[26] bl[211] br[211] vss 
+ write_mux 
* No parameters

xmux_212 
+ we[4] wmask[3] data[26] data_b[26] bl[212] br[212] vss 
+ write_mux 
* No parameters

xmux_213 
+ we[5] wmask[3] data[26] data_b[26] bl[213] br[213] vss 
+ write_mux 
* No parameters

xmux_214 
+ we[6] wmask[3] data[26] data_b[26] bl[214] br[214] vss 
+ write_mux 
* No parameters

xmux_215 
+ we[7] wmask[3] data[26] data_b[26] bl[215] br[215] vss 
+ write_mux 
* No parameters

xmux_216 
+ we[0] wmask[3] data[27] data_b[27] bl[216] br[216] vss 
+ write_mux 
* No parameters

xmux_217 
+ we[1] wmask[3] data[27] data_b[27] bl[217] br[217] vss 
+ write_mux 
* No parameters

xmux_218 
+ we[2] wmask[3] data[27] data_b[27] bl[218] br[218] vss 
+ write_mux 
* No parameters

xmux_219 
+ we[3] wmask[3] data[27] data_b[27] bl[219] br[219] vss 
+ write_mux 
* No parameters

xmux_220 
+ we[4] wmask[3] data[27] data_b[27] bl[220] br[220] vss 
+ write_mux 
* No parameters

xmux_221 
+ we[5] wmask[3] data[27] data_b[27] bl[221] br[221] vss 
+ write_mux 
* No parameters

xmux_222 
+ we[6] wmask[3] data[27] data_b[27] bl[222] br[222] vss 
+ write_mux 
* No parameters

xmux_223 
+ we[7] wmask[3] data[27] data_b[27] bl[223] br[223] vss 
+ write_mux 
* No parameters

xmux_224 
+ we[0] wmask[3] data[28] data_b[28] bl[224] br[224] vss 
+ write_mux 
* No parameters

xmux_225 
+ we[1] wmask[3] data[28] data_b[28] bl[225] br[225] vss 
+ write_mux 
* No parameters

xmux_226 
+ we[2] wmask[3] data[28] data_b[28] bl[226] br[226] vss 
+ write_mux 
* No parameters

xmux_227 
+ we[3] wmask[3] data[28] data_b[28] bl[227] br[227] vss 
+ write_mux 
* No parameters

xmux_228 
+ we[4] wmask[3] data[28] data_b[28] bl[228] br[228] vss 
+ write_mux 
* No parameters

xmux_229 
+ we[5] wmask[3] data[28] data_b[28] bl[229] br[229] vss 
+ write_mux 
* No parameters

xmux_230 
+ we[6] wmask[3] data[28] data_b[28] bl[230] br[230] vss 
+ write_mux 
* No parameters

xmux_231 
+ we[7] wmask[3] data[28] data_b[28] bl[231] br[231] vss 
+ write_mux 
* No parameters

xmux_232 
+ we[0] wmask[3] data[29] data_b[29] bl[232] br[232] vss 
+ write_mux 
* No parameters

xmux_233 
+ we[1] wmask[3] data[29] data_b[29] bl[233] br[233] vss 
+ write_mux 
* No parameters

xmux_234 
+ we[2] wmask[3] data[29] data_b[29] bl[234] br[234] vss 
+ write_mux 
* No parameters

xmux_235 
+ we[3] wmask[3] data[29] data_b[29] bl[235] br[235] vss 
+ write_mux 
* No parameters

xmux_236 
+ we[4] wmask[3] data[29] data_b[29] bl[236] br[236] vss 
+ write_mux 
* No parameters

xmux_237 
+ we[5] wmask[3] data[29] data_b[29] bl[237] br[237] vss 
+ write_mux 
* No parameters

xmux_238 
+ we[6] wmask[3] data[29] data_b[29] bl[238] br[238] vss 
+ write_mux 
* No parameters

xmux_239 
+ we[7] wmask[3] data[29] data_b[29] bl[239] br[239] vss 
+ write_mux 
* No parameters

xmux_240 
+ we[0] wmask[3] data[30] data_b[30] bl[240] br[240] vss 
+ write_mux 
* No parameters

xmux_241 
+ we[1] wmask[3] data[30] data_b[30] bl[241] br[241] vss 
+ write_mux 
* No parameters

xmux_242 
+ we[2] wmask[3] data[30] data_b[30] bl[242] br[242] vss 
+ write_mux 
* No parameters

xmux_243 
+ we[3] wmask[3] data[30] data_b[30] bl[243] br[243] vss 
+ write_mux 
* No parameters

xmux_244 
+ we[4] wmask[3] data[30] data_b[30] bl[244] br[244] vss 
+ write_mux 
* No parameters

xmux_245 
+ we[5] wmask[3] data[30] data_b[30] bl[245] br[245] vss 
+ write_mux 
* No parameters

xmux_246 
+ we[6] wmask[3] data[30] data_b[30] bl[246] br[246] vss 
+ write_mux 
* No parameters

xmux_247 
+ we[7] wmask[3] data[30] data_b[30] bl[247] br[247] vss 
+ write_mux 
* No parameters

xmux_248 
+ we[0] wmask[3] data[31] data_b[31] bl[248] br[248] vss 
+ write_mux 
* No parameters

xmux_249 
+ we[1] wmask[3] data[31] data_b[31] bl[249] br[249] vss 
+ write_mux 
* No parameters

xmux_250 
+ we[2] wmask[3] data[31] data_b[31] bl[250] br[250] vss 
+ write_mux 
* No parameters

xmux_251 
+ we[3] wmask[3] data[31] data_b[31] bl[251] br[251] vss 
+ write_mux 
* No parameters

xmux_252 
+ we[4] wmask[3] data[31] data_b[31] bl[252] br[252] vss 
+ write_mux 
* No parameters

xmux_253 
+ we[5] wmask[3] data[31] data_b[31] bl[253] br[253] vss 
+ write_mux 
* No parameters

xmux_254 
+ we[6] wmask[3] data[31] data_b[31] bl[254] br[254] vss 
+ write_mux 
* No parameters

xmux_255 
+ we[7] wmask[3] data[31] data_b[31] bl[255] br[255] vss 
+ write_mux 
* No parameters

.ENDS

.SUBCKT data_dff_array 
+ vdd vss clk d[31] d[30] d[29] d[28] d[27] d[26] d[25] d[24] d[23] d[22] d[21] d[20] d[19] d[18] d[17] d[16] d[15] d[14] d[13] d[12] d[11] d[10] d[9] d[8] d[7] d[6] d[5] d[4] d[3] d[2] d[1] d[0] q[31] q[30] q[29] q[28] q[27] q[26] q[25] q[24] q[23] q[22] q[21] q[20] q[19] q[18] q[17] q[16] q[15] q[14] q[13] q[12] q[11] q[10] q[9] q[8] q[7] q[6] q[5] q[4] q[3] q[2] q[1] q[0] q_b[31] q_b[30] q_b[29] q_b[28] q_b[27] q_b[26] q_b[25] q_b[24] q_b[23] q_b[22] q_b[21] q_b[20] q_b[19] q_b[18] q_b[17] q_b[16] q_b[15] q_b[14] q_b[13] q_b[12] q_b[11] q_b[10] q_b[9] q_b[8] q_b[7] q_b[6] q_b[5] q_b[4] q_b[3] q_b[2] q_b[1] q_b[0] 

xdff_0 
+ vdd vss clk d[0] q[0] q_b[0] 
+ openram_dff 
* No parameters

xdff_1 
+ vdd vss clk d[1] q[1] q_b[1] 
+ openram_dff 
* No parameters

xdff_2 
+ vdd vss clk d[2] q[2] q_b[2] 
+ openram_dff 
* No parameters

xdff_3 
+ vdd vss clk d[3] q[3] q_b[3] 
+ openram_dff 
* No parameters

xdff_4 
+ vdd vss clk d[4] q[4] q_b[4] 
+ openram_dff 
* No parameters

xdff_5 
+ vdd vss clk d[5] q[5] q_b[5] 
+ openram_dff 
* No parameters

xdff_6 
+ vdd vss clk d[6] q[6] q_b[6] 
+ openram_dff 
* No parameters

xdff_7 
+ vdd vss clk d[7] q[7] q_b[7] 
+ openram_dff 
* No parameters

xdff_8 
+ vdd vss clk d[8] q[8] q_b[8] 
+ openram_dff 
* No parameters

xdff_9 
+ vdd vss clk d[9] q[9] q_b[9] 
+ openram_dff 
* No parameters

xdff_10 
+ vdd vss clk d[10] q[10] q_b[10] 
+ openram_dff 
* No parameters

xdff_11 
+ vdd vss clk d[11] q[11] q_b[11] 
+ openram_dff 
* No parameters

xdff_12 
+ vdd vss clk d[12] q[12] q_b[12] 
+ openram_dff 
* No parameters

xdff_13 
+ vdd vss clk d[13] q[13] q_b[13] 
+ openram_dff 
* No parameters

xdff_14 
+ vdd vss clk d[14] q[14] q_b[14] 
+ openram_dff 
* No parameters

xdff_15 
+ vdd vss clk d[15] q[15] q_b[15] 
+ openram_dff 
* No parameters

xdff_16 
+ vdd vss clk d[16] q[16] q_b[16] 
+ openram_dff 
* No parameters

xdff_17 
+ vdd vss clk d[17] q[17] q_b[17] 
+ openram_dff 
* No parameters

xdff_18 
+ vdd vss clk d[18] q[18] q_b[18] 
+ openram_dff 
* No parameters

xdff_19 
+ vdd vss clk d[19] q[19] q_b[19] 
+ openram_dff 
* No parameters

xdff_20 
+ vdd vss clk d[20] q[20] q_b[20] 
+ openram_dff 
* No parameters

xdff_21 
+ vdd vss clk d[21] q[21] q_b[21] 
+ openram_dff 
* No parameters

xdff_22 
+ vdd vss clk d[22] q[22] q_b[22] 
+ openram_dff 
* No parameters

xdff_23 
+ vdd vss clk d[23] q[23] q_b[23] 
+ openram_dff 
* No parameters

xdff_24 
+ vdd vss clk d[24] q[24] q_b[24] 
+ openram_dff 
* No parameters

xdff_25 
+ vdd vss clk d[25] q[25] q_b[25] 
+ openram_dff 
* No parameters

xdff_26 
+ vdd vss clk d[26] q[26] q_b[26] 
+ openram_dff 
* No parameters

xdff_27 
+ vdd vss clk d[27] q[27] q_b[27] 
+ openram_dff 
* No parameters

xdff_28 
+ vdd vss clk d[28] q[28] q_b[28] 
+ openram_dff 
* No parameters

xdff_29 
+ vdd vss clk d[29] q[29] q_b[29] 
+ openram_dff 
* No parameters

xdff_30 
+ vdd vss clk d[30] q[30] q_b[30] 
+ openram_dff 
* No parameters

xdff_31 
+ vdd vss clk d[31] q[31] q_b[31] 
+ openram_dff 
* No parameters

.ENDS

.SUBCKT addr_dff_array 
+ vdd vss clk d[9] d[8] d[7] d[6] d[5] d[4] d[3] d[2] d[1] d[0] q[9] q[8] q[7] q[6] q[5] q[4] q[3] q[2] q[1] q[0] q_b[9] q_b[8] q_b[7] q_b[6] q_b[5] q_b[4] q_b[3] q_b[2] q_b[1] q_b[0] 

xdff_0 
+ vdd vss clk d[0] q[0] q_b[0] 
+ openram_dff 
* No parameters

xdff_1 
+ vdd vss clk d[1] q[1] q_b[1] 
+ openram_dff 
* No parameters

xdff_2 
+ vdd vss clk d[2] q[2] q_b[2] 
+ openram_dff 
* No parameters

xdff_3 
+ vdd vss clk d[3] q[3] q_b[3] 
+ openram_dff 
* No parameters

xdff_4 
+ vdd vss clk d[4] q[4] q_b[4] 
+ openram_dff 
* No parameters

xdff_5 
+ vdd vss clk d[5] q[5] q_b[5] 
+ openram_dff 
* No parameters

xdff_6 
+ vdd vss clk d[6] q[6] q_b[6] 
+ openram_dff 
* No parameters

xdff_7 
+ vdd vss clk d[7] q[7] q_b[7] 
+ openram_dff 
* No parameters

xdff_8 
+ vdd vss clk d[8] q[8] q_b[8] 
+ openram_dff 
* No parameters

xdff_9 
+ vdd vss clk d[9] q[9] q_b[9] 
+ openram_dff 
* No parameters

.ENDS

.SUBCKT wmask_dff_array 
+ vdd vss clk d[3] d[2] d[1] d[0] q[3] q[2] q[1] q[0] q_b[3] q_b[2] q_b[1] q_b[0] 

xdff_0 
+ vdd vss clk d[0] q[0] q_b[0] 
+ openram_dff 
* No parameters

xdff_1 
+ vdd vss clk d[1] q[1] q_b[1] 
+ openram_dff 
* No parameters

xdff_2 
+ vdd vss clk d[2] q[2] q_b[2] 
+ openram_dff 
* No parameters

xdff_3 
+ vdd vss clk d[3] q[3] q_b[3] 
+ openram_dff 
* No parameters

.ENDS

.SUBCKT col_data_inv 
+ din din_b vdd vss 

xMP0 
+ din_b din vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.6' l='0.15' 

xMN0 
+ din_b din vss vss 
+ sky130_fd_pr__nfet_01v8 
+ w='1.4' l='0.15' 

.ENDS

.SUBCKT col_inv_array 
+ din[31] din[30] din[29] din[28] din[27] din[26] din[25] din[24] din[23] din[22] din[21] din[20] din[19] din[18] din[17] din[16] din[15] din[14] din[13] din[12] din[11] din[10] din[9] din[8] din[7] din[6] din[5] din[4] din[3] din[2] din[1] din[0] din_b[31] din_b[30] din_b[29] din_b[28] din_b[27] din_b[26] din_b[25] din_b[24] din_b[23] din_b[22] din_b[21] din_b[20] din_b[19] din_b[18] din_b[17] din_b[16] din_b[15] din_b[14] din_b[13] din_b[12] din_b[11] din_b[10] din_b[9] din_b[8] din_b[7] din_b[6] din_b[5] din_b[4] din_b[3] din_b[2] din_b[1] din_b[0] vdd vss 

xinv_0 
+ din[0] din_b[0] vdd vss 
+ col_data_inv 
* No parameters

xinv_1 
+ din[1] din_b[1] vdd vss 
+ col_data_inv 
* No parameters

xinv_2 
+ din[2] din_b[2] vdd vss 
+ col_data_inv 
* No parameters

xinv_3 
+ din[3] din_b[3] vdd vss 
+ col_data_inv 
* No parameters

xinv_4 
+ din[4] din_b[4] vdd vss 
+ col_data_inv 
* No parameters

xinv_5 
+ din[5] din_b[5] vdd vss 
+ col_data_inv 
* No parameters

xinv_6 
+ din[6] din_b[6] vdd vss 
+ col_data_inv 
* No parameters

xinv_7 
+ din[7] din_b[7] vdd vss 
+ col_data_inv 
* No parameters

xinv_8 
+ din[8] din_b[8] vdd vss 
+ col_data_inv 
* No parameters

xinv_9 
+ din[9] din_b[9] vdd vss 
+ col_data_inv 
* No parameters

xinv_10 
+ din[10] din_b[10] vdd vss 
+ col_data_inv 
* No parameters

xinv_11 
+ din[11] din_b[11] vdd vss 
+ col_data_inv 
* No parameters

xinv_12 
+ din[12] din_b[12] vdd vss 
+ col_data_inv 
* No parameters

xinv_13 
+ din[13] din_b[13] vdd vss 
+ col_data_inv 
* No parameters

xinv_14 
+ din[14] din_b[14] vdd vss 
+ col_data_inv 
* No parameters

xinv_15 
+ din[15] din_b[15] vdd vss 
+ col_data_inv 
* No parameters

xinv_16 
+ din[16] din_b[16] vdd vss 
+ col_data_inv 
* No parameters

xinv_17 
+ din[17] din_b[17] vdd vss 
+ col_data_inv 
* No parameters

xinv_18 
+ din[18] din_b[18] vdd vss 
+ col_data_inv 
* No parameters

xinv_19 
+ din[19] din_b[19] vdd vss 
+ col_data_inv 
* No parameters

xinv_20 
+ din[20] din_b[20] vdd vss 
+ col_data_inv 
* No parameters

xinv_21 
+ din[21] din_b[21] vdd vss 
+ col_data_inv 
* No parameters

xinv_22 
+ din[22] din_b[22] vdd vss 
+ col_data_inv 
* No parameters

xinv_23 
+ din[23] din_b[23] vdd vss 
+ col_data_inv 
* No parameters

xinv_24 
+ din[24] din_b[24] vdd vss 
+ col_data_inv 
* No parameters

xinv_25 
+ din[25] din_b[25] vdd vss 
+ col_data_inv 
* No parameters

xinv_26 
+ din[26] din_b[26] vdd vss 
+ col_data_inv 
* No parameters

xinv_27 
+ din[27] din_b[27] vdd vss 
+ col_data_inv 
* No parameters

xinv_28 
+ din[28] din_b[28] vdd vss 
+ col_data_inv 
* No parameters

xinv_29 
+ din[29] din_b[29] vdd vss 
+ col_data_inv 
* No parameters

xinv_30 
+ din[30] din_b[30] vdd vss 
+ col_data_inv 
* No parameters

xinv_31 
+ din[31] din_b[31] vdd vss 
+ col_data_inv 
* No parameters

.ENDS

.SUBCKT sense_amp_array 
+ vdd vss clk bl[31] bl[30] bl[29] bl[28] bl[27] bl[26] bl[25] bl[24] bl[23] bl[22] bl[21] bl[20] bl[19] bl[18] bl[17] bl[16] bl[15] bl[14] bl[13] bl[12] bl[11] bl[10] bl[9] bl[8] bl[7] bl[6] bl[5] bl[4] bl[3] bl[2] bl[1] bl[0] br[31] br[30] br[29] br[28] br[27] br[26] br[25] br[24] br[23] br[22] br[21] br[20] br[19] br[18] br[17] br[16] br[15] br[14] br[13] br[12] br[11] br[10] br[9] br[8] br[7] br[6] br[5] br[4] br[3] br[2] br[1] br[0] data[31] data[30] data[29] data[28] data[27] data[26] data[25] data[24] data[23] data[22] data[21] data[20] data[19] data[18] data[17] data[16] data[15] data[14] data[13] data[12] data[11] data[10] data[9] data[8] data[7] data[6] data[5] data[4] data[3] data[2] data[1] data[0] data_b[31] data_b[30] data_b[29] data_b[28] data_b[27] data_b[26] data_b[25] data_b[24] data_b[23] data_b[22] data_b[21] data_b[20] data_b[19] data_b[18] data_b[17] data_b[16] data_b[15] data_b[14] data_b[13] data_b[12] data_b[11] data_b[10] data_b[9] data_b[8] data_b[7] data_b[6] data_b[5] data_b[4] data_b[3] data_b[2] data_b[1] data_b[0] 

xsense_amp_0 
+ clk br[0] bl[0] data_b[0] data[0] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_1 
+ clk br[1] bl[1] data_b[1] data[1] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_2 
+ clk br[2] bl[2] data_b[2] data[2] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_3 
+ clk br[3] bl[3] data_b[3] data[3] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_4 
+ clk br[4] bl[4] data_b[4] data[4] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_5 
+ clk br[5] bl[5] data_b[5] data[5] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_6 
+ clk br[6] bl[6] data_b[6] data[6] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_7 
+ clk br[7] bl[7] data_b[7] data[7] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_8 
+ clk br[8] bl[8] data_b[8] data[8] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_9 
+ clk br[9] bl[9] data_b[9] data[9] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_10 
+ clk br[10] bl[10] data_b[10] data[10] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_11 
+ clk br[11] bl[11] data_b[11] data[11] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_12 
+ clk br[12] bl[12] data_b[12] data[12] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_13 
+ clk br[13] bl[13] data_b[13] data[13] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_14 
+ clk br[14] bl[14] data_b[14] data[14] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_15 
+ clk br[15] bl[15] data_b[15] data[15] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_16 
+ clk br[16] bl[16] data_b[16] data[16] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_17 
+ clk br[17] bl[17] data_b[17] data[17] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_18 
+ clk br[18] bl[18] data_b[18] data[18] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_19 
+ clk br[19] bl[19] data_b[19] data[19] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_20 
+ clk br[20] bl[20] data_b[20] data[20] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_21 
+ clk br[21] bl[21] data_b[21] data[21] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_22 
+ clk br[22] bl[22] data_b[22] data[22] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_23 
+ clk br[23] bl[23] data_b[23] data[23] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_24 
+ clk br[24] bl[24] data_b[24] data[24] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_25 
+ clk br[25] bl[25] data_b[25] data[25] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_26 
+ clk br[26] bl[26] data_b[26] data[26] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_27 
+ clk br[27] bl[27] data_b[27] data[27] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_28 
+ clk br[28] bl[28] data_b[28] data[28] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_29 
+ clk br[29] bl[29] data_b[29] data[29] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_30 
+ clk br[30] bl[30] data_b[30] data[30] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_31 
+ clk br[31] bl[31] data_b[31] data[31] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

.ENDS

.SUBCKT dout_buf 
+ din1 din2 dout1 dout2 vdd vss 

xMP11 
+ x1 din1 vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='1.6' l='0.15' 

xMN11 
+ x1 din1 vss vss 
+ sky130_fd_pr__nfet_01v8 
+ w='1.0' l='0.15' 

xMP21 
+ dout1 x1 vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='3.2' l='0.15' 

xMN21 
+ dout1 x1 vss vss 
+ sky130_fd_pr__nfet_01v8 
+ w='2.0' l='0.15' 

xMP12 
+ x2 din2 vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='1.6' l='0.15' 

xMN12 
+ x2 din2 vss vss 
+ sky130_fd_pr__nfet_01v8 
+ w='1.0' l='0.15' 

xMP22 
+ dout2 x2 vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='3.2' l='0.15' 

xMN22 
+ dout2 x2 vss vss 
+ sky130_fd_pr__nfet_01v8 
+ w='2.0' l='0.15' 

.ENDS

.SUBCKT dout_buf_array 
+ din1[31] din1[30] din1[29] din1[28] din1[27] din1[26] din1[25] din1[24] din1[23] din1[22] din1[21] din1[20] din1[19] din1[18] din1[17] din1[16] din1[15] din1[14] din1[13] din1[12] din1[11] din1[10] din1[9] din1[8] din1[7] din1[6] din1[5] din1[4] din1[3] din1[2] din1[1] din1[0] din2[31] din2[30] din2[29] din2[28] din2[27] din2[26] din2[25] din2[24] din2[23] din2[22] din2[21] din2[20] din2[19] din2[18] din2[17] din2[16] din2[15] din2[14] din2[13] din2[12] din2[11] din2[10] din2[9] din2[8] din2[7] din2[6] din2[5] din2[4] din2[3] din2[2] din2[1] din2[0] dout1[31] dout1[30] dout1[29] dout1[28] dout1[27] dout1[26] dout1[25] dout1[24] dout1[23] dout1[22] dout1[21] dout1[20] dout1[19] dout1[18] dout1[17] dout1[16] dout1[15] dout1[14] dout1[13] dout1[12] dout1[11] dout1[10] dout1[9] dout1[8] dout1[7] dout1[6] dout1[5] dout1[4] dout1[3] dout1[2] dout1[1] dout1[0] dout2[31] dout2[30] dout2[29] dout2[28] dout2[27] dout2[26] dout2[25] dout2[24] dout2[23] dout2[22] dout2[21] dout2[20] dout2[19] dout2[18] dout2[17] dout2[16] dout2[15] dout2[14] dout2[13] dout2[12] dout2[11] dout2[10] dout2[9] dout2[8] dout2[7] dout2[6] dout2[5] dout2[4] dout2[3] dout2[2] dout2[1] dout2[0] vdd vss 

xbuf_0 
+ din1[0] din2[0] dout1[0] dout2[0] vdd vss 
+ dout_buf 
* No parameters

xbuf_1 
+ din1[1] din2[1] dout1[1] dout2[1] vdd vss 
+ dout_buf 
* No parameters

xbuf_2 
+ din1[2] din2[2] dout1[2] dout2[2] vdd vss 
+ dout_buf 
* No parameters

xbuf_3 
+ din1[3] din2[3] dout1[3] dout2[3] vdd vss 
+ dout_buf 
* No parameters

xbuf_4 
+ din1[4] din2[4] dout1[4] dout2[4] vdd vss 
+ dout_buf 
* No parameters

xbuf_5 
+ din1[5] din2[5] dout1[5] dout2[5] vdd vss 
+ dout_buf 
* No parameters

xbuf_6 
+ din1[6] din2[6] dout1[6] dout2[6] vdd vss 
+ dout_buf 
* No parameters

xbuf_7 
+ din1[7] din2[7] dout1[7] dout2[7] vdd vss 
+ dout_buf 
* No parameters

xbuf_8 
+ din1[8] din2[8] dout1[8] dout2[8] vdd vss 
+ dout_buf 
* No parameters

xbuf_9 
+ din1[9] din2[9] dout1[9] dout2[9] vdd vss 
+ dout_buf 
* No parameters

xbuf_10 
+ din1[10] din2[10] dout1[10] dout2[10] vdd vss 
+ dout_buf 
* No parameters

xbuf_11 
+ din1[11] din2[11] dout1[11] dout2[11] vdd vss 
+ dout_buf 
* No parameters

xbuf_12 
+ din1[12] din2[12] dout1[12] dout2[12] vdd vss 
+ dout_buf 
* No parameters

xbuf_13 
+ din1[13] din2[13] dout1[13] dout2[13] vdd vss 
+ dout_buf 
* No parameters

xbuf_14 
+ din1[14] din2[14] dout1[14] dout2[14] vdd vss 
+ dout_buf 
* No parameters

xbuf_15 
+ din1[15] din2[15] dout1[15] dout2[15] vdd vss 
+ dout_buf 
* No parameters

xbuf_16 
+ din1[16] din2[16] dout1[16] dout2[16] vdd vss 
+ dout_buf 
* No parameters

xbuf_17 
+ din1[17] din2[17] dout1[17] dout2[17] vdd vss 
+ dout_buf 
* No parameters

xbuf_18 
+ din1[18] din2[18] dout1[18] dout2[18] vdd vss 
+ dout_buf 
* No parameters

xbuf_19 
+ din1[19] din2[19] dout1[19] dout2[19] vdd vss 
+ dout_buf 
* No parameters

xbuf_20 
+ din1[20] din2[20] dout1[20] dout2[20] vdd vss 
+ dout_buf 
* No parameters

xbuf_21 
+ din1[21] din2[21] dout1[21] dout2[21] vdd vss 
+ dout_buf 
* No parameters

xbuf_22 
+ din1[22] din2[22] dout1[22] dout2[22] vdd vss 
+ dout_buf 
* No parameters

xbuf_23 
+ din1[23] din2[23] dout1[23] dout2[23] vdd vss 
+ dout_buf 
* No parameters

xbuf_24 
+ din1[24] din2[24] dout1[24] dout2[24] vdd vss 
+ dout_buf 
* No parameters

xbuf_25 
+ din1[25] din2[25] dout1[25] dout2[25] vdd vss 
+ dout_buf 
* No parameters

xbuf_26 
+ din1[26] din2[26] dout1[26] dout2[26] vdd vss 
+ dout_buf 
* No parameters

xbuf_27 
+ din1[27] din2[27] dout1[27] dout2[27] vdd vss 
+ dout_buf 
* No parameters

xbuf_28 
+ din1[28] din2[28] dout1[28] dout2[28] vdd vss 
+ dout_buf 
* No parameters

xbuf_29 
+ din1[29] din2[29] dout1[29] dout2[29] vdd vss 
+ dout_buf 
* No parameters

xbuf_30 
+ din1[30] din2[30] dout1[30] dout2[30] vdd vss 
+ dout_buf 
* No parameters

xbuf_31 
+ din1[31] din2[31] dout1[31] dout2[31] vdd vss 
+ dout_buf 
* No parameters

.ENDS

.SUBCKT we_control_and2_nand 
+ gnd vdd a b y 

xn1 
+ x a gnd gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='3.0' l='0.15' 

xn2 
+ y b x gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='3.0' l='0.15' 

xp1 
+ y a vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='4.0' l='0.15' 

xp2 
+ y b vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='4.0' l='0.15' 

.ENDS

.SUBCKT we_control_and2_inv 
+ gnd vdd din din_b 

xn 
+ din_b din gnd gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='8.0' l='0.15' 

xp 
+ din_b din vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='12.0' l='0.15' 

.ENDS

.SUBCKT we_control_and2 
+ a b y vdd vss 

xnand 
+ vss vdd a b tmp 
+ we_control_and2_nand 
* No parameters

xinv 
+ vss vdd tmp y 
+ we_control_and2_inv 
* No parameters

.ENDS

.SUBCKT we_control 
+ wr_en sel[7] sel[6] sel[5] sel[4] sel[3] sel[2] sel[1] sel[0] write_driver_en[7] write_driver_en[6] write_driver_en[5] write_driver_en[4] write_driver_en[3] write_driver_en[2] write_driver_en[1] write_driver_en[0] vdd vss 

xand2_0 
+ sel[0] wr_en write_driver_en[0] vdd vss 
+ we_control_and2 
* No parameters

xand2_1 
+ sel[1] wr_en write_driver_en[1] vdd vss 
+ we_control_and2 
* No parameters

xand2_2 
+ sel[2] wr_en write_driver_en[2] vdd vss 
+ we_control_and2 
* No parameters

xand2_3 
+ sel[3] wr_en write_driver_en[3] vdd vss 
+ we_control_and2 
* No parameters

xand2_4 
+ sel[4] wr_en write_driver_en[4] vdd vss 
+ we_control_and2 
* No parameters

xand2_5 
+ sel[5] wr_en write_driver_en[5] vdd vss 
+ we_control_and2 
* No parameters

xand2_6 
+ sel[6] wr_en write_driver_en[6] vdd vss 
+ we_control_and2 
* No parameters

xand2_7 
+ sel[7] wr_en write_driver_en[7] vdd vss 
+ we_control_and2 
* No parameters

.ENDS

.SUBCKT control_logic_delay_chain 
+ din dout vdd vss 

xinv_0 
+ din int[0] vdd vss 
+ control_logic_inv 
* No parameters

xinv_1 
+ int[0] int[1] vdd vss 
+ control_logic_inv 
* No parameters

xinv_2 
+ int[1] int[2] vdd vss 
+ control_logic_inv 
* No parameters

xinv_3 
+ int[2] int[3] vdd vss 
+ control_logic_inv 
* No parameters

xinv_4 
+ int[3] int[4] vdd vss 
+ control_logic_inv 
* No parameters

xinv_5 
+ int[4] int[5] vdd vss 
+ control_logic_inv 
* No parameters

xinv_6 
+ int[5] int[6] vdd vss 
+ control_logic_inv 
* No parameters

xinv_7 
+ int[6] int[7] vdd vss 
+ control_logic_inv 
* No parameters

xinv_8 
+ int[7] int[8] vdd vss 
+ control_logic_inv 
* No parameters

xinv_9 
+ int[8] int[9] vdd vss 
+ control_logic_inv 
* No parameters

xinv_10 
+ int[9] int[10] vdd vss 
+ control_logic_inv 
* No parameters

xinv_11 
+ int[10] int[11] vdd vss 
+ control_logic_inv 
* No parameters

xinv_12 
+ int[11] int[12] vdd vss 
+ control_logic_inv 
* No parameters

xinv_13 
+ int[12] int[13] vdd vss 
+ control_logic_inv 
* No parameters

xinv_14 
+ int[13] int[14] vdd vss 
+ control_logic_inv 
* No parameters

xinv_15 
+ int[14] int[15] vdd vss 
+ control_logic_inv 
* No parameters

xinv_16 
+ int[15] int[16] vdd vss 
+ control_logic_inv 
* No parameters

xinv_17 
+ int[16] int[17] vdd vss 
+ control_logic_inv 
* No parameters

xinv_18 
+ int[17] int[18] vdd vss 
+ control_logic_inv 
* No parameters

xinv_19 
+ int[18] int[19] vdd vss 
+ control_logic_inv 
* No parameters

xinv_20 
+ int[19] int[20] vdd vss 
+ control_logic_inv 
* No parameters

xinv_21 
+ int[20] int[21] vdd vss 
+ control_logic_inv 
* No parameters

xinv_22 
+ int[21] int[22] vdd vss 
+ control_logic_inv 
* No parameters

xinv_23 
+ int[22] int[23] vdd vss 
+ control_logic_inv 
* No parameters

xinv_24 
+ int[23] int[24] vdd vss 
+ control_logic_inv 
* No parameters

xinv_25 
+ int[24] int[25] vdd vss 
+ control_logic_inv 
* No parameters

xinv_26 
+ int[25] int[26] vdd vss 
+ control_logic_inv 
* No parameters

xinv_27 
+ int[26] int[27] vdd vss 
+ control_logic_inv 
* No parameters

xinv_28 
+ int[27] int[28] vdd vss 
+ control_logic_inv 
* No parameters

xinv_29 
+ int[28] int[29] vdd vss 
+ control_logic_inv 
* No parameters

xinv_30 
+ int[29] int[30] vdd vss 
+ control_logic_inv 
* No parameters

xinv_31 
+ int[30] int[31] vdd vss 
+ control_logic_inv 
* No parameters

xinv_32 
+ int[31] int[32] vdd vss 
+ control_logic_inv 
* No parameters

xinv_33 
+ int[32] int[33] vdd vss 
+ control_logic_inv 
* No parameters

xinv_34 
+ int[33] int[34] vdd vss 
+ control_logic_inv 
* No parameters

xinv_35 
+ int[34] int[35] vdd vss 
+ control_logic_inv 
* No parameters

xinv_36 
+ int[35] int[36] vdd vss 
+ control_logic_inv 
* No parameters

xinv_37 
+ int[36] int[37] vdd vss 
+ control_logic_inv 
* No parameters

xinv_38 
+ int[37] int[38] vdd vss 
+ control_logic_inv 
* No parameters

xinv_39 
+ int[38] int[39] vdd vss 
+ control_logic_inv 
* No parameters

xinv_40 
+ int[39] int[40] vdd vss 
+ control_logic_inv 
* No parameters

xinv_41 
+ int[40] int[41] vdd vss 
+ control_logic_inv 
* No parameters

xinv_42 
+ int[41] int[42] vdd vss 
+ control_logic_inv 
* No parameters

xinv_43 
+ int[42] int[43] vdd vss 
+ control_logic_inv 
* No parameters

xinv_44 
+ int[43] dout vdd vss 
+ control_logic_inv 
* No parameters

.ENDS

.SUBCKT sramgen_sram_1024x32m8w8_replica_v1 
+ vdd vss clk din[31] din[30] din[29] din[28] din[27] din[26] din[25] din[24] din[23] din[22] din[21] din[20] din[19] din[18] din[17] din[16] din[15] din[14] din[13] din[12] din[11] din[10] din[9] din[8] din[7] din[6] din[5] din[4] din[3] din[2] din[1] din[0] dout[31] dout[30] dout[29] dout[28] dout[27] dout[26] dout[25] dout[24] dout[23] dout[22] dout[21] dout[20] dout[19] dout[18] dout[17] dout[16] dout[15] dout[14] dout[13] dout[12] dout[11] dout[10] dout[9] dout[8] dout[7] dout[6] dout[5] dout[4] dout[3] dout[2] dout[1] dout[0] we addr[9] addr[8] addr[7] addr[6] addr[5] addr[4] addr[3] addr[2] addr[1] addr[0] wmask[3] wmask[2] wmask[1] wmask[0] 

xdin_dffs 
+ vdd vss clk din[31] din[30] din[29] din[28] din[27] din[26] din[25] din[24] din[23] din[22] din[21] din[20] din[19] din[18] din[17] din[16] din[15] din[14] din[13] din[12] din[11] din[10] din[9] din[8] din[7] din[6] din[5] din[4] din[3] din[2] din[1] din[0] bank_din[31] bank_din[30] bank_din[29] bank_din[28] bank_din[27] bank_din[26] bank_din[25] bank_din[24] bank_din[23] bank_din[22] bank_din[21] bank_din[20] bank_din[19] bank_din[18] bank_din[17] bank_din[16] bank_din[15] bank_din[14] bank_din[13] bank_din[12] bank_din[11] bank_din[10] bank_din[9] bank_din[8] bank_din[7] bank_din[6] bank_din[5] bank_din[4] bank_din[3] bank_din[2] bank_din[1] bank_din[0] dff_din_b[31] dff_din_b[30] dff_din_b[29] dff_din_b[28] dff_din_b[27] dff_din_b[26] dff_din_b[25] dff_din_b[24] dff_din_b[23] dff_din_b[22] dff_din_b[21] dff_din_b[20] dff_din_b[19] dff_din_b[18] dff_din_b[17] dff_din_b[16] dff_din_b[15] dff_din_b[14] dff_din_b[13] dff_din_b[12] dff_din_b[11] dff_din_b[10] dff_din_b[9] dff_din_b[8] dff_din_b[7] dff_din_b[6] dff_din_b[5] dff_din_b[4] dff_din_b[3] dff_din_b[2] dff_din_b[1] dff_din_b[0] 
+ data_dff_array 
* No parameters

xaddr_dffs 
+ vdd vss clk addr[9] addr[8] addr[7] addr[6] addr[5] addr[4] addr[3] addr[2] addr[1] addr[0] bank_addr[9] bank_addr[8] bank_addr[7] bank_addr[6] bank_addr[5] bank_addr[4] bank_addr[3] bank_addr[2] bank_addr[1] bank_addr[0] bank_addr_b[9] bank_addr_b[8] bank_addr_b[7] bank_addr_b[6] bank_addr_b[5] bank_addr_b[4] bank_addr_b[3] bank_addr_b[2] bank_addr_b[1] bank_addr_b[0] 
+ addr_dff_array 
* No parameters

xwmask_dffs 
+ vdd vss clk wmask[3] wmask[2] wmask[1] wmask[0] bank_wmask[3] bank_wmask[2] bank_wmask[1] bank_wmask[0] bank_wmask_b[3] bank_wmask_b[2] bank_wmask_b[1] bank_wmask_b[0] 
+ wmask_dff_array 
* No parameters

xwe_dff 
+ vdd vss clk we bank_we bank_we_b 
+ openram_dff 
* No parameters

xdecoder 
+ vdd vss bank_addr[9] bank_addr[8] bank_addr[7] bank_addr[6] bank_addr[5] bank_addr[4] bank_addr[3] bank_addr_b[9] bank_addr_b[8] bank_addr_b[7] bank_addr_b[6] bank_addr_b[5] bank_addr_b[4] bank_addr_b[3] wl_data[127] wl_data[126] wl_data[125] wl_data[124] wl_data[123] wl_data[122] wl_data[121] wl_data[120] wl_data[119] wl_data[118] wl_data[117] wl_data[116] wl_data[115] wl_data[114] wl_data[113] wl_data[112] wl_data[111] wl_data[110] wl_data[109] wl_data[108] wl_data[107] wl_data[106] wl_data[105] wl_data[104] wl_data[103] wl_data[102] wl_data[101] wl_data[100] wl_data[99] wl_data[98] wl_data[97] wl_data[96] wl_data[95] wl_data[94] wl_data[93] wl_data[92] wl_data[91] wl_data[90] wl_data[89] wl_data[88] wl_data[87] wl_data[86] wl_data[85] wl_data[84] wl_data[83] wl_data[82] wl_data[81] wl_data[80] wl_data[79] wl_data[78] wl_data[77] wl_data[76] wl_data[75] wl_data[74] wl_data[73] wl_data[72] wl_data[71] wl_data[70] wl_data[69] wl_data[68] wl_data[67] wl_data[66] wl_data[65] wl_data[64] wl_data[63] wl_data[62] wl_data[61] wl_data[60] wl_data[59] wl_data[58] wl_data[57] wl_data[56] wl_data[55] wl_data[54] wl_data[53] wl_data[52] wl_data[51] wl_data[50] wl_data[49] wl_data[48] wl_data[47] wl_data[46] wl_data[45] wl_data[44] wl_data[43] wl_data[42] wl_data[41] wl_data[40] wl_data[39] wl_data[38] wl_data[37] wl_data[36] wl_data[35] wl_data[34] wl_data[33] wl_data[32] wl_data[31] wl_data[30] wl_data[29] wl_data[28] wl_data[27] wl_data[26] wl_data[25] wl_data[24] wl_data[23] wl_data[22] wl_data[21] wl_data[20] wl_data[19] wl_data[18] wl_data[17] wl_data[16] wl_data[15] wl_data[14] wl_data[13] wl_data[12] wl_data[11] wl_data[10] wl_data[9] wl_data[8] wl_data[7] wl_data[6] wl_data[5] wl_data[4] wl_data[3] wl_data[2] wl_data[1] wl_data[0] wl_data_b[127] wl_data_b[126] wl_data_b[125] wl_data_b[124] wl_data_b[123] wl_data_b[122] wl_data_b[121] wl_data_b[120] wl_data_b[119] wl_data_b[118] wl_data_b[117] wl_data_b[116] wl_data_b[115] wl_data_b[114] wl_data_b[113] wl_data_b[112] wl_data_b[111] wl_data_b[110] wl_data_b[109] wl_data_b[108] wl_data_b[107] wl_data_b[106] wl_data_b[105] wl_data_b[104] wl_data_b[103] wl_data_b[102] wl_data_b[101] wl_data_b[100] wl_data_b[99] wl_data_b[98] wl_data_b[97] wl_data_b[96] wl_data_b[95] wl_data_b[94] wl_data_b[93] wl_data_b[92] wl_data_b[91] wl_data_b[90] wl_data_b[89] wl_data_b[88] wl_data_b[87] wl_data_b[86] wl_data_b[85] wl_data_b[84] wl_data_b[83] wl_data_b[82] wl_data_b[81] wl_data_b[80] wl_data_b[79] wl_data_b[78] wl_data_b[77] wl_data_b[76] wl_data_b[75] wl_data_b[74] wl_data_b[73] wl_data_b[72] wl_data_b[71] wl_data_b[70] wl_data_b[69] wl_data_b[68] wl_data_b[67] wl_data_b[66] wl_data_b[65] wl_data_b[64] wl_data_b[63] wl_data_b[62] wl_data_b[61] wl_data_b[60] wl_data_b[59] wl_data_b[58] wl_data_b[57] wl_data_b[56] wl_data_b[55] wl_data_b[54] wl_data_b[53] wl_data_b[52] wl_data_b[51] wl_data_b[50] wl_data_b[49] wl_data_b[48] wl_data_b[47] wl_data_b[46] wl_data_b[45] wl_data_b[44] wl_data_b[43] wl_data_b[42] wl_data_b[41] wl_data_b[40] wl_data_b[39] wl_data_b[38] wl_data_b[37] wl_data_b[36] wl_data_b[35] wl_data_b[34] wl_data_b[33] wl_data_b[32] wl_data_b[31] wl_data_b[30] wl_data_b[29] wl_data_b[28] wl_data_b[27] wl_data_b[26] wl_data_b[25] wl_data_b[24] wl_data_b[23] wl_data_b[22] wl_data_b[21] wl_data_b[20] wl_data_b[19] wl_data_b[18] wl_data_b[17] wl_data_b[16] wl_data_b[15] wl_data_b[14] wl_data_b[13] wl_data_b[12] wl_data_b[11] wl_data_b[10] wl_data_b[9] wl_data_b[8] wl_data_b[7] wl_data_b[6] wl_data_b[5] wl_data_b[4] wl_data_b[3] wl_data_b[2] wl_data_b[1] wl_data_b[0] 
+ hierarchical_decoder 
* No parameters

xwl_driver_array 
+ vdd vss wl_data[127] wl_data[126] wl_data[125] wl_data[124] wl_data[123] wl_data[122] wl_data[121] wl_data[120] wl_data[119] wl_data[118] wl_data[117] wl_data[116] wl_data[115] wl_data[114] wl_data[113] wl_data[112] wl_data[111] wl_data[110] wl_data[109] wl_data[108] wl_data[107] wl_data[106] wl_data[105] wl_data[104] wl_data[103] wl_data[102] wl_data[101] wl_data[100] wl_data[99] wl_data[98] wl_data[97] wl_data[96] wl_data[95] wl_data[94] wl_data[93] wl_data[92] wl_data[91] wl_data[90] wl_data[89] wl_data[88] wl_data[87] wl_data[86] wl_data[85] wl_data[84] wl_data[83] wl_data[82] wl_data[81] wl_data[80] wl_data[79] wl_data[78] wl_data[77] wl_data[76] wl_data[75] wl_data[74] wl_data[73] wl_data[72] wl_data[71] wl_data[70] wl_data[69] wl_data[68] wl_data[67] wl_data[66] wl_data[65] wl_data[64] wl_data[63] wl_data[62] wl_data[61] wl_data[60] wl_data[59] wl_data[58] wl_data[57] wl_data[56] wl_data[55] wl_data[54] wl_data[53] wl_data[52] wl_data[51] wl_data[50] wl_data[49] wl_data[48] wl_data[47] wl_data[46] wl_data[45] wl_data[44] wl_data[43] wl_data[42] wl_data[41] wl_data[40] wl_data[39] wl_data[38] wl_data[37] wl_data[36] wl_data[35] wl_data[34] wl_data[33] wl_data[32] wl_data[31] wl_data[30] wl_data[29] wl_data[28] wl_data[27] wl_data[26] wl_data[25] wl_data[24] wl_data[23] wl_data[22] wl_data[21] wl_data[20] wl_data[19] wl_data[18] wl_data[17] wl_data[16] wl_data[15] wl_data[14] wl_data[13] wl_data[12] wl_data[11] wl_data[10] wl_data[9] wl_data[8] wl_data[7] wl_data[6] wl_data[5] wl_data[4] wl_data[3] wl_data[2] wl_data[1] wl_data[0] wl_en wl[127] wl[126] wl[125] wl[124] wl[123] wl[122] wl[121] wl[120] wl[119] wl[118] wl[117] wl[116] wl[115] wl[114] wl[113] wl[112] wl[111] wl[110] wl[109] wl[108] wl[107] wl[106] wl[105] wl[104] wl[103] wl[102] wl[101] wl[100] wl[99] wl[98] wl[97] wl[96] wl[95] wl[94] wl[93] wl[92] wl[91] wl[90] wl[89] wl[88] wl[87] wl[86] wl[85] wl[84] wl[83] wl[82] wl[81] wl[80] wl[79] wl[78] wl[77] wl[76] wl[75] wl[74] wl[73] wl[72] wl[71] wl[70] wl[69] wl[68] wl[67] wl[66] wl[65] wl[64] wl[63] wl[62] wl[61] wl[60] wl[59] wl[58] wl[57] wl[56] wl[55] wl[54] wl[53] wl[52] wl[51] wl[50] wl[49] wl[48] wl[47] wl[46] wl[45] wl[44] wl[43] wl[42] wl[41] wl[40] wl[39] wl[38] wl[37] wl[36] wl[35] wl[34] wl[33] wl[32] wl[31] wl[30] wl[29] wl[28] wl[27] wl[26] wl[25] wl[24] wl[23] wl[22] wl[21] wl[20] wl[19] wl[18] wl[17] wl[16] wl[15] wl[14] wl[13] wl[12] wl[11] wl[10] wl[9] wl[8] wl[7] wl[6] wl[5] wl[4] wl[3] wl[2] wl[1] wl[0] 
+ wordline_driver_array 
* No parameters

xbitcells 
+ vdd vss bl[255] bl[254] bl[253] bl[252] bl[251] bl[250] bl[249] bl[248] bl[247] bl[246] bl[245] bl[244] bl[243] bl[242] bl[241] bl[240] bl[239] bl[238] bl[237] bl[236] bl[235] bl[234] bl[233] bl[232] bl[231] bl[230] bl[229] bl[228] bl[227] bl[226] bl[225] bl[224] bl[223] bl[222] bl[221] bl[220] bl[219] bl[218] bl[217] bl[216] bl[215] bl[214] bl[213] bl[212] bl[211] bl[210] bl[209] bl[208] bl[207] bl[206] bl[205] bl[204] bl[203] bl[202] bl[201] bl[200] bl[199] bl[198] bl[197] bl[196] bl[195] bl[194] bl[193] bl[192] bl[191] bl[190] bl[189] bl[188] bl[187] bl[186] bl[185] bl[184] bl[183] bl[182] bl[181] bl[180] bl[179] bl[178] bl[177] bl[176] bl[175] bl[174] bl[173] bl[172] bl[171] bl[170] bl[169] bl[168] bl[167] bl[166] bl[165] bl[164] bl[163] bl[162] bl[161] bl[160] bl[159] bl[158] bl[157] bl[156] bl[155] bl[154] bl[153] bl[152] bl[151] bl[150] bl[149] bl[148] bl[147] bl[146] bl[145] bl[144] bl[143] bl[142] bl[141] bl[140] bl[139] bl[138] bl[137] bl[136] bl[135] bl[134] bl[133] bl[132] bl[131] bl[130] bl[129] bl[128] bl[127] bl[126] bl[125] bl[124] bl[123] bl[122] bl[121] bl[120] bl[119] bl[118] bl[117] bl[116] bl[115] bl[114] bl[113] bl[112] bl[111] bl[110] bl[109] bl[108] bl[107] bl[106] bl[105] bl[104] bl[103] bl[102] bl[101] bl[100] bl[99] bl[98] bl[97] bl[96] bl[95] bl[94] bl[93] bl[92] bl[91] bl[90] bl[89] bl[88] bl[87] bl[86] bl[85] bl[84] bl[83] bl[82] bl[81] bl[80] bl[79] bl[78] bl[77] bl[76] bl[75] bl[74] bl[73] bl[72] bl[71] bl[70] bl[69] bl[68] bl[67] bl[66] bl[65] bl[64] bl[63] bl[62] bl[61] bl[60] bl[59] bl[58] bl[57] bl[56] bl[55] bl[54] bl[53] bl[52] bl[51] bl[50] bl[49] bl[48] bl[47] bl[46] bl[45] bl[44] bl[43] bl[42] bl[41] bl[40] bl[39] bl[38] bl[37] bl[36] bl[35] bl[34] bl[33] bl[32] bl[31] bl[30] bl[29] bl[28] bl[27] bl[26] bl[25] bl[24] bl[23] bl[22] bl[21] bl[20] bl[19] bl[18] bl[17] bl[16] bl[15] bl[14] bl[13] bl[12] bl[11] bl[10] bl[9] bl[8] bl[7] bl[6] bl[5] bl[4] bl[3] bl[2] bl[1] bl[0] br[255] br[254] br[253] br[252] br[251] br[250] br[249] br[248] br[247] br[246] br[245] br[244] br[243] br[242] br[241] br[240] br[239] br[238] br[237] br[236] br[235] br[234] br[233] br[232] br[231] br[230] br[229] br[228] br[227] br[226] br[225] br[224] br[223] br[222] br[221] br[220] br[219] br[218] br[217] br[216] br[215] br[214] br[213] br[212] br[211] br[210] br[209] br[208] br[207] br[206] br[205] br[204] br[203] br[202] br[201] br[200] br[199] br[198] br[197] br[196] br[195] br[194] br[193] br[192] br[191] br[190] br[189] br[188] br[187] br[186] br[185] br[184] br[183] br[182] br[181] br[180] br[179] br[178] br[177] br[176] br[175] br[174] br[173] br[172] br[171] br[170] br[169] br[168] br[167] br[166] br[165] br[164] br[163] br[162] br[161] br[160] br[159] br[158] br[157] br[156] br[155] br[154] br[153] br[152] br[151] br[150] br[149] br[148] br[147] br[146] br[145] br[144] br[143] br[142] br[141] br[140] br[139] br[138] br[137] br[136] br[135] br[134] br[133] br[132] br[131] br[130] br[129] br[128] br[127] br[126] br[125] br[124] br[123] br[122] br[121] br[120] br[119] br[118] br[117] br[116] br[115] br[114] br[113] br[112] br[111] br[110] br[109] br[108] br[107] br[106] br[105] br[104] br[103] br[102] br[101] br[100] br[99] br[98] br[97] br[96] br[95] br[94] br[93] br[92] br[91] br[90] br[89] br[88] br[87] br[86] br[85] br[84] br[83] br[82] br[81] br[80] br[79] br[78] br[77] br[76] br[75] br[74] br[73] br[72] br[71] br[70] br[69] br[68] br[67] br[66] br[65] br[64] br[63] br[62] br[61] br[60] br[59] br[58] br[57] br[56] br[55] br[54] br[53] br[52] br[51] br[50] br[49] br[48] br[47] br[46] br[45] br[44] br[43] br[42] br[41] br[40] br[39] br[38] br[37] br[36] br[35] br[34] br[33] br[32] br[31] br[30] br[29] br[28] br[27] br[26] br[25] br[24] br[23] br[22] br[21] br[20] br[19] br[18] br[17] br[16] br[15] br[14] br[13] br[12] br[11] br[10] br[9] br[8] br[7] br[6] br[5] br[4] br[3] br[2] br[1] br[0] wl[127] wl[126] wl[125] wl[124] wl[123] wl[122] wl[121] wl[120] wl[119] wl[118] wl[117] wl[116] wl[115] wl[114] wl[113] wl[112] wl[111] wl[110] wl[109] wl[108] wl[107] wl[106] wl[105] wl[104] wl[103] wl[102] wl[101] wl[100] wl[99] wl[98] wl[97] wl[96] wl[95] wl[94] wl[93] wl[92] wl[91] wl[90] wl[89] wl[88] wl[87] wl[86] wl[85] wl[84] wl[83] wl[82] wl[81] wl[80] wl[79] wl[78] wl[77] wl[76] wl[75] wl[74] wl[73] wl[72] wl[71] wl[70] wl[69] wl[68] wl[67] wl[66] wl[65] wl[64] wl[63] wl[62] wl[61] wl[60] wl[59] wl[58] wl[57] wl[56] wl[55] wl[54] wl[53] wl[52] wl[51] wl[50] wl[49] wl[48] wl[47] wl[46] wl[45] wl[44] wl[43] wl[42] wl[41] wl[40] wl[39] wl[38] wl[37] wl[36] wl[35] wl[34] wl[33] wl[32] wl[31] wl[30] wl[29] wl[28] wl[27] wl[26] wl[25] wl[24] wl[23] wl[22] wl[21] wl[20] wl[19] wl[18] wl[17] wl[16] wl[15] wl[14] wl[13] wl[12] wl[11] wl[10] wl[9] wl[8] wl[7] wl[6] wl[5] wl[4] wl[3] wl[2] wl[1] wl[0] vss vdd rbl rbr 
+ bitcell_array 
* No parameters

xprecharge_array 
+ vdd pc_b rbl bl[255] bl[254] bl[253] bl[252] bl[251] bl[250] bl[249] bl[248] bl[247] bl[246] bl[245] bl[244] bl[243] bl[242] bl[241] bl[240] bl[239] bl[238] bl[237] bl[236] bl[235] bl[234] bl[233] bl[232] bl[231] bl[230] bl[229] bl[228] bl[227] bl[226] bl[225] bl[224] bl[223] bl[222] bl[221] bl[220] bl[219] bl[218] bl[217] bl[216] bl[215] bl[214] bl[213] bl[212] bl[211] bl[210] bl[209] bl[208] bl[207] bl[206] bl[205] bl[204] bl[203] bl[202] bl[201] bl[200] bl[199] bl[198] bl[197] bl[196] bl[195] bl[194] bl[193] bl[192] bl[191] bl[190] bl[189] bl[188] bl[187] bl[186] bl[185] bl[184] bl[183] bl[182] bl[181] bl[180] bl[179] bl[178] bl[177] bl[176] bl[175] bl[174] bl[173] bl[172] bl[171] bl[170] bl[169] bl[168] bl[167] bl[166] bl[165] bl[164] bl[163] bl[162] bl[161] bl[160] bl[159] bl[158] bl[157] bl[156] bl[155] bl[154] bl[153] bl[152] bl[151] bl[150] bl[149] bl[148] bl[147] bl[146] bl[145] bl[144] bl[143] bl[142] bl[141] bl[140] bl[139] bl[138] bl[137] bl[136] bl[135] bl[134] bl[133] bl[132] bl[131] bl[130] bl[129] bl[128] bl[127] bl[126] bl[125] bl[124] bl[123] bl[122] bl[121] bl[120] bl[119] bl[118] bl[117] bl[116] bl[115] bl[114] bl[113] bl[112] bl[111] bl[110] bl[109] bl[108] bl[107] bl[106] bl[105] bl[104] bl[103] bl[102] bl[101] bl[100] bl[99] bl[98] bl[97] bl[96] bl[95] bl[94] bl[93] bl[92] bl[91] bl[90] bl[89] bl[88] bl[87] bl[86] bl[85] bl[84] bl[83] bl[82] bl[81] bl[80] bl[79] bl[78] bl[77] bl[76] bl[75] bl[74] bl[73] bl[72] bl[71] bl[70] bl[69] bl[68] bl[67] bl[66] bl[65] bl[64] bl[63] bl[62] bl[61] bl[60] bl[59] bl[58] bl[57] bl[56] bl[55] bl[54] bl[53] bl[52] bl[51] bl[50] bl[49] bl[48] bl[47] bl[46] bl[45] bl[44] bl[43] bl[42] bl[41] bl[40] bl[39] bl[38] bl[37] bl[36] bl[35] bl[34] bl[33] bl[32] bl[31] bl[30] bl[29] bl[28] bl[27] bl[26] bl[25] bl[24] bl[23] bl[22] bl[21] bl[20] bl[19] bl[18] bl[17] bl[16] bl[15] bl[14] bl[13] bl[12] bl[11] bl[10] bl[9] bl[8] bl[7] bl[6] bl[5] bl[4] bl[3] bl[2] bl[1] bl[0]  rbr br[255] br[254] br[253] br[252] br[251] br[250] br[249] br[248] br[247] br[246] br[245] br[244] br[243] br[242] br[241] br[240] br[239] br[238] br[237] br[236] br[235] br[234] br[233] br[232] br[231] br[230] br[229] br[228] br[227] br[226] br[225] br[224] br[223] br[222] br[221] br[220] br[219] br[218] br[217] br[216] br[215] br[214] br[213] br[212] br[211] br[210] br[209] br[208] br[207] br[206] br[205] br[204] br[203] br[202] br[201] br[200] br[199] br[198] br[197] br[196] br[195] br[194] br[193] br[192] br[191] br[190] br[189] br[188] br[187] br[186] br[185] br[184] br[183] br[182] br[181] br[180] br[179] br[178] br[177] br[176] br[175] br[174] br[173] br[172] br[171] br[170] br[169] br[168] br[167] br[166] br[165] br[164] br[163] br[162] br[161] br[160] br[159] br[158] br[157] br[156] br[155] br[154] br[153] br[152] br[151] br[150] br[149] br[148] br[147] br[146] br[145] br[144] br[143] br[142] br[141] br[140] br[139] br[138] br[137] br[136] br[135] br[134] br[133] br[132] br[131] br[130] br[129] br[128] br[127] br[126] br[125] br[124] br[123] br[122] br[121] br[120] br[119] br[118] br[117] br[116] br[115] br[114] br[113] br[112] br[111] br[110] br[109] br[108] br[107] br[106] br[105] br[104] br[103] br[102] br[101] br[100] br[99] br[98] br[97] br[96] br[95] br[94] br[93] br[92] br[91] br[90] br[89] br[88] br[87] br[86] br[85] br[84] br[83] br[82] br[81] br[80] br[79] br[78] br[77] br[76] br[75] br[74] br[73] br[72] br[71] br[70] br[69] br[68] br[67] br[66] br[65] br[64] br[63] br[62] br[61] br[60] br[59] br[58] br[57] br[56] br[55] br[54] br[53] br[52] br[51] br[50] br[49] br[48] br[47] br[46] br[45] br[44] br[43] br[42] br[41] br[40] br[39] br[38] br[37] br[36] br[35] br[34] br[33] br[32] br[31] br[30] br[29] br[28] br[27] br[26] br[25] br[24] br[23] br[22] br[21] br[20] br[19] br[18] br[17] br[16] br[15] br[14] br[13] br[12] br[11] br[10] br[9] br[8] br[7] br[6] br[5] br[4] br[3] br[2] br[1] br[0]  
+ precharge_array 
* No parameters

xwrite_mux_array 
+ write_driver_en[7] write_driver_en[6] write_driver_en[5] write_driver_en[4] write_driver_en[3] write_driver_en[2] write_driver_en[1] write_driver_en[0] bank_wmask[3] bank_wmask[2] bank_wmask[1] bank_wmask[0] bank_din[31] bank_din[30] bank_din[29] bank_din[28] bank_din[27] bank_din[26] bank_din[25] bank_din[24] bank_din[23] bank_din[22] bank_din[21] bank_din[20] bank_din[19] bank_din[18] bank_din[17] bank_din[16] bank_din[15] bank_din[14] bank_din[13] bank_din[12] bank_din[11] bank_din[10] bank_din[9] bank_din[8] bank_din[7] bank_din[6] bank_din[5] bank_din[4] bank_din[3] bank_din[2] bank_din[1] bank_din[0] bank_din_b[31] bank_din_b[30] bank_din_b[29] bank_din_b[28] bank_din_b[27] bank_din_b[26] bank_din_b[25] bank_din_b[24] bank_din_b[23] bank_din_b[22] bank_din_b[21] bank_din_b[20] bank_din_b[19] bank_din_b[18] bank_din_b[17] bank_din_b[16] bank_din_b[15] bank_din_b[14] bank_din_b[13] bank_din_b[12] bank_din_b[11] bank_din_b[10] bank_din_b[9] bank_din_b[8] bank_din_b[7] bank_din_b[6] bank_din_b[5] bank_din_b[4] bank_din_b[3] bank_din_b[2] bank_din_b[1] bank_din_b[0] bl[255] bl[254] bl[253] bl[252] bl[251] bl[250] bl[249] bl[248] bl[247] bl[246] bl[245] bl[244] bl[243] bl[242] bl[241] bl[240] bl[239] bl[238] bl[237] bl[236] bl[235] bl[234] bl[233] bl[232] bl[231] bl[230] bl[229] bl[228] bl[227] bl[226] bl[225] bl[224] bl[223] bl[222] bl[221] bl[220] bl[219] bl[218] bl[217] bl[216] bl[215] bl[214] bl[213] bl[212] bl[211] bl[210] bl[209] bl[208] bl[207] bl[206] bl[205] bl[204] bl[203] bl[202] bl[201] bl[200] bl[199] bl[198] bl[197] bl[196] bl[195] bl[194] bl[193] bl[192] bl[191] bl[190] bl[189] bl[188] bl[187] bl[186] bl[185] bl[184] bl[183] bl[182] bl[181] bl[180] bl[179] bl[178] bl[177] bl[176] bl[175] bl[174] bl[173] bl[172] bl[171] bl[170] bl[169] bl[168] bl[167] bl[166] bl[165] bl[164] bl[163] bl[162] bl[161] bl[160] bl[159] bl[158] bl[157] bl[156] bl[155] bl[154] bl[153] bl[152] bl[151] bl[150] bl[149] bl[148] bl[147] bl[146] bl[145] bl[144] bl[143] bl[142] bl[141] bl[140] bl[139] bl[138] bl[137] bl[136] bl[135] bl[134] bl[133] bl[132] bl[131] bl[130] bl[129] bl[128] bl[127] bl[126] bl[125] bl[124] bl[123] bl[122] bl[121] bl[120] bl[119] bl[118] bl[117] bl[116] bl[115] bl[114] bl[113] bl[112] bl[111] bl[110] bl[109] bl[108] bl[107] bl[106] bl[105] bl[104] bl[103] bl[102] bl[101] bl[100] bl[99] bl[98] bl[97] bl[96] bl[95] bl[94] bl[93] bl[92] bl[91] bl[90] bl[89] bl[88] bl[87] bl[86] bl[85] bl[84] bl[83] bl[82] bl[81] bl[80] bl[79] bl[78] bl[77] bl[76] bl[75] bl[74] bl[73] bl[72] bl[71] bl[70] bl[69] bl[68] bl[67] bl[66] bl[65] bl[64] bl[63] bl[62] bl[61] bl[60] bl[59] bl[58] bl[57] bl[56] bl[55] bl[54] bl[53] bl[52] bl[51] bl[50] bl[49] bl[48] bl[47] bl[46] bl[45] bl[44] bl[43] bl[42] bl[41] bl[40] bl[39] bl[38] bl[37] bl[36] bl[35] bl[34] bl[33] bl[32] bl[31] bl[30] bl[29] bl[28] bl[27] bl[26] bl[25] bl[24] bl[23] bl[22] bl[21] bl[20] bl[19] bl[18] bl[17] bl[16] bl[15] bl[14] bl[13] bl[12] bl[11] bl[10] bl[9] bl[8] bl[7] bl[6] bl[5] bl[4] bl[3] bl[2] bl[1] bl[0] br[255] br[254] br[253] br[252] br[251] br[250] br[249] br[248] br[247] br[246] br[245] br[244] br[243] br[242] br[241] br[240] br[239] br[238] br[237] br[236] br[235] br[234] br[233] br[232] br[231] br[230] br[229] br[228] br[227] br[226] br[225] br[224] br[223] br[222] br[221] br[220] br[219] br[218] br[217] br[216] br[215] br[214] br[213] br[212] br[211] br[210] br[209] br[208] br[207] br[206] br[205] br[204] br[203] br[202] br[201] br[200] br[199] br[198] br[197] br[196] br[195] br[194] br[193] br[192] br[191] br[190] br[189] br[188] br[187] br[186] br[185] br[184] br[183] br[182] br[181] br[180] br[179] br[178] br[177] br[176] br[175] br[174] br[173] br[172] br[171] br[170] br[169] br[168] br[167] br[166] br[165] br[164] br[163] br[162] br[161] br[160] br[159] br[158] br[157] br[156] br[155] br[154] br[153] br[152] br[151] br[150] br[149] br[148] br[147] br[146] br[145] br[144] br[143] br[142] br[141] br[140] br[139] br[138] br[137] br[136] br[135] br[134] br[133] br[132] br[131] br[130] br[129] br[128] br[127] br[126] br[125] br[124] br[123] br[122] br[121] br[120] br[119] br[118] br[117] br[116] br[115] br[114] br[113] br[112] br[111] br[110] br[109] br[108] br[107] br[106] br[105] br[104] br[103] br[102] br[101] br[100] br[99] br[98] br[97] br[96] br[95] br[94] br[93] br[92] br[91] br[90] br[89] br[88] br[87] br[86] br[85] br[84] br[83] br[82] br[81] br[80] br[79] br[78] br[77] br[76] br[75] br[74] br[73] br[72] br[71] br[70] br[69] br[68] br[67] br[66] br[65] br[64] br[63] br[62] br[61] br[60] br[59] br[58] br[57] br[56] br[55] br[54] br[53] br[52] br[51] br[50] br[49] br[48] br[47] br[46] br[45] br[44] br[43] br[42] br[41] br[40] br[39] br[38] br[37] br[36] br[35] br[34] br[33] br[32] br[31] br[30] br[29] br[28] br[27] br[26] br[25] br[24] br[23] br[22] br[21] br[20] br[19] br[18] br[17] br[16] br[15] br[14] br[13] br[12] br[11] br[10] br[9] br[8] br[7] br[6] br[5] br[4] br[3] br[2] br[1] br[0] vss 
+ write_mux_array 
* No parameters

xread_mux_array 
+ col_sel_b[7] col_sel_b[6] col_sel_b[5] col_sel_b[4] col_sel_b[3] col_sel_b[2] col_sel_b[1] col_sel_b[0] bl[255] bl[254] bl[253] bl[252] bl[251] bl[250] bl[249] bl[248] bl[247] bl[246] bl[245] bl[244] bl[243] bl[242] bl[241] bl[240] bl[239] bl[238] bl[237] bl[236] bl[235] bl[234] bl[233] bl[232] bl[231] bl[230] bl[229] bl[228] bl[227] bl[226] bl[225] bl[224] bl[223] bl[222] bl[221] bl[220] bl[219] bl[218] bl[217] bl[216] bl[215] bl[214] bl[213] bl[212] bl[211] bl[210] bl[209] bl[208] bl[207] bl[206] bl[205] bl[204] bl[203] bl[202] bl[201] bl[200] bl[199] bl[198] bl[197] bl[196] bl[195] bl[194] bl[193] bl[192] bl[191] bl[190] bl[189] bl[188] bl[187] bl[186] bl[185] bl[184] bl[183] bl[182] bl[181] bl[180] bl[179] bl[178] bl[177] bl[176] bl[175] bl[174] bl[173] bl[172] bl[171] bl[170] bl[169] bl[168] bl[167] bl[166] bl[165] bl[164] bl[163] bl[162] bl[161] bl[160] bl[159] bl[158] bl[157] bl[156] bl[155] bl[154] bl[153] bl[152] bl[151] bl[150] bl[149] bl[148] bl[147] bl[146] bl[145] bl[144] bl[143] bl[142] bl[141] bl[140] bl[139] bl[138] bl[137] bl[136] bl[135] bl[134] bl[133] bl[132] bl[131] bl[130] bl[129] bl[128] bl[127] bl[126] bl[125] bl[124] bl[123] bl[122] bl[121] bl[120] bl[119] bl[118] bl[117] bl[116] bl[115] bl[114] bl[113] bl[112] bl[111] bl[110] bl[109] bl[108] bl[107] bl[106] bl[105] bl[104] bl[103] bl[102] bl[101] bl[100] bl[99] bl[98] bl[97] bl[96] bl[95] bl[94] bl[93] bl[92] bl[91] bl[90] bl[89] bl[88] bl[87] bl[86] bl[85] bl[84] bl[83] bl[82] bl[81] bl[80] bl[79] bl[78] bl[77] bl[76] bl[75] bl[74] bl[73] bl[72] bl[71] bl[70] bl[69] bl[68] bl[67] bl[66] bl[65] bl[64] bl[63] bl[62] bl[61] bl[60] bl[59] bl[58] bl[57] bl[56] bl[55] bl[54] bl[53] bl[52] bl[51] bl[50] bl[49] bl[48] bl[47] bl[46] bl[45] bl[44] bl[43] bl[42] bl[41] bl[40] bl[39] bl[38] bl[37] bl[36] bl[35] bl[34] bl[33] bl[32] bl[31] bl[30] bl[29] bl[28] bl[27] bl[26] bl[25] bl[24] bl[23] bl[22] bl[21] bl[20] bl[19] bl[18] bl[17] bl[16] bl[15] bl[14] bl[13] bl[12] bl[11] bl[10] bl[9] bl[8] bl[7] bl[6] bl[5] bl[4] bl[3] bl[2] bl[1] bl[0] br[255] br[254] br[253] br[252] br[251] br[250] br[249] br[248] br[247] br[246] br[245] br[244] br[243] br[242] br[241] br[240] br[239] br[238] br[237] br[236] br[235] br[234] br[233] br[232] br[231] br[230] br[229] br[228] br[227] br[226] br[225] br[224] br[223] br[222] br[221] br[220] br[219] br[218] br[217] br[216] br[215] br[214] br[213] br[212] br[211] br[210] br[209] br[208] br[207] br[206] br[205] br[204] br[203] br[202] br[201] br[200] br[199] br[198] br[197] br[196] br[195] br[194] br[193] br[192] br[191] br[190] br[189] br[188] br[187] br[186] br[185] br[184] br[183] br[182] br[181] br[180] br[179] br[178] br[177] br[176] br[175] br[174] br[173] br[172] br[171] br[170] br[169] br[168] br[167] br[166] br[165] br[164] br[163] br[162] br[161] br[160] br[159] br[158] br[157] br[156] br[155] br[154] br[153] br[152] br[151] br[150] br[149] br[148] br[147] br[146] br[145] br[144] br[143] br[142] br[141] br[140] br[139] br[138] br[137] br[136] br[135] br[134] br[133] br[132] br[131] br[130] br[129] br[128] br[127] br[126] br[125] br[124] br[123] br[122] br[121] br[120] br[119] br[118] br[117] br[116] br[115] br[114] br[113] br[112] br[111] br[110] br[109] br[108] br[107] br[106] br[105] br[104] br[103] br[102] br[101] br[100] br[99] br[98] br[97] br[96] br[95] br[94] br[93] br[92] br[91] br[90] br[89] br[88] br[87] br[86] br[85] br[84] br[83] br[82] br[81] br[80] br[79] br[78] br[77] br[76] br[75] br[74] br[73] br[72] br[71] br[70] br[69] br[68] br[67] br[66] br[65] br[64] br[63] br[62] br[61] br[60] br[59] br[58] br[57] br[56] br[55] br[54] br[53] br[52] br[51] br[50] br[49] br[48] br[47] br[46] br[45] br[44] br[43] br[42] br[41] br[40] br[39] br[38] br[37] br[36] br[35] br[34] br[33] br[32] br[31] br[30] br[29] br[28] br[27] br[26] br[25] br[24] br[23] br[22] br[21] br[20] br[19] br[18] br[17] br[16] br[15] br[14] br[13] br[12] br[11] br[10] br[9] br[8] br[7] br[6] br[5] br[4] br[3] br[2] br[1] br[0] bl_read[31] bl_read[30] bl_read[29] bl_read[28] bl_read[27] bl_read[26] bl_read[25] bl_read[24] bl_read[23] bl_read[22] bl_read[21] bl_read[20] bl_read[19] bl_read[18] bl_read[17] bl_read[16] bl_read[15] bl_read[14] bl_read[13] bl_read[12] bl_read[11] bl_read[10] bl_read[9] bl_read[8] bl_read[7] bl_read[6] bl_read[5] bl_read[4] bl_read[3] bl_read[2] bl_read[1] bl_read[0] br_read[31] br_read[30] br_read[29] br_read[28] br_read[27] br_read[26] br_read[25] br_read[24] br_read[23] br_read[22] br_read[21] br_read[20] br_read[19] br_read[18] br_read[17] br_read[16] br_read[15] br_read[14] br_read[13] br_read[12] br_read[11] br_read[10] br_read[9] br_read[8] br_read[7] br_read[6] br_read[5] br_read[4] br_read[3] br_read[2] br_read[1] br_read[0] vdd 
+ read_mux_array 
* No parameters

xcol_inv_array 
+ bank_din[31] bank_din[30] bank_din[29] bank_din[28] bank_din[27] bank_din[26] bank_din[25] bank_din[24] bank_din[23] bank_din[22] bank_din[21] bank_din[20] bank_din[19] bank_din[18] bank_din[17] bank_din[16] bank_din[15] bank_din[14] bank_din[13] bank_din[12] bank_din[11] bank_din[10] bank_din[9] bank_din[8] bank_din[7] bank_din[6] bank_din[5] bank_din[4] bank_din[3] bank_din[2] bank_din[1] bank_din[0] bank_din_b[31] bank_din_b[30] bank_din_b[29] bank_din_b[28] bank_din_b[27] bank_din_b[26] bank_din_b[25] bank_din_b[24] bank_din_b[23] bank_din_b[22] bank_din_b[21] bank_din_b[20] bank_din_b[19] bank_din_b[18] bank_din_b[17] bank_din_b[16] bank_din_b[15] bank_din_b[14] bank_din_b[13] bank_din_b[12] bank_din_b[11] bank_din_b[10] bank_din_b[9] bank_din_b[8] bank_din_b[7] bank_din_b[6] bank_din_b[5] bank_din_b[4] bank_din_b[3] bank_din_b[2] bank_din_b[1] bank_din_b[0] vdd vss 
+ col_inv_array 
* No parameters

xsense_amp_array 
+ vdd vss sense_amp_en bl_read[31] bl_read[30] bl_read[29] bl_read[28] bl_read[27] bl_read[26] bl_read[25] bl_read[24] bl_read[23] bl_read[22] bl_read[21] bl_read[20] bl_read[19] bl_read[18] bl_read[17] bl_read[16] bl_read[15] bl_read[14] bl_read[13] bl_read[12] bl_read[11] bl_read[10] bl_read[9] bl_read[8] bl_read[7] bl_read[6] bl_read[5] bl_read[4] bl_read[3] bl_read[2] bl_read[1] bl_read[0] br_read[31] br_read[30] br_read[29] br_read[28] br_read[27] br_read[26] br_read[25] br_read[24] br_read[23] br_read[22] br_read[21] br_read[20] br_read[19] br_read[18] br_read[17] br_read[16] br_read[15] br_read[14] br_read[13] br_read[12] br_read[11] br_read[10] br_read[9] br_read[8] br_read[7] br_read[6] br_read[5] br_read[4] br_read[3] br_read[2] br_read[1] br_read[0] sa_outp[31] sa_outp[30] sa_outp[29] sa_outp[28] sa_outp[27] sa_outp[26] sa_outp[25] sa_outp[24] sa_outp[23] sa_outp[22] sa_outp[21] sa_outp[20] sa_outp[19] sa_outp[18] sa_outp[17] sa_outp[16] sa_outp[15] sa_outp[14] sa_outp[13] sa_outp[12] sa_outp[11] sa_outp[10] sa_outp[9] sa_outp[8] sa_outp[7] sa_outp[6] sa_outp[5] sa_outp[4] sa_outp[3] sa_outp[2] sa_outp[1] sa_outp[0] sa_outn[31] sa_outn[30] sa_outn[29] sa_outn[28] sa_outn[27] sa_outn[26] sa_outn[25] sa_outn[24] sa_outn[23] sa_outn[22] sa_outn[21] sa_outn[20] sa_outn[19] sa_outn[18] sa_outn[17] sa_outn[16] sa_outn[15] sa_outn[14] sa_outn[13] sa_outn[12] sa_outn[11] sa_outn[10] sa_outn[9] sa_outn[8] sa_outn[7] sa_outn[6] sa_outn[5] sa_outn[4] sa_outn[3] sa_outn[2] sa_outn[1] sa_outn[0] 
+ sense_amp_array 
* No parameters

xdout_buf_array 
+ sa_outp[31] sa_outp[30] sa_outp[29] sa_outp[28] sa_outp[27] sa_outp[26] sa_outp[25] sa_outp[24] sa_outp[23] sa_outp[22] sa_outp[21] sa_outp[20] sa_outp[19] sa_outp[18] sa_outp[17] sa_outp[16] sa_outp[15] sa_outp[14] sa_outp[13] sa_outp[12] sa_outp[11] sa_outp[10] sa_outp[9] sa_outp[8] sa_outp[7] sa_outp[6] sa_outp[5] sa_outp[4] sa_outp[3] sa_outp[2] sa_outp[1] sa_outp[0] sa_outn[31] sa_outn[30] sa_outn[29] sa_outn[28] sa_outn[27] sa_outn[26] sa_outn[25] sa_outn[24] sa_outn[23] sa_outn[22] sa_outn[21] sa_outn[20] sa_outn[19] sa_outn[18] sa_outn[17] sa_outn[16] sa_outn[15] sa_outn[14] sa_outn[13] sa_outn[12] sa_outn[11] sa_outn[10] sa_outn[9] sa_outn[8] sa_outn[7] sa_outn[6] sa_outn[5] sa_outn[4] sa_outn[3] sa_outn[2] sa_outn[1] sa_outn[0] dout[31] dout[30] dout[29] dout[28] dout[27] dout[26] dout[25] dout[24] dout[23] dout[22] dout[21] dout[20] dout[19] dout[18] dout[17] dout[16] dout[15] dout[14] dout[13] dout[12] dout[11] dout[10] dout[9] dout[8] dout[7] dout[6] dout[5] dout[4] dout[3] dout[2] dout[1] dout[0] dout_b[31] dout_b[30] dout_b[29] dout_b[28] dout_b[27] dout_b[26] dout_b[25] dout_b[24] dout_b[23] dout_b[22] dout_b[21] dout_b[20] dout_b[19] dout_b[18] dout_b[17] dout_b[16] dout_b[15] dout_b[14] dout_b[13] dout_b[12] dout_b[11] dout_b[10] dout_b[9] dout_b[8] dout_b[7] dout_b[6] dout_b[5] dout_b[4] dout_b[3] dout_b[2] dout_b[1] dout_b[0] vdd vss 
+ dout_buf_array 
* No parameters

xcontrol_logic 
+ clk bank_we rbl pc_b wl_en wr_en sense_amp_en vdd vss 
+ sramgen_control_replica_v1 
* No parameters

xcolumn_decoder 
+ vdd vss bank_addr[2] bank_addr[1] bank_addr[0] bank_addr_b[2] bank_addr_b[1] bank_addr_b[0] col_sel[7] col_sel[6] col_sel[5] col_sel[4] col_sel[3] col_sel[2] col_sel[1] col_sel[0] col_sel_b[7] col_sel_b[6] col_sel_b[5] col_sel_b[4] col_sel_b[3] col_sel_b[2] col_sel_b[1] col_sel_b[0] 
+ column_decoder 
* No parameters

xwe_control 
+ wr_en col_sel[7] col_sel[6] col_sel[5] col_sel[4] col_sel[3] col_sel[2] col_sel[1] col_sel[0] write_driver_en[7] write_driver_en[6] write_driver_en[5] write_driver_en[4] write_driver_en[3] write_driver_en[2] write_driver_en[1] write_driver_en[0] vdd vss 
+ we_control 
* No parameters

.ENDS

