VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sram22_512x64m4w8
  CLASS BLOCK ;
  ORIGIN 80.225 183.565 ;
  FOREIGN sram22_512x64m4w8 -80.225 -183.565 ;
  SIZE 488.21 BY 429.01 ;
  SYMMETRY X Y R90 ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 398.995 244.04 399.325 245.17 ;
        RECT 398.995 239.875 399.325 240.205 ;
        RECT 398.995 238.515 399.325 238.845 ;
        RECT 398.995 237.155 399.325 237.485 ;
        RECT 398.995 235.17 399.325 235.5 ;
        RECT 398.995 232.995 399.325 233.325 ;
        RECT 398.995 231.415 399.325 231.745 ;
        RECT 398.995 230.565 399.325 230.895 ;
        RECT 398.995 228.255 399.325 228.585 ;
        RECT 398.995 227.405 399.325 227.735 ;
        RECT 398.995 225.095 399.325 225.425 ;
        RECT 398.995 224.245 399.325 224.575 ;
        RECT 398.995 221.935 399.325 222.265 ;
        RECT 398.995 221.085 399.325 221.415 ;
        RECT 398.995 218.775 399.325 219.105 ;
        RECT 398.995 217.195 399.325 217.525 ;
        RECT 398.995 216.345 399.325 216.675 ;
        RECT 398.995 214.035 399.325 214.365 ;
        RECT 398.995 213.185 399.325 213.515 ;
        RECT 398.995 210.875 399.325 211.205 ;
        RECT 398.995 210.025 399.325 210.355 ;
        RECT 398.995 207.715 399.325 208.045 ;
        RECT 398.995 206.865 399.325 207.195 ;
        RECT 398.995 204.555 399.325 204.885 ;
        RECT 398.995 202.975 399.325 203.305 ;
        RECT 398.995 202.125 399.325 202.455 ;
        RECT 398.995 199.815 399.325 200.145 ;
        RECT 398.995 198.965 399.325 199.295 ;
        RECT 398.995 196.655 399.325 196.985 ;
        RECT 398.995 195.805 399.325 196.135 ;
        RECT 398.995 193.495 399.325 193.825 ;
        RECT 398.995 192.645 399.325 192.975 ;
        RECT 398.995 190.335 399.325 190.665 ;
        RECT 398.995 188.755 399.325 189.085 ;
        RECT 398.995 187.905 399.325 188.235 ;
        RECT 398.995 185.595 399.325 185.925 ;
        RECT 398.995 184.745 399.325 185.075 ;
        RECT 398.995 182.435 399.325 182.765 ;
        RECT 398.995 181.585 399.325 181.915 ;
        RECT 398.995 179.275 399.325 179.605 ;
        RECT 398.995 178.425 399.325 178.755 ;
        RECT 398.995 176.115 399.325 176.445 ;
        RECT 398.995 174.535 399.325 174.865 ;
        RECT 398.995 173.685 399.325 174.015 ;
        RECT 398.995 171.375 399.325 171.705 ;
        RECT 398.995 170.525 399.325 170.855 ;
        RECT 398.995 168.215 399.325 168.545 ;
        RECT 398.995 167.365 399.325 167.695 ;
        RECT 398.995 165.055 399.325 165.385 ;
        RECT 398.995 164.205 399.325 164.535 ;
        RECT 398.995 161.895 399.325 162.225 ;
        RECT 398.995 160.315 399.325 160.645 ;
        RECT 398.995 159.465 399.325 159.795 ;
        RECT 398.995 157.155 399.325 157.485 ;
        RECT 398.995 156.305 399.325 156.635 ;
        RECT 398.995 153.995 399.325 154.325 ;
        RECT 398.995 153.145 399.325 153.475 ;
        RECT 398.995 150.835 399.325 151.165 ;
        RECT 398.995 149.985 399.325 150.315 ;
        RECT 398.995 147.675 399.325 148.005 ;
        RECT 398.995 146.095 399.325 146.425 ;
        RECT 398.995 145.245 399.325 145.575 ;
        RECT 398.995 142.935 399.325 143.265 ;
        RECT 398.995 142.085 399.325 142.415 ;
        RECT 398.995 139.775 399.325 140.105 ;
        RECT 398.995 138.925 399.325 139.255 ;
        RECT 398.995 136.615 399.325 136.945 ;
        RECT 398.995 135.765 399.325 136.095 ;
        RECT 398.995 133.455 399.325 133.785 ;
        RECT 398.995 131.875 399.325 132.205 ;
        RECT 398.995 131.025 399.325 131.355 ;
        RECT 398.995 128.715 399.325 129.045 ;
        RECT 398.995 127.865 399.325 128.195 ;
        RECT 398.995 125.555 399.325 125.885 ;
        RECT 398.995 124.705 399.325 125.035 ;
        RECT 398.995 122.395 399.325 122.725 ;
        RECT 398.995 121.545 399.325 121.875 ;
        RECT 398.995 119.235 399.325 119.565 ;
        RECT 398.995 117.655 399.325 117.985 ;
        RECT 398.995 116.805 399.325 117.135 ;
        RECT 398.995 114.495 399.325 114.825 ;
        RECT 398.995 113.645 399.325 113.975 ;
        RECT 398.995 111.335 399.325 111.665 ;
        RECT 398.995 110.485 399.325 110.815 ;
        RECT 398.995 108.175 399.325 108.505 ;
        RECT 398.995 107.325 399.325 107.655 ;
        RECT 398.995 105.015 399.325 105.345 ;
        RECT 398.995 103.435 399.325 103.765 ;
        RECT 398.995 102.585 399.325 102.915 ;
        RECT 398.995 100.275 399.325 100.605 ;
        RECT 398.995 99.425 399.325 99.755 ;
        RECT 398.995 97.115 399.325 97.445 ;
        RECT 398.995 96.265 399.325 96.595 ;
        RECT 398.995 93.955 399.325 94.285 ;
        RECT 398.995 93.105 399.325 93.435 ;
        RECT 398.995 90.795 399.325 91.125 ;
        RECT 398.995 89.215 399.325 89.545 ;
        RECT 398.995 88.365 399.325 88.695 ;
        RECT 398.995 86.055 399.325 86.385 ;
        RECT 398.995 85.205 399.325 85.535 ;
        RECT 398.995 82.895 399.325 83.225 ;
        RECT 398.995 82.045 399.325 82.375 ;
        RECT 398.995 79.735 399.325 80.065 ;
        RECT 398.995 78.885 399.325 79.215 ;
        RECT 398.995 76.575 399.325 76.905 ;
        RECT 398.995 74.995 399.325 75.325 ;
        RECT 398.995 74.145 399.325 74.475 ;
        RECT 398.995 71.835 399.325 72.165 ;
        RECT 398.995 70.985 399.325 71.315 ;
        RECT 398.995 68.675 399.325 69.005 ;
        RECT 398.995 67.825 399.325 68.155 ;
        RECT 398.995 65.515 399.325 65.845 ;
        RECT 398.995 64.665 399.325 64.995 ;
        RECT 398.995 62.355 399.325 62.685 ;
        RECT 398.995 60.775 399.325 61.105 ;
        RECT 398.995 59.925 399.325 60.255 ;
        RECT 398.995 57.615 399.325 57.945 ;
        RECT 398.995 56.765 399.325 57.095 ;
        RECT 398.995 54.455 399.325 54.785 ;
        RECT 398.995 53.605 399.325 53.935 ;
        RECT 398.995 51.295 399.325 51.625 ;
        RECT 398.995 50.445 399.325 50.775 ;
        RECT 398.995 48.135 399.325 48.465 ;
        RECT 398.995 46.555 399.325 46.885 ;
        RECT 398.995 45.705 399.325 46.035 ;
        RECT 398.995 43.395 399.325 43.725 ;
        RECT 398.995 42.545 399.325 42.875 ;
        RECT 398.995 40.235 399.325 40.565 ;
        RECT 398.995 39.385 399.325 39.715 ;
        RECT 398.995 37.075 399.325 37.405 ;
        RECT 398.995 36.225 399.325 36.555 ;
        RECT 398.995 33.915 399.325 34.245 ;
        RECT 398.995 32.335 399.325 32.665 ;
        RECT 398.995 31.485 399.325 31.815 ;
        RECT 398.995 29.175 399.325 29.505 ;
        RECT 398.995 28.325 399.325 28.655 ;
        RECT 398.995 26.015 399.325 26.345 ;
        RECT 398.995 25.165 399.325 25.495 ;
        RECT 398.995 22.855 399.325 23.185 ;
        RECT 398.995 22.005 399.325 22.335 ;
        RECT 398.995 19.695 399.325 20.025 ;
        RECT 398.995 18.115 399.325 18.445 ;
        RECT 398.995 17.265 399.325 17.595 ;
        RECT 398.995 14.955 399.325 15.285 ;
        RECT 398.995 14.105 399.325 14.435 ;
        RECT 398.995 11.795 399.325 12.125 ;
        RECT 398.995 10.945 399.325 11.275 ;
        RECT 398.995 8.635 399.325 8.965 ;
        RECT 398.995 7.785 399.325 8.115 ;
        RECT 398.995 5.475 399.325 5.805 ;
        RECT 398.995 3.895 399.325 4.225 ;
        RECT 398.995 3.045 399.325 3.375 ;
        RECT 398.995 0.87 399.325 1.2 ;
        RECT 398.995 -0.845 399.325 -0.515 ;
        RECT 398.995 -2.205 399.325 -1.875 ;
        RECT 398.995 -3.565 399.325 -3.235 ;
        RECT 398.995 -4.925 399.325 -4.595 ;
        RECT 398.995 -6.285 399.325 -5.955 ;
        RECT 398.995 -7.645 399.325 -7.315 ;
        RECT 398.995 -9.005 399.325 -8.675 ;
        RECT 398.995 -10.365 399.325 -10.035 ;
        RECT 398.995 -11.725 399.325 -11.395 ;
        RECT 398.995 -13.085 399.325 -12.755 ;
        RECT 398.995 -14.445 399.325 -14.115 ;
        RECT 398.995 -15.805 399.325 -15.475 ;
        RECT 398.995 -17.165 399.325 -16.835 ;
        RECT 398.995 -18.525 399.325 -18.195 ;
        RECT 398.995 -19.885 399.325 -19.555 ;
        RECT 398.995 -21.245 399.325 -20.915 ;
        RECT 398.995 -22.605 399.325 -22.275 ;
        RECT 398.995 -23.965 399.325 -23.635 ;
        RECT 398.995 -25.325 399.325 -24.995 ;
        RECT 398.995 -26.685 399.325 -26.355 ;
        RECT 398.995 -28.045 399.325 -27.715 ;
        RECT 398.995 -29.405 399.325 -29.075 ;
        RECT 398.995 -30.765 399.325 -30.435 ;
        RECT 398.995 -32.125 399.325 -31.795 ;
        RECT 398.995 -33.485 399.325 -33.155 ;
        RECT 398.995 -34.845 399.325 -34.515 ;
        RECT 398.995 -36.205 399.325 -35.875 ;
        RECT 398.995 -37.565 399.325 -37.235 ;
        RECT 398.995 -38.925 399.325 -38.595 ;
        RECT 398.995 -40.285 399.325 -39.955 ;
        RECT 398.995 -41.645 399.325 -41.315 ;
        RECT 398.995 -43.005 399.325 -42.675 ;
        RECT 398.995 -44.365 399.325 -44.035 ;
        RECT 398.995 -45.725 399.325 -45.395 ;
        RECT 398.995 -47.085 399.325 -46.755 ;
        RECT 398.995 -48.445 399.325 -48.115 ;
        RECT 398.995 -49.805 399.325 -49.475 ;
        RECT 398.995 -51.165 399.325 -50.835 ;
        RECT 398.995 -52.525 399.325 -52.195 ;
        RECT 398.995 -53.885 399.325 -53.555 ;
        RECT 398.995 -55.245 399.325 -54.915 ;
        RECT 398.995 -56.605 399.325 -56.275 ;
        RECT 398.995 -57.965 399.325 -57.635 ;
        RECT 398.995 -59.325 399.325 -58.995 ;
        RECT 398.995 -60.685 399.325 -60.355 ;
        RECT 398.995 -62.045 399.325 -61.715 ;
        RECT 398.995 -63.405 399.325 -63.075 ;
        RECT 398.995 -64.765 399.325 -64.435 ;
        RECT 398.995 -66.125 399.325 -65.795 ;
        RECT 398.995 -67.485 399.325 -67.155 ;
        RECT 398.995 -68.845 399.325 -68.515 ;
        RECT 398.995 -70.205 399.325 -69.875 ;
        RECT 398.995 -71.565 399.325 -71.235 ;
        RECT 398.995 -72.925 399.325 -72.595 ;
        RECT 398.995 -74.285 399.325 -73.955 ;
        RECT 398.995 -75.645 399.325 -75.315 ;
        RECT 398.995 -77.005 399.325 -76.675 ;
        RECT 398.995 -78.365 399.325 -78.035 ;
        RECT 398.995 -79.725 399.325 -79.395 ;
        RECT 398.995 -81.085 399.325 -80.755 ;
        RECT 398.995 -82.445 399.325 -82.115 ;
        RECT 398.995 -83.805 399.325 -83.475 ;
        RECT 398.995 -85.165 399.325 -84.835 ;
        RECT 398.995 -86.525 399.325 -86.195 ;
        RECT 398.995 -87.885 399.325 -87.555 ;
        RECT 398.995 -89.245 399.325 -88.915 ;
        RECT 398.995 -90.605 399.325 -90.275 ;
        RECT 398.995 -91.965 399.325 -91.635 ;
        RECT 398.995 -93.325 399.325 -92.995 ;
        RECT 398.995 -94.685 399.325 -94.355 ;
        RECT 398.995 -96.045 399.325 -95.715 ;
        RECT 398.995 -97.405 399.325 -97.075 ;
        RECT 398.995 -98.765 399.325 -98.435 ;
        RECT 398.995 -100.125 399.325 -99.795 ;
        RECT 398.995 -101.485 399.325 -101.155 ;
        RECT 398.995 -102.845 399.325 -102.515 ;
        RECT 398.995 -104.205 399.325 -103.875 ;
        RECT 398.995 -105.565 399.325 -105.235 ;
        RECT 398.995 -106.925 399.325 -106.595 ;
        RECT 398.995 -108.285 399.325 -107.955 ;
        RECT 398.995 -109.645 399.325 -109.315 ;
        RECT 398.995 -111.005 399.325 -110.675 ;
        RECT 398.995 -112.365 399.325 -112.035 ;
        RECT 398.995 -113.725 399.325 -113.395 ;
        RECT 398.995 -115.085 399.325 -114.755 ;
        RECT 398.995 -116.445 399.325 -116.115 ;
        RECT 398.995 -117.805 399.325 -117.475 ;
        RECT 398.995 -119.165 399.325 -118.835 ;
        RECT 398.995 -120.525 399.325 -120.195 ;
        RECT 398.995 -121.885 399.325 -121.555 ;
        RECT 398.995 -123.245 399.325 -122.915 ;
        RECT 398.995 -124.605 399.325 -124.275 ;
        RECT 398.995 -125.965 399.325 -125.635 ;
        RECT 398.995 -127.325 399.325 -126.995 ;
        RECT 398.995 -128.685 399.325 -128.355 ;
        RECT 398.995 -130.045 399.325 -129.715 ;
        RECT 398.995 -131.405 399.325 -131.075 ;
        RECT 398.995 -132.765 399.325 -132.435 ;
        RECT 398.995 -134.125 399.325 -133.795 ;
        RECT 398.995 -135.485 399.325 -135.155 ;
        RECT 398.995 -136.845 399.325 -136.515 ;
        RECT 398.995 -138.205 399.325 -137.875 ;
        RECT 398.995 -139.565 399.325 -139.235 ;
        RECT 398.995 -140.925 399.325 -140.595 ;
        RECT 398.995 -142.285 399.325 -141.955 ;
        RECT 398.995 -143.645 399.325 -143.315 ;
        RECT 398.995 -145.005 399.325 -144.675 ;
        RECT 398.995 -146.365 399.325 -146.035 ;
        RECT 398.995 -147.725 399.325 -147.395 ;
        RECT 398.995 -149.085 399.325 -148.755 ;
        RECT 398.995 -150.445 399.325 -150.115 ;
        RECT 398.995 -151.805 399.325 -151.475 ;
        RECT 398.995 -153.165 399.325 -152.835 ;
        RECT 398.995 -154.525 399.325 -154.195 ;
        RECT 398.995 -155.885 399.325 -155.555 ;
        RECT 398.995 -157.245 399.325 -156.915 ;
        RECT 398.995 -158.605 399.325 -158.275 ;
        RECT 398.995 -159.965 399.325 -159.635 ;
        RECT 398.995 -161.325 399.325 -160.995 ;
        RECT 398.995 -162.685 399.325 -162.355 ;
        RECT 398.995 -164.045 399.325 -163.715 ;
        RECT 398.995 -165.405 399.325 -165.075 ;
        RECT 398.995 -166.765 399.325 -166.435 ;
        RECT 398.995 -168.125 399.325 -167.795 ;
        RECT 398.995 -169.485 399.325 -169.155 ;
        RECT 398.995 -170.845 399.325 -170.515 ;
        RECT 398.995 -172.205 399.325 -171.875 ;
        RECT 398.995 -173.565 399.325 -173.235 ;
        RECT 398.995 -174.925 399.325 -174.595 ;
        RECT 398.995 -176.285 399.325 -175.955 ;
        RECT 398.995 -177.645 399.325 -177.315 ;
        RECT 398.995 -183.29 399.325 -182.16 ;
        RECT 399 -183.405 399.32 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 400.355 244.04 400.685 245.17 ;
        RECT 400.355 239.875 400.685 240.205 ;
        RECT 400.355 238.515 400.685 238.845 ;
        RECT 400.355 237.155 400.685 237.485 ;
        RECT 400.355 235.17 400.685 235.5 ;
        RECT 400.355 232.995 400.685 233.325 ;
        RECT 400.355 231.415 400.685 231.745 ;
        RECT 400.355 230.565 400.685 230.895 ;
        RECT 400.355 228.255 400.685 228.585 ;
        RECT 400.355 227.405 400.685 227.735 ;
        RECT 400.355 225.095 400.685 225.425 ;
        RECT 400.355 224.245 400.685 224.575 ;
        RECT 400.355 221.935 400.685 222.265 ;
        RECT 400.355 221.085 400.685 221.415 ;
        RECT 400.355 218.775 400.685 219.105 ;
        RECT 400.355 217.195 400.685 217.525 ;
        RECT 400.355 216.345 400.685 216.675 ;
        RECT 400.355 214.035 400.685 214.365 ;
        RECT 400.355 213.185 400.685 213.515 ;
        RECT 400.355 210.875 400.685 211.205 ;
        RECT 400.355 210.025 400.685 210.355 ;
        RECT 400.355 207.715 400.685 208.045 ;
        RECT 400.355 206.865 400.685 207.195 ;
        RECT 400.355 204.555 400.685 204.885 ;
        RECT 400.355 202.975 400.685 203.305 ;
        RECT 400.355 202.125 400.685 202.455 ;
        RECT 400.355 199.815 400.685 200.145 ;
        RECT 400.355 198.965 400.685 199.295 ;
        RECT 400.355 196.655 400.685 196.985 ;
        RECT 400.355 195.805 400.685 196.135 ;
        RECT 400.355 193.495 400.685 193.825 ;
        RECT 400.355 192.645 400.685 192.975 ;
        RECT 400.355 190.335 400.685 190.665 ;
        RECT 400.355 188.755 400.685 189.085 ;
        RECT 400.355 187.905 400.685 188.235 ;
        RECT 400.355 185.595 400.685 185.925 ;
        RECT 400.355 184.745 400.685 185.075 ;
        RECT 400.355 182.435 400.685 182.765 ;
        RECT 400.355 181.585 400.685 181.915 ;
        RECT 400.355 179.275 400.685 179.605 ;
        RECT 400.355 178.425 400.685 178.755 ;
        RECT 400.355 176.115 400.685 176.445 ;
        RECT 400.355 174.535 400.685 174.865 ;
        RECT 400.355 173.685 400.685 174.015 ;
        RECT 400.355 171.375 400.685 171.705 ;
        RECT 400.355 170.525 400.685 170.855 ;
        RECT 400.355 168.215 400.685 168.545 ;
        RECT 400.355 167.365 400.685 167.695 ;
        RECT 400.355 165.055 400.685 165.385 ;
        RECT 400.355 164.205 400.685 164.535 ;
        RECT 400.355 161.895 400.685 162.225 ;
        RECT 400.355 160.315 400.685 160.645 ;
        RECT 400.355 159.465 400.685 159.795 ;
        RECT 400.355 157.155 400.685 157.485 ;
        RECT 400.355 156.305 400.685 156.635 ;
        RECT 400.355 153.995 400.685 154.325 ;
        RECT 400.355 153.145 400.685 153.475 ;
        RECT 400.355 150.835 400.685 151.165 ;
        RECT 400.355 149.985 400.685 150.315 ;
        RECT 400.355 147.675 400.685 148.005 ;
        RECT 400.355 146.095 400.685 146.425 ;
        RECT 400.355 145.245 400.685 145.575 ;
        RECT 400.355 142.935 400.685 143.265 ;
        RECT 400.355 142.085 400.685 142.415 ;
        RECT 400.355 139.775 400.685 140.105 ;
        RECT 400.355 138.925 400.685 139.255 ;
        RECT 400.355 136.615 400.685 136.945 ;
        RECT 400.355 135.765 400.685 136.095 ;
        RECT 400.355 133.455 400.685 133.785 ;
        RECT 400.355 131.875 400.685 132.205 ;
        RECT 400.355 131.025 400.685 131.355 ;
        RECT 400.355 128.715 400.685 129.045 ;
        RECT 400.355 127.865 400.685 128.195 ;
        RECT 400.355 125.555 400.685 125.885 ;
        RECT 400.355 124.705 400.685 125.035 ;
        RECT 400.355 122.395 400.685 122.725 ;
        RECT 400.355 121.545 400.685 121.875 ;
        RECT 400.355 119.235 400.685 119.565 ;
        RECT 400.355 117.655 400.685 117.985 ;
        RECT 400.355 116.805 400.685 117.135 ;
        RECT 400.355 114.495 400.685 114.825 ;
        RECT 400.355 113.645 400.685 113.975 ;
        RECT 400.355 111.335 400.685 111.665 ;
        RECT 400.355 110.485 400.685 110.815 ;
        RECT 400.355 108.175 400.685 108.505 ;
        RECT 400.355 107.325 400.685 107.655 ;
        RECT 400.355 105.015 400.685 105.345 ;
        RECT 400.355 103.435 400.685 103.765 ;
        RECT 400.355 102.585 400.685 102.915 ;
        RECT 400.355 100.275 400.685 100.605 ;
        RECT 400.355 99.425 400.685 99.755 ;
        RECT 400.355 97.115 400.685 97.445 ;
        RECT 400.355 96.265 400.685 96.595 ;
        RECT 400.355 93.955 400.685 94.285 ;
        RECT 400.355 93.105 400.685 93.435 ;
        RECT 400.355 90.795 400.685 91.125 ;
        RECT 400.355 89.215 400.685 89.545 ;
        RECT 400.355 88.365 400.685 88.695 ;
        RECT 400.355 86.055 400.685 86.385 ;
        RECT 400.355 85.205 400.685 85.535 ;
        RECT 400.355 82.895 400.685 83.225 ;
        RECT 400.355 82.045 400.685 82.375 ;
        RECT 400.355 79.735 400.685 80.065 ;
        RECT 400.355 78.885 400.685 79.215 ;
        RECT 400.355 76.575 400.685 76.905 ;
        RECT 400.355 74.995 400.685 75.325 ;
        RECT 400.355 74.145 400.685 74.475 ;
        RECT 400.355 71.835 400.685 72.165 ;
        RECT 400.355 70.985 400.685 71.315 ;
        RECT 400.355 68.675 400.685 69.005 ;
        RECT 400.355 67.825 400.685 68.155 ;
        RECT 400.355 65.515 400.685 65.845 ;
        RECT 400.355 64.665 400.685 64.995 ;
        RECT 400.355 62.355 400.685 62.685 ;
        RECT 400.355 60.775 400.685 61.105 ;
        RECT 400.355 59.925 400.685 60.255 ;
        RECT 400.355 57.615 400.685 57.945 ;
        RECT 400.355 56.765 400.685 57.095 ;
        RECT 400.355 54.455 400.685 54.785 ;
        RECT 400.355 53.605 400.685 53.935 ;
        RECT 400.355 51.295 400.685 51.625 ;
        RECT 400.355 50.445 400.685 50.775 ;
        RECT 400.355 48.135 400.685 48.465 ;
        RECT 400.355 46.555 400.685 46.885 ;
        RECT 400.355 45.705 400.685 46.035 ;
        RECT 400.355 43.395 400.685 43.725 ;
        RECT 400.355 42.545 400.685 42.875 ;
        RECT 400.355 40.235 400.685 40.565 ;
        RECT 400.355 39.385 400.685 39.715 ;
        RECT 400.355 37.075 400.685 37.405 ;
        RECT 400.355 36.225 400.685 36.555 ;
        RECT 400.355 33.915 400.685 34.245 ;
        RECT 400.355 32.335 400.685 32.665 ;
        RECT 400.355 31.485 400.685 31.815 ;
        RECT 400.355 29.175 400.685 29.505 ;
        RECT 400.355 28.325 400.685 28.655 ;
        RECT 400.355 26.015 400.685 26.345 ;
        RECT 400.355 25.165 400.685 25.495 ;
        RECT 400.355 22.855 400.685 23.185 ;
        RECT 400.355 22.005 400.685 22.335 ;
        RECT 400.355 19.695 400.685 20.025 ;
        RECT 400.355 18.115 400.685 18.445 ;
        RECT 400.355 17.265 400.685 17.595 ;
        RECT 400.355 14.955 400.685 15.285 ;
        RECT 400.355 14.105 400.685 14.435 ;
        RECT 400.355 11.795 400.685 12.125 ;
        RECT 400.355 10.945 400.685 11.275 ;
        RECT 400.355 8.635 400.685 8.965 ;
        RECT 400.355 7.785 400.685 8.115 ;
        RECT 400.355 5.475 400.685 5.805 ;
        RECT 400.355 3.895 400.685 4.225 ;
        RECT 400.355 3.045 400.685 3.375 ;
        RECT 400.355 0.87 400.685 1.2 ;
        RECT 400.355 -0.845 400.685 -0.515 ;
        RECT 400.355 -2.205 400.685 -1.875 ;
        RECT 400.355 -3.565 400.685 -3.235 ;
        RECT 400.355 -4.925 400.685 -4.595 ;
        RECT 400.355 -6.285 400.685 -5.955 ;
        RECT 400.355 -7.645 400.685 -7.315 ;
        RECT 400.355 -9.005 400.685 -8.675 ;
        RECT 400.355 -10.365 400.685 -10.035 ;
        RECT 400.355 -11.725 400.685 -11.395 ;
        RECT 400.355 -13.085 400.685 -12.755 ;
        RECT 400.355 -14.445 400.685 -14.115 ;
        RECT 400.355 -15.805 400.685 -15.475 ;
        RECT 400.355 -17.165 400.685 -16.835 ;
        RECT 400.355 -18.525 400.685 -18.195 ;
        RECT 400.355 -19.885 400.685 -19.555 ;
        RECT 400.355 -21.245 400.685 -20.915 ;
        RECT 400.355 -22.605 400.685 -22.275 ;
        RECT 400.355 -23.965 400.685 -23.635 ;
        RECT 400.355 -25.325 400.685 -24.995 ;
        RECT 400.355 -26.685 400.685 -26.355 ;
        RECT 400.355 -28.045 400.685 -27.715 ;
        RECT 400.355 -29.405 400.685 -29.075 ;
        RECT 400.355 -30.765 400.685 -30.435 ;
        RECT 400.355 -32.125 400.685 -31.795 ;
        RECT 400.355 -33.485 400.685 -33.155 ;
        RECT 400.355 -34.845 400.685 -34.515 ;
        RECT 400.355 -36.205 400.685 -35.875 ;
        RECT 400.355 -37.565 400.685 -37.235 ;
        RECT 400.355 -38.925 400.685 -38.595 ;
        RECT 400.355 -40.285 400.685 -39.955 ;
        RECT 400.355 -41.645 400.685 -41.315 ;
        RECT 400.355 -43.005 400.685 -42.675 ;
        RECT 400.355 -44.365 400.685 -44.035 ;
        RECT 400.355 -45.725 400.685 -45.395 ;
        RECT 400.355 -47.085 400.685 -46.755 ;
        RECT 400.355 -48.445 400.685 -48.115 ;
        RECT 400.355 -49.805 400.685 -49.475 ;
        RECT 400.355 -51.165 400.685 -50.835 ;
        RECT 400.355 -52.525 400.685 -52.195 ;
        RECT 400.355 -53.885 400.685 -53.555 ;
        RECT 400.355 -55.245 400.685 -54.915 ;
        RECT 400.355 -56.605 400.685 -56.275 ;
        RECT 400.355 -57.965 400.685 -57.635 ;
        RECT 400.355 -59.325 400.685 -58.995 ;
        RECT 400.355 -60.685 400.685 -60.355 ;
        RECT 400.355 -62.045 400.685 -61.715 ;
        RECT 400.355 -63.405 400.685 -63.075 ;
        RECT 400.355 -64.765 400.685 -64.435 ;
        RECT 400.355 -66.125 400.685 -65.795 ;
        RECT 400.355 -67.485 400.685 -67.155 ;
        RECT 400.355 -68.845 400.685 -68.515 ;
        RECT 400.355 -70.205 400.685 -69.875 ;
        RECT 400.355 -71.565 400.685 -71.235 ;
        RECT 400.355 -72.925 400.685 -72.595 ;
        RECT 400.355 -74.285 400.685 -73.955 ;
        RECT 400.355 -75.645 400.685 -75.315 ;
        RECT 400.355 -77.005 400.685 -76.675 ;
        RECT 400.355 -78.365 400.685 -78.035 ;
        RECT 400.355 -79.725 400.685 -79.395 ;
        RECT 400.355 -81.085 400.685 -80.755 ;
        RECT 400.355 -82.445 400.685 -82.115 ;
        RECT 400.355 -83.805 400.685 -83.475 ;
        RECT 400.355 -85.165 400.685 -84.835 ;
        RECT 400.355 -86.525 400.685 -86.195 ;
        RECT 400.355 -87.885 400.685 -87.555 ;
        RECT 400.355 -89.245 400.685 -88.915 ;
        RECT 400.355 -90.605 400.685 -90.275 ;
        RECT 400.355 -91.965 400.685 -91.635 ;
        RECT 400.355 -93.325 400.685 -92.995 ;
        RECT 400.355 -94.685 400.685 -94.355 ;
        RECT 400.355 -96.045 400.685 -95.715 ;
        RECT 400.355 -97.405 400.685 -97.075 ;
        RECT 400.355 -98.765 400.685 -98.435 ;
        RECT 400.355 -100.125 400.685 -99.795 ;
        RECT 400.355 -101.485 400.685 -101.155 ;
        RECT 400.355 -102.845 400.685 -102.515 ;
        RECT 400.355 -104.205 400.685 -103.875 ;
        RECT 400.355 -105.565 400.685 -105.235 ;
        RECT 400.355 -106.925 400.685 -106.595 ;
        RECT 400.355 -108.285 400.685 -107.955 ;
        RECT 400.355 -109.645 400.685 -109.315 ;
        RECT 400.355 -111.005 400.685 -110.675 ;
        RECT 400.355 -112.365 400.685 -112.035 ;
        RECT 400.355 -113.725 400.685 -113.395 ;
        RECT 400.355 -115.085 400.685 -114.755 ;
        RECT 400.355 -116.445 400.685 -116.115 ;
        RECT 400.355 -117.805 400.685 -117.475 ;
        RECT 400.355 -119.165 400.685 -118.835 ;
        RECT 400.355 -120.525 400.685 -120.195 ;
        RECT 400.355 -121.885 400.685 -121.555 ;
        RECT 400.355 -123.245 400.685 -122.915 ;
        RECT 400.355 -124.605 400.685 -124.275 ;
        RECT 400.355 -125.965 400.685 -125.635 ;
        RECT 400.355 -127.325 400.685 -126.995 ;
        RECT 400.355 -128.685 400.685 -128.355 ;
        RECT 400.355 -130.045 400.685 -129.715 ;
        RECT 400.355 -131.405 400.685 -131.075 ;
        RECT 400.355 -132.765 400.685 -132.435 ;
        RECT 400.355 -134.125 400.685 -133.795 ;
        RECT 400.355 -135.485 400.685 -135.155 ;
        RECT 400.355 -136.845 400.685 -136.515 ;
        RECT 400.355 -138.205 400.685 -137.875 ;
        RECT 400.355 -139.565 400.685 -139.235 ;
        RECT 400.355 -140.925 400.685 -140.595 ;
        RECT 400.355 -142.285 400.685 -141.955 ;
        RECT 400.355 -143.645 400.685 -143.315 ;
        RECT 400.355 -145.005 400.685 -144.675 ;
        RECT 400.355 -146.365 400.685 -146.035 ;
        RECT 400.355 -147.725 400.685 -147.395 ;
        RECT 400.355 -149.085 400.685 -148.755 ;
        RECT 400.355 -150.445 400.685 -150.115 ;
        RECT 400.355 -151.805 400.685 -151.475 ;
        RECT 400.355 -153.165 400.685 -152.835 ;
        RECT 400.355 -154.525 400.685 -154.195 ;
        RECT 400.355 -155.885 400.685 -155.555 ;
        RECT 400.355 -157.245 400.685 -156.915 ;
        RECT 400.355 -158.605 400.685 -158.275 ;
        RECT 400.355 -159.965 400.685 -159.635 ;
        RECT 400.355 -161.325 400.685 -160.995 ;
        RECT 400.355 -162.685 400.685 -162.355 ;
        RECT 400.355 -164.045 400.685 -163.715 ;
        RECT 400.355 -165.405 400.685 -165.075 ;
        RECT 400.355 -166.765 400.685 -166.435 ;
        RECT 400.355 -168.125 400.685 -167.795 ;
        RECT 400.355 -169.485 400.685 -169.155 ;
        RECT 400.355 -170.845 400.685 -170.515 ;
        RECT 400.355 -172.205 400.685 -171.875 ;
        RECT 400.355 -173.565 400.685 -173.235 ;
        RECT 400.355 -174.925 400.685 -174.595 ;
        RECT 400.355 -176.285 400.685 -175.955 ;
        RECT 400.355 -177.645 400.685 -177.315 ;
        RECT 400.355 -183.29 400.685 -182.16 ;
        RECT 400.36 -183.405 400.68 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 401.715 244.04 402.045 245.17 ;
        RECT 401.715 239.875 402.045 240.205 ;
        RECT 401.715 238.515 402.045 238.845 ;
        RECT 401.715 237.155 402.045 237.485 ;
        RECT 401.715 235.17 402.045 235.5 ;
        RECT 401.715 232.995 402.045 233.325 ;
        RECT 401.715 231.415 402.045 231.745 ;
        RECT 401.715 230.565 402.045 230.895 ;
        RECT 401.715 228.255 402.045 228.585 ;
        RECT 401.715 227.405 402.045 227.735 ;
        RECT 401.715 225.095 402.045 225.425 ;
        RECT 401.715 224.245 402.045 224.575 ;
        RECT 401.715 221.935 402.045 222.265 ;
        RECT 401.715 221.085 402.045 221.415 ;
        RECT 401.715 218.775 402.045 219.105 ;
        RECT 401.715 217.195 402.045 217.525 ;
        RECT 401.715 216.345 402.045 216.675 ;
        RECT 401.715 214.035 402.045 214.365 ;
        RECT 401.715 213.185 402.045 213.515 ;
        RECT 401.715 210.875 402.045 211.205 ;
        RECT 401.715 210.025 402.045 210.355 ;
        RECT 401.715 207.715 402.045 208.045 ;
        RECT 401.715 206.865 402.045 207.195 ;
        RECT 401.715 204.555 402.045 204.885 ;
        RECT 401.715 202.975 402.045 203.305 ;
        RECT 401.715 202.125 402.045 202.455 ;
        RECT 401.715 199.815 402.045 200.145 ;
        RECT 401.715 198.965 402.045 199.295 ;
        RECT 401.715 196.655 402.045 196.985 ;
        RECT 401.715 195.805 402.045 196.135 ;
        RECT 401.715 193.495 402.045 193.825 ;
        RECT 401.715 192.645 402.045 192.975 ;
        RECT 401.715 190.335 402.045 190.665 ;
        RECT 401.715 188.755 402.045 189.085 ;
        RECT 401.715 187.905 402.045 188.235 ;
        RECT 401.715 185.595 402.045 185.925 ;
        RECT 401.715 184.745 402.045 185.075 ;
        RECT 401.715 182.435 402.045 182.765 ;
        RECT 401.715 181.585 402.045 181.915 ;
        RECT 401.715 179.275 402.045 179.605 ;
        RECT 401.715 178.425 402.045 178.755 ;
        RECT 401.715 176.115 402.045 176.445 ;
        RECT 401.715 174.535 402.045 174.865 ;
        RECT 401.715 173.685 402.045 174.015 ;
        RECT 401.715 171.375 402.045 171.705 ;
        RECT 401.715 170.525 402.045 170.855 ;
        RECT 401.715 168.215 402.045 168.545 ;
        RECT 401.715 167.365 402.045 167.695 ;
        RECT 401.715 165.055 402.045 165.385 ;
        RECT 401.715 164.205 402.045 164.535 ;
        RECT 401.715 161.895 402.045 162.225 ;
        RECT 401.715 160.315 402.045 160.645 ;
        RECT 401.715 159.465 402.045 159.795 ;
        RECT 401.715 157.155 402.045 157.485 ;
        RECT 401.715 156.305 402.045 156.635 ;
        RECT 401.715 153.995 402.045 154.325 ;
        RECT 401.715 153.145 402.045 153.475 ;
        RECT 401.715 150.835 402.045 151.165 ;
        RECT 401.715 149.985 402.045 150.315 ;
        RECT 401.715 147.675 402.045 148.005 ;
        RECT 401.715 146.095 402.045 146.425 ;
        RECT 401.715 145.245 402.045 145.575 ;
        RECT 401.715 142.935 402.045 143.265 ;
        RECT 401.715 142.085 402.045 142.415 ;
        RECT 401.715 139.775 402.045 140.105 ;
        RECT 401.715 138.925 402.045 139.255 ;
        RECT 401.715 136.615 402.045 136.945 ;
        RECT 401.715 135.765 402.045 136.095 ;
        RECT 401.715 133.455 402.045 133.785 ;
        RECT 401.715 131.875 402.045 132.205 ;
        RECT 401.715 131.025 402.045 131.355 ;
        RECT 401.715 128.715 402.045 129.045 ;
        RECT 401.715 127.865 402.045 128.195 ;
        RECT 401.715 125.555 402.045 125.885 ;
        RECT 401.715 124.705 402.045 125.035 ;
        RECT 401.715 122.395 402.045 122.725 ;
        RECT 401.715 121.545 402.045 121.875 ;
        RECT 401.715 119.235 402.045 119.565 ;
        RECT 401.715 117.655 402.045 117.985 ;
        RECT 401.715 116.805 402.045 117.135 ;
        RECT 401.715 114.495 402.045 114.825 ;
        RECT 401.715 113.645 402.045 113.975 ;
        RECT 401.715 111.335 402.045 111.665 ;
        RECT 401.715 110.485 402.045 110.815 ;
        RECT 401.715 108.175 402.045 108.505 ;
        RECT 401.715 107.325 402.045 107.655 ;
        RECT 401.715 105.015 402.045 105.345 ;
        RECT 401.715 103.435 402.045 103.765 ;
        RECT 401.715 102.585 402.045 102.915 ;
        RECT 401.715 100.275 402.045 100.605 ;
        RECT 401.715 99.425 402.045 99.755 ;
        RECT 401.715 97.115 402.045 97.445 ;
        RECT 401.715 96.265 402.045 96.595 ;
        RECT 401.715 93.955 402.045 94.285 ;
        RECT 401.715 93.105 402.045 93.435 ;
        RECT 401.715 90.795 402.045 91.125 ;
        RECT 401.715 89.215 402.045 89.545 ;
        RECT 401.715 88.365 402.045 88.695 ;
        RECT 401.715 86.055 402.045 86.385 ;
        RECT 401.715 85.205 402.045 85.535 ;
        RECT 401.715 82.895 402.045 83.225 ;
        RECT 401.715 82.045 402.045 82.375 ;
        RECT 401.715 79.735 402.045 80.065 ;
        RECT 401.715 78.885 402.045 79.215 ;
        RECT 401.715 76.575 402.045 76.905 ;
        RECT 401.715 74.995 402.045 75.325 ;
        RECT 401.715 74.145 402.045 74.475 ;
        RECT 401.715 71.835 402.045 72.165 ;
        RECT 401.715 70.985 402.045 71.315 ;
        RECT 401.715 68.675 402.045 69.005 ;
        RECT 401.715 67.825 402.045 68.155 ;
        RECT 401.715 65.515 402.045 65.845 ;
        RECT 401.715 64.665 402.045 64.995 ;
        RECT 401.715 62.355 402.045 62.685 ;
        RECT 401.715 60.775 402.045 61.105 ;
        RECT 401.715 59.925 402.045 60.255 ;
        RECT 401.715 57.615 402.045 57.945 ;
        RECT 401.715 56.765 402.045 57.095 ;
        RECT 401.715 54.455 402.045 54.785 ;
        RECT 401.715 53.605 402.045 53.935 ;
        RECT 401.715 51.295 402.045 51.625 ;
        RECT 401.715 50.445 402.045 50.775 ;
        RECT 401.715 48.135 402.045 48.465 ;
        RECT 401.715 46.555 402.045 46.885 ;
        RECT 401.715 45.705 402.045 46.035 ;
        RECT 401.715 43.395 402.045 43.725 ;
        RECT 401.715 42.545 402.045 42.875 ;
        RECT 401.715 40.235 402.045 40.565 ;
        RECT 401.715 39.385 402.045 39.715 ;
        RECT 401.715 37.075 402.045 37.405 ;
        RECT 401.715 36.225 402.045 36.555 ;
        RECT 401.715 33.915 402.045 34.245 ;
        RECT 401.715 32.335 402.045 32.665 ;
        RECT 401.715 31.485 402.045 31.815 ;
        RECT 401.715 29.175 402.045 29.505 ;
        RECT 401.715 28.325 402.045 28.655 ;
        RECT 401.715 26.015 402.045 26.345 ;
        RECT 401.715 25.165 402.045 25.495 ;
        RECT 401.715 22.855 402.045 23.185 ;
        RECT 401.715 22.005 402.045 22.335 ;
        RECT 401.715 19.695 402.045 20.025 ;
        RECT 401.715 18.115 402.045 18.445 ;
        RECT 401.715 17.265 402.045 17.595 ;
        RECT 401.715 14.955 402.045 15.285 ;
        RECT 401.715 14.105 402.045 14.435 ;
        RECT 401.715 11.795 402.045 12.125 ;
        RECT 401.715 10.945 402.045 11.275 ;
        RECT 401.715 8.635 402.045 8.965 ;
        RECT 401.715 7.785 402.045 8.115 ;
        RECT 401.715 5.475 402.045 5.805 ;
        RECT 401.715 3.895 402.045 4.225 ;
        RECT 401.715 3.045 402.045 3.375 ;
        RECT 401.715 0.87 402.045 1.2 ;
        RECT 401.715 -0.845 402.045 -0.515 ;
        RECT 401.715 -2.205 402.045 -1.875 ;
        RECT 401.715 -3.565 402.045 -3.235 ;
        RECT 401.715 -4.925 402.045 -4.595 ;
        RECT 401.715 -6.285 402.045 -5.955 ;
        RECT 401.715 -7.645 402.045 -7.315 ;
        RECT 401.715 -9.005 402.045 -8.675 ;
        RECT 401.715 -10.365 402.045 -10.035 ;
        RECT 401.715 -11.725 402.045 -11.395 ;
        RECT 401.715 -13.085 402.045 -12.755 ;
        RECT 401.715 -14.445 402.045 -14.115 ;
        RECT 401.715 -15.805 402.045 -15.475 ;
        RECT 401.715 -17.165 402.045 -16.835 ;
        RECT 401.715 -18.525 402.045 -18.195 ;
        RECT 401.715 -19.885 402.045 -19.555 ;
        RECT 401.715 -21.245 402.045 -20.915 ;
        RECT 401.715 -22.605 402.045 -22.275 ;
        RECT 401.715 -23.965 402.045 -23.635 ;
        RECT 401.715 -25.325 402.045 -24.995 ;
        RECT 401.715 -26.685 402.045 -26.355 ;
        RECT 401.715 -28.045 402.045 -27.715 ;
        RECT 401.715 -29.405 402.045 -29.075 ;
        RECT 401.715 -30.765 402.045 -30.435 ;
        RECT 401.715 -32.125 402.045 -31.795 ;
        RECT 401.715 -33.485 402.045 -33.155 ;
        RECT 401.715 -34.845 402.045 -34.515 ;
        RECT 401.715 -36.205 402.045 -35.875 ;
        RECT 401.715 -37.565 402.045 -37.235 ;
        RECT 401.715 -38.925 402.045 -38.595 ;
        RECT 401.715 -40.285 402.045 -39.955 ;
        RECT 401.715 -41.645 402.045 -41.315 ;
        RECT 401.715 -43.005 402.045 -42.675 ;
        RECT 401.715 -44.365 402.045 -44.035 ;
        RECT 401.715 -45.725 402.045 -45.395 ;
        RECT 401.715 -47.085 402.045 -46.755 ;
        RECT 401.715 -48.445 402.045 -48.115 ;
        RECT 401.715 -49.805 402.045 -49.475 ;
        RECT 401.715 -51.165 402.045 -50.835 ;
        RECT 401.715 -52.525 402.045 -52.195 ;
        RECT 401.715 -53.885 402.045 -53.555 ;
        RECT 401.715 -55.245 402.045 -54.915 ;
        RECT 401.715 -56.605 402.045 -56.275 ;
        RECT 401.715 -57.965 402.045 -57.635 ;
        RECT 401.715 -59.325 402.045 -58.995 ;
        RECT 401.715 -60.685 402.045 -60.355 ;
        RECT 401.715 -62.045 402.045 -61.715 ;
        RECT 401.715 -63.405 402.045 -63.075 ;
        RECT 401.715 -64.765 402.045 -64.435 ;
        RECT 401.715 -66.125 402.045 -65.795 ;
        RECT 401.715 -67.485 402.045 -67.155 ;
        RECT 401.715 -68.845 402.045 -68.515 ;
        RECT 401.715 -70.205 402.045 -69.875 ;
        RECT 401.715 -71.565 402.045 -71.235 ;
        RECT 401.715 -72.925 402.045 -72.595 ;
        RECT 401.715 -74.285 402.045 -73.955 ;
        RECT 401.715 -75.645 402.045 -75.315 ;
        RECT 401.715 -77.005 402.045 -76.675 ;
        RECT 401.715 -78.365 402.045 -78.035 ;
        RECT 401.715 -79.725 402.045 -79.395 ;
        RECT 401.715 -81.085 402.045 -80.755 ;
        RECT 401.715 -82.445 402.045 -82.115 ;
        RECT 401.715 -83.805 402.045 -83.475 ;
        RECT 401.715 -85.165 402.045 -84.835 ;
        RECT 401.715 -86.525 402.045 -86.195 ;
        RECT 401.715 -87.885 402.045 -87.555 ;
        RECT 401.715 -89.245 402.045 -88.915 ;
        RECT 401.715 -90.605 402.045 -90.275 ;
        RECT 401.715 -91.965 402.045 -91.635 ;
        RECT 401.715 -93.325 402.045 -92.995 ;
        RECT 401.715 -94.685 402.045 -94.355 ;
        RECT 401.715 -96.045 402.045 -95.715 ;
        RECT 401.715 -97.405 402.045 -97.075 ;
        RECT 401.715 -98.765 402.045 -98.435 ;
        RECT 401.715 -100.125 402.045 -99.795 ;
        RECT 401.715 -101.485 402.045 -101.155 ;
        RECT 401.715 -102.845 402.045 -102.515 ;
        RECT 401.715 -104.205 402.045 -103.875 ;
        RECT 401.715 -105.565 402.045 -105.235 ;
        RECT 401.715 -106.925 402.045 -106.595 ;
        RECT 401.715 -108.285 402.045 -107.955 ;
        RECT 401.715 -109.645 402.045 -109.315 ;
        RECT 401.715 -111.005 402.045 -110.675 ;
        RECT 401.715 -112.365 402.045 -112.035 ;
        RECT 401.715 -113.725 402.045 -113.395 ;
        RECT 401.715 -115.085 402.045 -114.755 ;
        RECT 401.715 -116.445 402.045 -116.115 ;
        RECT 401.715 -117.805 402.045 -117.475 ;
        RECT 401.715 -119.165 402.045 -118.835 ;
        RECT 401.715 -120.525 402.045 -120.195 ;
        RECT 401.715 -121.885 402.045 -121.555 ;
        RECT 401.715 -123.245 402.045 -122.915 ;
        RECT 401.715 -124.605 402.045 -124.275 ;
        RECT 401.715 -125.965 402.045 -125.635 ;
        RECT 401.715 -127.325 402.045 -126.995 ;
        RECT 401.715 -128.685 402.045 -128.355 ;
        RECT 401.715 -130.045 402.045 -129.715 ;
        RECT 401.715 -131.405 402.045 -131.075 ;
        RECT 401.715 -132.765 402.045 -132.435 ;
        RECT 401.715 -134.125 402.045 -133.795 ;
        RECT 401.715 -135.485 402.045 -135.155 ;
        RECT 401.715 -136.845 402.045 -136.515 ;
        RECT 401.715 -138.205 402.045 -137.875 ;
        RECT 401.715 -139.565 402.045 -139.235 ;
        RECT 401.715 -140.925 402.045 -140.595 ;
        RECT 401.715 -142.285 402.045 -141.955 ;
        RECT 401.715 -143.645 402.045 -143.315 ;
        RECT 401.715 -145.005 402.045 -144.675 ;
        RECT 401.715 -146.365 402.045 -146.035 ;
        RECT 401.715 -147.725 402.045 -147.395 ;
        RECT 401.715 -149.085 402.045 -148.755 ;
        RECT 401.715 -150.445 402.045 -150.115 ;
        RECT 401.715 -151.805 402.045 -151.475 ;
        RECT 401.715 -153.165 402.045 -152.835 ;
        RECT 401.715 -154.525 402.045 -154.195 ;
        RECT 401.715 -155.885 402.045 -155.555 ;
        RECT 401.715 -157.245 402.045 -156.915 ;
        RECT 401.715 -158.605 402.045 -158.275 ;
        RECT 401.715 -159.965 402.045 -159.635 ;
        RECT 401.715 -161.325 402.045 -160.995 ;
        RECT 401.715 -162.685 402.045 -162.355 ;
        RECT 401.715 -164.045 402.045 -163.715 ;
        RECT 401.715 -165.405 402.045 -165.075 ;
        RECT 401.715 -166.765 402.045 -166.435 ;
        RECT 401.715 -168.125 402.045 -167.795 ;
        RECT 401.715 -169.485 402.045 -169.155 ;
        RECT 401.715 -170.845 402.045 -170.515 ;
        RECT 401.715 -172.205 402.045 -171.875 ;
        RECT 401.715 -173.565 402.045 -173.235 ;
        RECT 401.715 -174.925 402.045 -174.595 ;
        RECT 401.715 -176.285 402.045 -175.955 ;
        RECT 401.715 -177.645 402.045 -177.315 ;
        RECT 401.715 -183.29 402.045 -182.16 ;
        RECT 401.72 -183.405 402.04 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 374.515 244.04 374.845 245.17 ;
        RECT 374.515 239.875 374.845 240.205 ;
        RECT 374.515 238.515 374.845 238.845 ;
        RECT 374.515 237.155 374.845 237.485 ;
        RECT 374.52 237.155 374.84 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 374.515 -96.045 374.845 -95.715 ;
        RECT 374.515 -97.405 374.845 -97.075 ;
        RECT 374.515 -98.765 374.845 -98.435 ;
        RECT 374.515 -100.125 374.845 -99.795 ;
        RECT 374.515 -101.485 374.845 -101.155 ;
        RECT 374.515 -102.845 374.845 -102.515 ;
        RECT 374.515 -104.205 374.845 -103.875 ;
        RECT 374.515 -105.565 374.845 -105.235 ;
        RECT 374.515 -106.925 374.845 -106.595 ;
        RECT 374.515 -108.285 374.845 -107.955 ;
        RECT 374.515 -109.645 374.845 -109.315 ;
        RECT 374.515 -111.005 374.845 -110.675 ;
        RECT 374.515 -112.365 374.845 -112.035 ;
        RECT 374.515 -113.725 374.845 -113.395 ;
        RECT 374.515 -115.085 374.845 -114.755 ;
        RECT 374.515 -116.445 374.845 -116.115 ;
        RECT 374.515 -117.805 374.845 -117.475 ;
        RECT 374.515 -119.165 374.845 -118.835 ;
        RECT 374.515 -120.525 374.845 -120.195 ;
        RECT 374.515 -121.885 374.845 -121.555 ;
        RECT 374.515 -123.245 374.845 -122.915 ;
        RECT 374.515 -124.605 374.845 -124.275 ;
        RECT 374.515 -125.965 374.845 -125.635 ;
        RECT 374.515 -127.325 374.845 -126.995 ;
        RECT 374.515 -128.685 374.845 -128.355 ;
        RECT 374.515 -130.045 374.845 -129.715 ;
        RECT 374.515 -131.405 374.845 -131.075 ;
        RECT 374.515 -132.765 374.845 -132.435 ;
        RECT 374.515 -134.125 374.845 -133.795 ;
        RECT 374.515 -135.485 374.845 -135.155 ;
        RECT 374.515 -136.845 374.845 -136.515 ;
        RECT 374.515 -138.205 374.845 -137.875 ;
        RECT 374.515 -139.565 374.845 -139.235 ;
        RECT 374.515 -140.925 374.845 -140.595 ;
        RECT 374.515 -142.285 374.845 -141.955 ;
        RECT 374.515 -143.645 374.845 -143.315 ;
        RECT 374.515 -145.005 374.845 -144.675 ;
        RECT 374.515 -146.365 374.845 -146.035 ;
        RECT 374.515 -147.725 374.845 -147.395 ;
        RECT 374.515 -149.085 374.845 -148.755 ;
        RECT 374.515 -150.445 374.845 -150.115 ;
        RECT 374.515 -151.805 374.845 -151.475 ;
        RECT 374.515 -153.165 374.845 -152.835 ;
        RECT 374.515 -154.525 374.845 -154.195 ;
        RECT 374.515 -155.885 374.845 -155.555 ;
        RECT 374.515 -157.245 374.845 -156.915 ;
        RECT 374.515 -158.605 374.845 -158.275 ;
        RECT 374.515 -159.965 374.845 -159.635 ;
        RECT 374.515 -161.325 374.845 -160.995 ;
        RECT 374.515 -162.685 374.845 -162.355 ;
        RECT 374.515 -164.045 374.845 -163.715 ;
        RECT 374.515 -165.405 374.845 -165.075 ;
        RECT 374.515 -166.765 374.845 -166.435 ;
        RECT 374.515 -168.125 374.845 -167.795 ;
        RECT 374.515 -169.485 374.845 -169.155 ;
        RECT 374.515 -170.845 374.845 -170.515 ;
        RECT 374.515 -172.205 374.845 -171.875 ;
        RECT 374.515 -173.565 374.845 -173.235 ;
        RECT 374.515 -174.925 374.845 -174.595 ;
        RECT 374.515 -176.285 374.845 -175.955 ;
        RECT 374.515 -177.645 374.845 -177.315 ;
        RECT 374.515 -183.29 374.845 -182.16 ;
        RECT 374.52 -183.405 374.84 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 374.76 -94.075 375.09 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 375.875 244.04 376.205 245.17 ;
        RECT 375.875 239.875 376.205 240.205 ;
        RECT 375.875 238.515 376.205 238.845 ;
        RECT 375.875 237.155 376.205 237.485 ;
        RECT 375.88 237.155 376.2 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 377.235 244.04 377.565 245.17 ;
        RECT 377.235 239.875 377.565 240.205 ;
        RECT 377.235 238.515 377.565 238.845 ;
        RECT 377.235 237.155 377.565 237.485 ;
        RECT 377.24 237.155 377.56 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 377.235 -0.845 377.565 -0.515 ;
        RECT 377.235 -2.205 377.565 -1.875 ;
        RECT 377.235 -3.565 377.565 -3.235 ;
        RECT 377.24 -3.565 377.56 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 378.595 244.04 378.925 245.17 ;
        RECT 378.595 239.875 378.925 240.205 ;
        RECT 378.595 238.515 378.925 238.845 ;
        RECT 378.595 237.155 378.925 237.485 ;
        RECT 378.6 237.155 378.92 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 378.595 -0.845 378.925 -0.515 ;
        RECT 378.595 -2.205 378.925 -1.875 ;
        RECT 378.595 -3.565 378.925 -3.235 ;
        RECT 378.6 -3.565 378.92 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 378.595 -91.965 378.925 -91.635 ;
        RECT 378.595 -93.325 378.925 -92.995 ;
        RECT 378.595 -94.685 378.925 -94.355 ;
        RECT 378.595 -96.045 378.925 -95.715 ;
        RECT 378.595 -97.405 378.925 -97.075 ;
        RECT 378.595 -98.765 378.925 -98.435 ;
        RECT 378.595 -100.125 378.925 -99.795 ;
        RECT 378.595 -101.485 378.925 -101.155 ;
        RECT 378.595 -102.845 378.925 -102.515 ;
        RECT 378.595 -104.205 378.925 -103.875 ;
        RECT 378.595 -105.565 378.925 -105.235 ;
        RECT 378.595 -106.925 378.925 -106.595 ;
        RECT 378.595 -108.285 378.925 -107.955 ;
        RECT 378.595 -109.645 378.925 -109.315 ;
        RECT 378.595 -111.005 378.925 -110.675 ;
        RECT 378.595 -112.365 378.925 -112.035 ;
        RECT 378.595 -113.725 378.925 -113.395 ;
        RECT 378.595 -115.085 378.925 -114.755 ;
        RECT 378.595 -116.445 378.925 -116.115 ;
        RECT 378.595 -117.805 378.925 -117.475 ;
        RECT 378.595 -119.165 378.925 -118.835 ;
        RECT 378.595 -120.525 378.925 -120.195 ;
        RECT 378.595 -121.885 378.925 -121.555 ;
        RECT 378.595 -123.245 378.925 -122.915 ;
        RECT 378.595 -124.605 378.925 -124.275 ;
        RECT 378.595 -125.965 378.925 -125.635 ;
        RECT 378.595 -127.325 378.925 -126.995 ;
        RECT 378.595 -128.685 378.925 -128.355 ;
        RECT 378.595 -130.045 378.925 -129.715 ;
        RECT 378.595 -131.405 378.925 -131.075 ;
        RECT 378.595 -132.765 378.925 -132.435 ;
        RECT 378.595 -134.125 378.925 -133.795 ;
        RECT 378.595 -135.485 378.925 -135.155 ;
        RECT 378.595 -136.845 378.925 -136.515 ;
        RECT 378.595 -138.205 378.925 -137.875 ;
        RECT 378.595 -139.565 378.925 -139.235 ;
        RECT 378.595 -140.925 378.925 -140.595 ;
        RECT 378.595 -142.285 378.925 -141.955 ;
        RECT 378.595 -143.645 378.925 -143.315 ;
        RECT 378.595 -145.005 378.925 -144.675 ;
        RECT 378.595 -146.365 378.925 -146.035 ;
        RECT 378.595 -147.725 378.925 -147.395 ;
        RECT 378.595 -149.085 378.925 -148.755 ;
        RECT 378.595 -150.445 378.925 -150.115 ;
        RECT 378.595 -151.805 378.925 -151.475 ;
        RECT 378.595 -153.165 378.925 -152.835 ;
        RECT 378.595 -154.525 378.925 -154.195 ;
        RECT 378.595 -155.885 378.925 -155.555 ;
        RECT 378.595 -157.245 378.925 -156.915 ;
        RECT 378.595 -158.605 378.925 -158.275 ;
        RECT 378.595 -159.965 378.925 -159.635 ;
        RECT 378.595 -161.325 378.925 -160.995 ;
        RECT 378.595 -162.685 378.925 -162.355 ;
        RECT 378.595 -164.045 378.925 -163.715 ;
        RECT 378.595 -165.405 378.925 -165.075 ;
        RECT 378.595 -166.765 378.925 -166.435 ;
        RECT 378.595 -168.125 378.925 -167.795 ;
        RECT 378.595 -169.485 378.925 -169.155 ;
        RECT 378.595 -170.845 378.925 -170.515 ;
        RECT 378.595 -172.205 378.925 -171.875 ;
        RECT 378.595 -173.565 378.925 -173.235 ;
        RECT 378.595 -174.925 378.925 -174.595 ;
        RECT 378.595 -176.285 378.925 -175.955 ;
        RECT 378.595 -177.645 378.925 -177.315 ;
        RECT 378.595 -183.29 378.925 -182.16 ;
        RECT 378.6 -183.405 378.92 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 379.955 244.04 380.285 245.17 ;
        RECT 379.955 239.875 380.285 240.205 ;
        RECT 379.955 238.515 380.285 238.845 ;
        RECT 379.955 237.155 380.285 237.485 ;
        RECT 379.96 237.155 380.28 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 379.955 -0.845 380.285 -0.515 ;
        RECT 379.955 -2.205 380.285 -1.875 ;
        RECT 379.955 -3.565 380.285 -3.235 ;
        RECT 379.96 -3.565 380.28 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 379.955 -91.965 380.285 -91.635 ;
        RECT 379.955 -93.325 380.285 -92.995 ;
        RECT 379.955 -94.685 380.285 -94.355 ;
        RECT 379.955 -96.045 380.285 -95.715 ;
        RECT 379.955 -97.405 380.285 -97.075 ;
        RECT 379.955 -98.765 380.285 -98.435 ;
        RECT 379.955 -100.125 380.285 -99.795 ;
        RECT 379.955 -101.485 380.285 -101.155 ;
        RECT 379.955 -102.845 380.285 -102.515 ;
        RECT 379.955 -104.205 380.285 -103.875 ;
        RECT 379.955 -105.565 380.285 -105.235 ;
        RECT 379.955 -106.925 380.285 -106.595 ;
        RECT 379.955 -108.285 380.285 -107.955 ;
        RECT 379.955 -109.645 380.285 -109.315 ;
        RECT 379.955 -111.005 380.285 -110.675 ;
        RECT 379.955 -112.365 380.285 -112.035 ;
        RECT 379.955 -113.725 380.285 -113.395 ;
        RECT 379.955 -115.085 380.285 -114.755 ;
        RECT 379.955 -116.445 380.285 -116.115 ;
        RECT 379.955 -117.805 380.285 -117.475 ;
        RECT 379.955 -119.165 380.285 -118.835 ;
        RECT 379.955 -120.525 380.285 -120.195 ;
        RECT 379.955 -121.885 380.285 -121.555 ;
        RECT 379.955 -123.245 380.285 -122.915 ;
        RECT 379.955 -124.605 380.285 -124.275 ;
        RECT 379.955 -125.965 380.285 -125.635 ;
        RECT 379.955 -127.325 380.285 -126.995 ;
        RECT 379.955 -128.685 380.285 -128.355 ;
        RECT 379.955 -130.045 380.285 -129.715 ;
        RECT 379.955 -131.405 380.285 -131.075 ;
        RECT 379.955 -132.765 380.285 -132.435 ;
        RECT 379.955 -134.125 380.285 -133.795 ;
        RECT 379.955 -135.485 380.285 -135.155 ;
        RECT 379.955 -136.845 380.285 -136.515 ;
        RECT 379.955 -138.205 380.285 -137.875 ;
        RECT 379.955 -139.565 380.285 -139.235 ;
        RECT 379.955 -140.925 380.285 -140.595 ;
        RECT 379.955 -142.285 380.285 -141.955 ;
        RECT 379.955 -143.645 380.285 -143.315 ;
        RECT 379.955 -145.005 380.285 -144.675 ;
        RECT 379.955 -146.365 380.285 -146.035 ;
        RECT 379.955 -147.725 380.285 -147.395 ;
        RECT 379.955 -149.085 380.285 -148.755 ;
        RECT 379.955 -150.445 380.285 -150.115 ;
        RECT 379.955 -151.805 380.285 -151.475 ;
        RECT 379.955 -153.165 380.285 -152.835 ;
        RECT 379.955 -154.525 380.285 -154.195 ;
        RECT 379.955 -155.885 380.285 -155.555 ;
        RECT 379.955 -157.245 380.285 -156.915 ;
        RECT 379.955 -158.605 380.285 -158.275 ;
        RECT 379.955 -159.965 380.285 -159.635 ;
        RECT 379.955 -161.325 380.285 -160.995 ;
        RECT 379.955 -162.685 380.285 -162.355 ;
        RECT 379.955 -164.045 380.285 -163.715 ;
        RECT 379.955 -165.405 380.285 -165.075 ;
        RECT 379.955 -166.765 380.285 -166.435 ;
        RECT 379.955 -168.125 380.285 -167.795 ;
        RECT 379.955 -169.485 380.285 -169.155 ;
        RECT 379.955 -170.845 380.285 -170.515 ;
        RECT 379.955 -172.205 380.285 -171.875 ;
        RECT 379.955 -173.565 380.285 -173.235 ;
        RECT 379.955 -174.925 380.285 -174.595 ;
        RECT 379.955 -176.285 380.285 -175.955 ;
        RECT 379.955 -177.645 380.285 -177.315 ;
        RECT 379.955 -183.29 380.285 -182.16 ;
        RECT 379.96 -183.405 380.28 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 380.86 -94.075 381.19 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 381.315 244.04 381.645 245.17 ;
        RECT 381.315 239.875 381.645 240.205 ;
        RECT 381.315 238.515 381.645 238.845 ;
        RECT 381.315 237.155 381.645 237.485 ;
        RECT 381.32 237.155 381.64 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 381.315 -96.045 381.645 -95.715 ;
        RECT 381.315 -97.405 381.645 -97.075 ;
        RECT 381.315 -98.765 381.645 -98.435 ;
        RECT 381.315 -100.125 381.645 -99.795 ;
        RECT 381.315 -101.485 381.645 -101.155 ;
        RECT 381.315 -102.845 381.645 -102.515 ;
        RECT 381.315 -104.205 381.645 -103.875 ;
        RECT 381.315 -105.565 381.645 -105.235 ;
        RECT 381.315 -106.925 381.645 -106.595 ;
        RECT 381.315 -108.285 381.645 -107.955 ;
        RECT 381.315 -109.645 381.645 -109.315 ;
        RECT 381.315 -111.005 381.645 -110.675 ;
        RECT 381.315 -112.365 381.645 -112.035 ;
        RECT 381.315 -113.725 381.645 -113.395 ;
        RECT 381.315 -115.085 381.645 -114.755 ;
        RECT 381.315 -116.445 381.645 -116.115 ;
        RECT 381.315 -117.805 381.645 -117.475 ;
        RECT 381.315 -119.165 381.645 -118.835 ;
        RECT 381.315 -120.525 381.645 -120.195 ;
        RECT 381.315 -121.885 381.645 -121.555 ;
        RECT 381.315 -123.245 381.645 -122.915 ;
        RECT 381.315 -124.605 381.645 -124.275 ;
        RECT 381.315 -125.965 381.645 -125.635 ;
        RECT 381.315 -127.325 381.645 -126.995 ;
        RECT 381.315 -128.685 381.645 -128.355 ;
        RECT 381.315 -130.045 381.645 -129.715 ;
        RECT 381.315 -131.405 381.645 -131.075 ;
        RECT 381.315 -132.765 381.645 -132.435 ;
        RECT 381.315 -134.125 381.645 -133.795 ;
        RECT 381.315 -135.485 381.645 -135.155 ;
        RECT 381.315 -136.845 381.645 -136.515 ;
        RECT 381.315 -138.205 381.645 -137.875 ;
        RECT 381.315 -139.565 381.645 -139.235 ;
        RECT 381.315 -140.925 381.645 -140.595 ;
        RECT 381.315 -142.285 381.645 -141.955 ;
        RECT 381.315 -143.645 381.645 -143.315 ;
        RECT 381.315 -145.005 381.645 -144.675 ;
        RECT 381.315 -146.365 381.645 -146.035 ;
        RECT 381.315 -147.725 381.645 -147.395 ;
        RECT 381.315 -149.085 381.645 -148.755 ;
        RECT 381.315 -150.445 381.645 -150.115 ;
        RECT 381.315 -151.805 381.645 -151.475 ;
        RECT 381.315 -153.165 381.645 -152.835 ;
        RECT 381.315 -154.525 381.645 -154.195 ;
        RECT 381.315 -155.885 381.645 -155.555 ;
        RECT 381.315 -157.245 381.645 -156.915 ;
        RECT 381.315 -158.605 381.645 -158.275 ;
        RECT 381.315 -159.965 381.645 -159.635 ;
        RECT 381.315 -161.325 381.645 -160.995 ;
        RECT 381.315 -162.685 381.645 -162.355 ;
        RECT 381.315 -164.045 381.645 -163.715 ;
        RECT 381.315 -165.405 381.645 -165.075 ;
        RECT 381.315 -166.765 381.645 -166.435 ;
        RECT 381.315 -168.125 381.645 -167.795 ;
        RECT 381.315 -169.485 381.645 -169.155 ;
        RECT 381.315 -170.845 381.645 -170.515 ;
        RECT 381.315 -172.205 381.645 -171.875 ;
        RECT 381.315 -173.565 381.645 -173.235 ;
        RECT 381.315 -174.925 381.645 -174.595 ;
        RECT 381.315 -176.285 381.645 -175.955 ;
        RECT 381.315 -177.645 381.645 -177.315 ;
        RECT 381.315 -183.29 381.645 -182.16 ;
        RECT 381.32 -183.405 381.64 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 382.675 244.04 383.005 245.17 ;
        RECT 382.675 239.875 383.005 240.205 ;
        RECT 382.675 238.515 383.005 238.845 ;
        RECT 382.675 237.155 383.005 237.485 ;
        RECT 382.68 237.155 383 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 382.675 -0.845 383.005 -0.515 ;
        RECT 382.675 -2.205 383.005 -1.875 ;
        RECT 382.675 -3.565 383.005 -3.235 ;
        RECT 382.68 -3.565 383 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 384.035 244.04 384.365 245.17 ;
        RECT 384.035 239.875 384.365 240.205 ;
        RECT 384.035 238.515 384.365 238.845 ;
        RECT 384.035 237.155 384.365 237.485 ;
        RECT 384.04 237.155 384.36 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 384.035 -0.845 384.365 -0.515 ;
        RECT 384.035 -2.205 384.365 -1.875 ;
        RECT 384.035 -3.565 384.365 -3.235 ;
        RECT 384.04 -3.565 384.36 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 385.395 244.04 385.725 245.17 ;
        RECT 385.395 239.875 385.725 240.205 ;
        RECT 385.395 238.515 385.725 238.845 ;
        RECT 385.395 237.155 385.725 237.485 ;
        RECT 385.4 237.155 385.72 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 385.395 -0.845 385.725 -0.515 ;
        RECT 385.395 -2.205 385.725 -1.875 ;
        RECT 385.395 -3.565 385.725 -3.235 ;
        RECT 385.4 -3.565 385.72 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 385.395 -91.965 385.725 -91.635 ;
        RECT 385.395 -93.325 385.725 -92.995 ;
        RECT 385.395 -94.685 385.725 -94.355 ;
        RECT 385.395 -96.045 385.725 -95.715 ;
        RECT 385.395 -97.405 385.725 -97.075 ;
        RECT 385.395 -98.765 385.725 -98.435 ;
        RECT 385.395 -100.125 385.725 -99.795 ;
        RECT 385.395 -101.485 385.725 -101.155 ;
        RECT 385.395 -102.845 385.725 -102.515 ;
        RECT 385.395 -104.205 385.725 -103.875 ;
        RECT 385.395 -105.565 385.725 -105.235 ;
        RECT 385.395 -106.925 385.725 -106.595 ;
        RECT 385.395 -108.285 385.725 -107.955 ;
        RECT 385.395 -109.645 385.725 -109.315 ;
        RECT 385.395 -111.005 385.725 -110.675 ;
        RECT 385.395 -112.365 385.725 -112.035 ;
        RECT 385.395 -113.725 385.725 -113.395 ;
        RECT 385.395 -115.085 385.725 -114.755 ;
        RECT 385.395 -116.445 385.725 -116.115 ;
        RECT 385.395 -117.805 385.725 -117.475 ;
        RECT 385.395 -119.165 385.725 -118.835 ;
        RECT 385.395 -120.525 385.725 -120.195 ;
        RECT 385.395 -121.885 385.725 -121.555 ;
        RECT 385.395 -123.245 385.725 -122.915 ;
        RECT 385.395 -124.605 385.725 -124.275 ;
        RECT 385.395 -125.965 385.725 -125.635 ;
        RECT 385.395 -127.325 385.725 -126.995 ;
        RECT 385.395 -128.685 385.725 -128.355 ;
        RECT 385.395 -130.045 385.725 -129.715 ;
        RECT 385.395 -131.405 385.725 -131.075 ;
        RECT 385.395 -132.765 385.725 -132.435 ;
        RECT 385.395 -134.125 385.725 -133.795 ;
        RECT 385.395 -135.485 385.725 -135.155 ;
        RECT 385.395 -136.845 385.725 -136.515 ;
        RECT 385.395 -138.205 385.725 -137.875 ;
        RECT 385.395 -139.565 385.725 -139.235 ;
        RECT 385.395 -140.925 385.725 -140.595 ;
        RECT 385.395 -142.285 385.725 -141.955 ;
        RECT 385.395 -143.645 385.725 -143.315 ;
        RECT 385.395 -145.005 385.725 -144.675 ;
        RECT 385.395 -146.365 385.725 -146.035 ;
        RECT 385.395 -147.725 385.725 -147.395 ;
        RECT 385.395 -149.085 385.725 -148.755 ;
        RECT 385.395 -150.445 385.725 -150.115 ;
        RECT 385.395 -151.805 385.725 -151.475 ;
        RECT 385.395 -153.165 385.725 -152.835 ;
        RECT 385.395 -154.525 385.725 -154.195 ;
        RECT 385.395 -155.885 385.725 -155.555 ;
        RECT 385.395 -157.245 385.725 -156.915 ;
        RECT 385.395 -158.605 385.725 -158.275 ;
        RECT 385.395 -159.965 385.725 -159.635 ;
        RECT 385.395 -161.325 385.725 -160.995 ;
        RECT 385.395 -162.685 385.725 -162.355 ;
        RECT 385.395 -164.045 385.725 -163.715 ;
        RECT 385.395 -165.405 385.725 -165.075 ;
        RECT 385.395 -166.765 385.725 -166.435 ;
        RECT 385.395 -168.125 385.725 -167.795 ;
        RECT 385.395 -169.485 385.725 -169.155 ;
        RECT 385.395 -170.845 385.725 -170.515 ;
        RECT 385.395 -172.205 385.725 -171.875 ;
        RECT 385.395 -173.565 385.725 -173.235 ;
        RECT 385.395 -174.925 385.725 -174.595 ;
        RECT 385.395 -176.285 385.725 -175.955 ;
        RECT 385.395 -177.645 385.725 -177.315 ;
        RECT 385.395 -183.29 385.725 -182.16 ;
        RECT 385.4 -183.405 385.72 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 386.755 244.04 387.085 245.17 ;
        RECT 386.755 239.875 387.085 240.205 ;
        RECT 386.755 238.515 387.085 238.845 ;
        RECT 386.755 237.155 387.085 237.485 ;
        RECT 386.76 237.155 387.08 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 386.755 -96.045 387.085 -95.715 ;
        RECT 386.755 -97.405 387.085 -97.075 ;
        RECT 386.755 -98.765 387.085 -98.435 ;
        RECT 386.755 -100.125 387.085 -99.795 ;
        RECT 386.755 -101.485 387.085 -101.155 ;
        RECT 386.755 -102.845 387.085 -102.515 ;
        RECT 386.755 -104.205 387.085 -103.875 ;
        RECT 386.755 -105.565 387.085 -105.235 ;
        RECT 386.755 -106.925 387.085 -106.595 ;
        RECT 386.755 -108.285 387.085 -107.955 ;
        RECT 386.755 -109.645 387.085 -109.315 ;
        RECT 386.755 -111.005 387.085 -110.675 ;
        RECT 386.755 -112.365 387.085 -112.035 ;
        RECT 386.755 -113.725 387.085 -113.395 ;
        RECT 386.755 -115.085 387.085 -114.755 ;
        RECT 386.755 -116.445 387.085 -116.115 ;
        RECT 386.755 -117.805 387.085 -117.475 ;
        RECT 386.755 -119.165 387.085 -118.835 ;
        RECT 386.755 -120.525 387.085 -120.195 ;
        RECT 386.755 -121.885 387.085 -121.555 ;
        RECT 386.755 -123.245 387.085 -122.915 ;
        RECT 386.755 -124.605 387.085 -124.275 ;
        RECT 386.755 -125.965 387.085 -125.635 ;
        RECT 386.755 -127.325 387.085 -126.995 ;
        RECT 386.755 -128.685 387.085 -128.355 ;
        RECT 386.755 -130.045 387.085 -129.715 ;
        RECT 386.755 -131.405 387.085 -131.075 ;
        RECT 386.755 -132.765 387.085 -132.435 ;
        RECT 386.755 -134.125 387.085 -133.795 ;
        RECT 386.755 -135.485 387.085 -135.155 ;
        RECT 386.755 -136.845 387.085 -136.515 ;
        RECT 386.755 -138.205 387.085 -137.875 ;
        RECT 386.755 -139.565 387.085 -139.235 ;
        RECT 386.755 -140.925 387.085 -140.595 ;
        RECT 386.755 -142.285 387.085 -141.955 ;
        RECT 386.755 -143.645 387.085 -143.315 ;
        RECT 386.755 -145.005 387.085 -144.675 ;
        RECT 386.755 -146.365 387.085 -146.035 ;
        RECT 386.755 -147.725 387.085 -147.395 ;
        RECT 386.755 -149.085 387.085 -148.755 ;
        RECT 386.755 -150.445 387.085 -150.115 ;
        RECT 386.755 -151.805 387.085 -151.475 ;
        RECT 386.755 -153.165 387.085 -152.835 ;
        RECT 386.755 -154.525 387.085 -154.195 ;
        RECT 386.755 -155.885 387.085 -155.555 ;
        RECT 386.755 -157.245 387.085 -156.915 ;
        RECT 386.755 -158.605 387.085 -158.275 ;
        RECT 386.755 -159.965 387.085 -159.635 ;
        RECT 386.755 -161.325 387.085 -160.995 ;
        RECT 386.755 -162.685 387.085 -162.355 ;
        RECT 386.755 -164.045 387.085 -163.715 ;
        RECT 386.755 -165.405 387.085 -165.075 ;
        RECT 386.755 -166.765 387.085 -166.435 ;
        RECT 386.755 -168.125 387.085 -167.795 ;
        RECT 386.755 -169.485 387.085 -169.155 ;
        RECT 386.755 -170.845 387.085 -170.515 ;
        RECT 386.755 -172.205 387.085 -171.875 ;
        RECT 386.755 -173.565 387.085 -173.235 ;
        RECT 386.755 -174.925 387.085 -174.595 ;
        RECT 386.755 -176.285 387.085 -175.955 ;
        RECT 386.755 -177.645 387.085 -177.315 ;
        RECT 386.755 -183.29 387.085 -182.16 ;
        RECT 386.76 -183.405 387.08 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 386.96 -94.075 387.29 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 388.115 244.04 388.445 245.17 ;
        RECT 388.115 239.875 388.445 240.205 ;
        RECT 388.115 238.515 388.445 238.845 ;
        RECT 388.115 237.155 388.445 237.485 ;
        RECT 388.12 237.155 388.44 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 389.475 244.04 389.805 245.17 ;
        RECT 389.475 239.875 389.805 240.205 ;
        RECT 389.475 238.515 389.805 238.845 ;
        RECT 389.475 237.155 389.805 237.485 ;
        RECT 389.48 237.155 389.8 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 389.475 -0.845 389.805 -0.515 ;
        RECT 389.475 -2.205 389.805 -1.875 ;
        RECT 389.475 -3.565 389.805 -3.235 ;
        RECT 389.48 -3.565 389.8 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 390.835 244.04 391.165 245.17 ;
        RECT 390.835 239.875 391.165 240.205 ;
        RECT 390.835 238.515 391.165 238.845 ;
        RECT 390.835 237.155 391.165 237.485 ;
        RECT 390.84 237.155 391.16 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 390.835 -0.845 391.165 -0.515 ;
        RECT 390.835 -2.205 391.165 -1.875 ;
        RECT 390.835 -3.565 391.165 -3.235 ;
        RECT 390.84 -3.565 391.16 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 390.835 -91.965 391.165 -91.635 ;
        RECT 390.835 -93.325 391.165 -92.995 ;
        RECT 390.835 -94.685 391.165 -94.355 ;
        RECT 390.835 -96.045 391.165 -95.715 ;
        RECT 390.835 -97.405 391.165 -97.075 ;
        RECT 390.835 -98.765 391.165 -98.435 ;
        RECT 390.835 -100.125 391.165 -99.795 ;
        RECT 390.835 -101.485 391.165 -101.155 ;
        RECT 390.835 -102.845 391.165 -102.515 ;
        RECT 390.835 -104.205 391.165 -103.875 ;
        RECT 390.835 -105.565 391.165 -105.235 ;
        RECT 390.835 -106.925 391.165 -106.595 ;
        RECT 390.835 -108.285 391.165 -107.955 ;
        RECT 390.835 -109.645 391.165 -109.315 ;
        RECT 390.835 -111.005 391.165 -110.675 ;
        RECT 390.835 -112.365 391.165 -112.035 ;
        RECT 390.835 -113.725 391.165 -113.395 ;
        RECT 390.835 -115.085 391.165 -114.755 ;
        RECT 390.835 -116.445 391.165 -116.115 ;
        RECT 390.835 -117.805 391.165 -117.475 ;
        RECT 390.835 -119.165 391.165 -118.835 ;
        RECT 390.835 -120.525 391.165 -120.195 ;
        RECT 390.835 -121.885 391.165 -121.555 ;
        RECT 390.835 -123.245 391.165 -122.915 ;
        RECT 390.835 -124.605 391.165 -124.275 ;
        RECT 390.835 -125.965 391.165 -125.635 ;
        RECT 390.835 -127.325 391.165 -126.995 ;
        RECT 390.835 -128.685 391.165 -128.355 ;
        RECT 390.835 -130.045 391.165 -129.715 ;
        RECT 390.835 -131.405 391.165 -131.075 ;
        RECT 390.835 -132.765 391.165 -132.435 ;
        RECT 390.835 -134.125 391.165 -133.795 ;
        RECT 390.835 -135.485 391.165 -135.155 ;
        RECT 390.835 -136.845 391.165 -136.515 ;
        RECT 390.835 -138.205 391.165 -137.875 ;
        RECT 390.835 -139.565 391.165 -139.235 ;
        RECT 390.835 -140.925 391.165 -140.595 ;
        RECT 390.835 -142.285 391.165 -141.955 ;
        RECT 390.835 -143.645 391.165 -143.315 ;
        RECT 390.835 -145.005 391.165 -144.675 ;
        RECT 390.835 -146.365 391.165 -146.035 ;
        RECT 390.835 -147.725 391.165 -147.395 ;
        RECT 390.835 -149.085 391.165 -148.755 ;
        RECT 390.835 -150.445 391.165 -150.115 ;
        RECT 390.835 -151.805 391.165 -151.475 ;
        RECT 390.835 -153.165 391.165 -152.835 ;
        RECT 390.835 -154.525 391.165 -154.195 ;
        RECT 390.835 -155.885 391.165 -155.555 ;
        RECT 390.835 -157.245 391.165 -156.915 ;
        RECT 390.835 -158.605 391.165 -158.275 ;
        RECT 390.835 -159.965 391.165 -159.635 ;
        RECT 390.835 -161.325 391.165 -160.995 ;
        RECT 390.835 -162.685 391.165 -162.355 ;
        RECT 390.835 -164.045 391.165 -163.715 ;
        RECT 390.835 -165.405 391.165 -165.075 ;
        RECT 390.835 -166.765 391.165 -166.435 ;
        RECT 390.835 -168.125 391.165 -167.795 ;
        RECT 390.835 -169.485 391.165 -169.155 ;
        RECT 390.835 -170.845 391.165 -170.515 ;
        RECT 390.835 -172.205 391.165 -171.875 ;
        RECT 390.835 -173.565 391.165 -173.235 ;
        RECT 390.835 -174.925 391.165 -174.595 ;
        RECT 390.835 -176.285 391.165 -175.955 ;
        RECT 390.835 -177.645 391.165 -177.315 ;
        RECT 390.835 -183.29 391.165 -182.16 ;
        RECT 390.84 -183.405 391.16 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 392.195 244.04 392.525 245.17 ;
        RECT 392.195 239.875 392.525 240.205 ;
        RECT 392.195 238.515 392.525 238.845 ;
        RECT 392.195 237.155 392.525 237.485 ;
        RECT 392.2 237.155 392.52 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 392.195 -0.845 392.525 -0.515 ;
        RECT 392.195 -2.205 392.525 -1.875 ;
        RECT 392.195 -3.565 392.525 -3.235 ;
        RECT 392.2 -3.565 392.52 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 392.195 -91.965 392.525 -91.635 ;
        RECT 392.195 -93.325 392.525 -92.995 ;
        RECT 392.195 -94.685 392.525 -94.355 ;
        RECT 392.195 -96.045 392.525 -95.715 ;
        RECT 392.195 -97.405 392.525 -97.075 ;
        RECT 392.195 -98.765 392.525 -98.435 ;
        RECT 392.195 -100.125 392.525 -99.795 ;
        RECT 392.195 -101.485 392.525 -101.155 ;
        RECT 392.195 -102.845 392.525 -102.515 ;
        RECT 392.195 -104.205 392.525 -103.875 ;
        RECT 392.195 -105.565 392.525 -105.235 ;
        RECT 392.195 -106.925 392.525 -106.595 ;
        RECT 392.195 -108.285 392.525 -107.955 ;
        RECT 392.195 -109.645 392.525 -109.315 ;
        RECT 392.195 -111.005 392.525 -110.675 ;
        RECT 392.195 -112.365 392.525 -112.035 ;
        RECT 392.195 -113.725 392.525 -113.395 ;
        RECT 392.195 -115.085 392.525 -114.755 ;
        RECT 392.195 -116.445 392.525 -116.115 ;
        RECT 392.195 -117.805 392.525 -117.475 ;
        RECT 392.195 -119.165 392.525 -118.835 ;
        RECT 392.195 -120.525 392.525 -120.195 ;
        RECT 392.195 -121.885 392.525 -121.555 ;
        RECT 392.195 -123.245 392.525 -122.915 ;
        RECT 392.195 -124.605 392.525 -124.275 ;
        RECT 392.195 -125.965 392.525 -125.635 ;
        RECT 392.195 -127.325 392.525 -126.995 ;
        RECT 392.195 -128.685 392.525 -128.355 ;
        RECT 392.195 -130.045 392.525 -129.715 ;
        RECT 392.195 -131.405 392.525 -131.075 ;
        RECT 392.195 -132.765 392.525 -132.435 ;
        RECT 392.195 -134.125 392.525 -133.795 ;
        RECT 392.195 -135.485 392.525 -135.155 ;
        RECT 392.195 -136.845 392.525 -136.515 ;
        RECT 392.195 -138.205 392.525 -137.875 ;
        RECT 392.195 -139.565 392.525 -139.235 ;
        RECT 392.195 -140.925 392.525 -140.595 ;
        RECT 392.195 -142.285 392.525 -141.955 ;
        RECT 392.195 -143.645 392.525 -143.315 ;
        RECT 392.195 -145.005 392.525 -144.675 ;
        RECT 392.195 -146.365 392.525 -146.035 ;
        RECT 392.195 -147.725 392.525 -147.395 ;
        RECT 392.195 -149.085 392.525 -148.755 ;
        RECT 392.195 -150.445 392.525 -150.115 ;
        RECT 392.195 -151.805 392.525 -151.475 ;
        RECT 392.195 -153.165 392.525 -152.835 ;
        RECT 392.195 -154.525 392.525 -154.195 ;
        RECT 392.195 -155.885 392.525 -155.555 ;
        RECT 392.195 -157.245 392.525 -156.915 ;
        RECT 392.195 -158.605 392.525 -158.275 ;
        RECT 392.195 -159.965 392.525 -159.635 ;
        RECT 392.195 -161.325 392.525 -160.995 ;
        RECT 392.195 -162.685 392.525 -162.355 ;
        RECT 392.195 -164.045 392.525 -163.715 ;
        RECT 392.195 -165.405 392.525 -165.075 ;
        RECT 392.195 -166.765 392.525 -166.435 ;
        RECT 392.195 -168.125 392.525 -167.795 ;
        RECT 392.195 -169.485 392.525 -169.155 ;
        RECT 392.195 -170.845 392.525 -170.515 ;
        RECT 392.195 -172.205 392.525 -171.875 ;
        RECT 392.195 -173.565 392.525 -173.235 ;
        RECT 392.195 -174.925 392.525 -174.595 ;
        RECT 392.195 -176.285 392.525 -175.955 ;
        RECT 392.195 -177.645 392.525 -177.315 ;
        RECT 392.195 -183.29 392.525 -182.16 ;
        RECT 392.2 -183.405 392.52 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 393.555 244.04 393.885 245.17 ;
        RECT 393.555 239.875 393.885 240.205 ;
        RECT 393.555 238.515 393.885 238.845 ;
        RECT 393.555 237.155 393.885 237.485 ;
        RECT 393.56 237.155 393.88 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 393.555 -96.045 393.885 -95.715 ;
        RECT 393.555 -97.405 393.885 -97.075 ;
        RECT 393.555 -98.765 393.885 -98.435 ;
        RECT 393.555 -100.125 393.885 -99.795 ;
        RECT 393.555 -101.485 393.885 -101.155 ;
        RECT 393.555 -102.845 393.885 -102.515 ;
        RECT 393.555 -104.205 393.885 -103.875 ;
        RECT 393.555 -105.565 393.885 -105.235 ;
        RECT 393.555 -106.925 393.885 -106.595 ;
        RECT 393.555 -108.285 393.885 -107.955 ;
        RECT 393.555 -109.645 393.885 -109.315 ;
        RECT 393.555 -111.005 393.885 -110.675 ;
        RECT 393.555 -112.365 393.885 -112.035 ;
        RECT 393.555 -113.725 393.885 -113.395 ;
        RECT 393.555 -115.085 393.885 -114.755 ;
        RECT 393.555 -116.445 393.885 -116.115 ;
        RECT 393.555 -117.805 393.885 -117.475 ;
        RECT 393.555 -119.165 393.885 -118.835 ;
        RECT 393.555 -120.525 393.885 -120.195 ;
        RECT 393.555 -121.885 393.885 -121.555 ;
        RECT 393.555 -123.245 393.885 -122.915 ;
        RECT 393.555 -124.605 393.885 -124.275 ;
        RECT 393.555 -125.965 393.885 -125.635 ;
        RECT 393.555 -127.325 393.885 -126.995 ;
        RECT 393.555 -128.685 393.885 -128.355 ;
        RECT 393.555 -130.045 393.885 -129.715 ;
        RECT 393.555 -131.405 393.885 -131.075 ;
        RECT 393.555 -132.765 393.885 -132.435 ;
        RECT 393.555 -134.125 393.885 -133.795 ;
        RECT 393.555 -135.485 393.885 -135.155 ;
        RECT 393.555 -136.845 393.885 -136.515 ;
        RECT 393.555 -138.205 393.885 -137.875 ;
        RECT 393.555 -139.565 393.885 -139.235 ;
        RECT 393.555 -140.925 393.885 -140.595 ;
        RECT 393.555 -142.285 393.885 -141.955 ;
        RECT 393.555 -143.645 393.885 -143.315 ;
        RECT 393.555 -145.005 393.885 -144.675 ;
        RECT 393.555 -146.365 393.885 -146.035 ;
        RECT 393.555 -147.725 393.885 -147.395 ;
        RECT 393.555 -149.085 393.885 -148.755 ;
        RECT 393.555 -150.445 393.885 -150.115 ;
        RECT 393.555 -151.805 393.885 -151.475 ;
        RECT 393.555 -153.165 393.885 -152.835 ;
        RECT 393.555 -154.525 393.885 -154.195 ;
        RECT 393.555 -155.885 393.885 -155.555 ;
        RECT 393.555 -157.245 393.885 -156.915 ;
        RECT 393.555 -158.605 393.885 -158.275 ;
        RECT 393.555 -159.965 393.885 -159.635 ;
        RECT 393.555 -161.325 393.885 -160.995 ;
        RECT 393.555 -162.685 393.885 -162.355 ;
        RECT 393.555 -164.045 393.885 -163.715 ;
        RECT 393.555 -165.405 393.885 -165.075 ;
        RECT 393.555 -166.765 393.885 -166.435 ;
        RECT 393.555 -168.125 393.885 -167.795 ;
        RECT 393.555 -169.485 393.885 -169.155 ;
        RECT 393.555 -170.845 393.885 -170.515 ;
        RECT 393.555 -172.205 393.885 -171.875 ;
        RECT 393.555 -173.565 393.885 -173.235 ;
        RECT 393.555 -174.925 393.885 -174.595 ;
        RECT 393.555 -176.285 393.885 -175.955 ;
        RECT 393.555 -177.645 393.885 -177.315 ;
        RECT 393.555 -183.29 393.885 -182.16 ;
        RECT 393.56 -183.405 393.88 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 393.71 -94.075 394.04 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 394.915 244.04 395.245 245.17 ;
        RECT 394.915 239.875 395.245 240.205 ;
        RECT 394.915 238.515 395.245 238.845 ;
        RECT 394.915 237.155 395.245 237.485 ;
        RECT 394.92 237.155 395.24 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 394.915 -0.845 395.245 -0.515 ;
        RECT 394.915 -2.205 395.245 -1.875 ;
        RECT 394.915 -3.565 395.245 -3.235 ;
        RECT 394.92 -3.565 395.24 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 394.915 -91.965 395.245 -91.635 ;
        RECT 394.915 -93.325 395.245 -92.995 ;
        RECT 394.915 -94.685 395.245 -94.355 ;
        RECT 394.915 -96.045 395.245 -95.715 ;
        RECT 394.915 -97.405 395.245 -97.075 ;
        RECT 394.915 -98.765 395.245 -98.435 ;
        RECT 394.915 -100.125 395.245 -99.795 ;
        RECT 394.915 -101.485 395.245 -101.155 ;
        RECT 394.915 -102.845 395.245 -102.515 ;
        RECT 394.915 -104.205 395.245 -103.875 ;
        RECT 394.915 -105.565 395.245 -105.235 ;
        RECT 394.915 -106.925 395.245 -106.595 ;
        RECT 394.915 -108.285 395.245 -107.955 ;
        RECT 394.915 -109.645 395.245 -109.315 ;
        RECT 394.915 -111.005 395.245 -110.675 ;
        RECT 394.915 -112.365 395.245 -112.035 ;
        RECT 394.915 -113.725 395.245 -113.395 ;
        RECT 394.915 -115.085 395.245 -114.755 ;
        RECT 394.915 -116.445 395.245 -116.115 ;
        RECT 394.915 -117.805 395.245 -117.475 ;
        RECT 394.915 -119.165 395.245 -118.835 ;
        RECT 394.915 -120.525 395.245 -120.195 ;
        RECT 394.915 -121.885 395.245 -121.555 ;
        RECT 394.915 -123.245 395.245 -122.915 ;
        RECT 394.915 -124.605 395.245 -124.275 ;
        RECT 394.915 -125.965 395.245 -125.635 ;
        RECT 394.915 -127.325 395.245 -126.995 ;
        RECT 394.915 -128.685 395.245 -128.355 ;
        RECT 394.915 -130.045 395.245 -129.715 ;
        RECT 394.915 -131.405 395.245 -131.075 ;
        RECT 394.915 -132.765 395.245 -132.435 ;
        RECT 394.915 -134.125 395.245 -133.795 ;
        RECT 394.915 -135.485 395.245 -135.155 ;
        RECT 394.915 -136.845 395.245 -136.515 ;
        RECT 394.915 -138.205 395.245 -137.875 ;
        RECT 394.915 -139.565 395.245 -139.235 ;
        RECT 394.915 -140.925 395.245 -140.595 ;
        RECT 394.915 -142.285 395.245 -141.955 ;
        RECT 394.915 -143.645 395.245 -143.315 ;
        RECT 394.915 -145.005 395.245 -144.675 ;
        RECT 394.915 -146.365 395.245 -146.035 ;
        RECT 394.915 -147.725 395.245 -147.395 ;
        RECT 394.915 -149.085 395.245 -148.755 ;
        RECT 394.915 -150.445 395.245 -150.115 ;
        RECT 394.915 -151.805 395.245 -151.475 ;
        RECT 394.915 -153.165 395.245 -152.835 ;
        RECT 394.915 -154.525 395.245 -154.195 ;
        RECT 394.915 -155.885 395.245 -155.555 ;
        RECT 394.915 -157.245 395.245 -156.915 ;
        RECT 394.915 -158.605 395.245 -158.275 ;
        RECT 394.915 -159.965 395.245 -159.635 ;
        RECT 394.915 -161.325 395.245 -160.995 ;
        RECT 394.915 -162.685 395.245 -162.355 ;
        RECT 394.915 -164.045 395.245 -163.715 ;
        RECT 394.915 -165.405 395.245 -165.075 ;
        RECT 394.915 -166.765 395.245 -166.435 ;
        RECT 394.915 -168.125 395.245 -167.795 ;
        RECT 394.915 -169.485 395.245 -169.155 ;
        RECT 394.915 -170.845 395.245 -170.515 ;
        RECT 394.915 -172.205 395.245 -171.875 ;
        RECT 394.915 -173.565 395.245 -173.235 ;
        RECT 394.915 -174.925 395.245 -174.595 ;
        RECT 394.915 -176.285 395.245 -175.955 ;
        RECT 394.915 -177.645 395.245 -177.315 ;
        RECT 394.915 -183.29 395.245 -182.16 ;
        RECT 394.92 -183.405 395.24 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 396.275 244.04 396.605 245.17 ;
        RECT 396.275 239.875 396.605 240.205 ;
        RECT 396.275 238.515 396.605 238.845 ;
        RECT 396.275 237.155 396.605 237.485 ;
        RECT 396.28 237.155 396.6 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 396.275 -0.845 396.605 -0.515 ;
        RECT 396.275 -2.205 396.605 -1.875 ;
        RECT 396.275 -3.565 396.605 -3.235 ;
        RECT 396.28 -3.565 396.6 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 396.275 -91.965 396.605 -91.635 ;
        RECT 396.275 -93.325 396.605 -92.995 ;
        RECT 396.275 -94.685 396.605 -94.355 ;
        RECT 396.275 -96.045 396.605 -95.715 ;
        RECT 396.275 -97.405 396.605 -97.075 ;
        RECT 396.275 -98.765 396.605 -98.435 ;
        RECT 396.275 -100.125 396.605 -99.795 ;
        RECT 396.275 -101.485 396.605 -101.155 ;
        RECT 396.275 -102.845 396.605 -102.515 ;
        RECT 396.275 -104.205 396.605 -103.875 ;
        RECT 396.275 -105.565 396.605 -105.235 ;
        RECT 396.275 -106.925 396.605 -106.595 ;
        RECT 396.275 -108.285 396.605 -107.955 ;
        RECT 396.275 -109.645 396.605 -109.315 ;
        RECT 396.275 -111.005 396.605 -110.675 ;
        RECT 396.275 -112.365 396.605 -112.035 ;
        RECT 396.275 -113.725 396.605 -113.395 ;
        RECT 396.275 -115.085 396.605 -114.755 ;
        RECT 396.275 -116.445 396.605 -116.115 ;
        RECT 396.275 -117.805 396.605 -117.475 ;
        RECT 396.275 -119.165 396.605 -118.835 ;
        RECT 396.275 -120.525 396.605 -120.195 ;
        RECT 396.275 -121.885 396.605 -121.555 ;
        RECT 396.275 -123.245 396.605 -122.915 ;
        RECT 396.275 -124.605 396.605 -124.275 ;
        RECT 396.275 -125.965 396.605 -125.635 ;
        RECT 396.275 -127.325 396.605 -126.995 ;
        RECT 396.275 -128.685 396.605 -128.355 ;
        RECT 396.275 -130.045 396.605 -129.715 ;
        RECT 396.275 -131.405 396.605 -131.075 ;
        RECT 396.275 -132.765 396.605 -132.435 ;
        RECT 396.275 -134.125 396.605 -133.795 ;
        RECT 396.275 -135.485 396.605 -135.155 ;
        RECT 396.275 -136.845 396.605 -136.515 ;
        RECT 396.275 -138.205 396.605 -137.875 ;
        RECT 396.275 -139.565 396.605 -139.235 ;
        RECT 396.275 -140.925 396.605 -140.595 ;
        RECT 396.275 -142.285 396.605 -141.955 ;
        RECT 396.275 -143.645 396.605 -143.315 ;
        RECT 396.275 -145.005 396.605 -144.675 ;
        RECT 396.275 -146.365 396.605 -146.035 ;
        RECT 396.275 -147.725 396.605 -147.395 ;
        RECT 396.275 -149.085 396.605 -148.755 ;
        RECT 396.275 -150.445 396.605 -150.115 ;
        RECT 396.275 -151.805 396.605 -151.475 ;
        RECT 396.275 -153.165 396.605 -152.835 ;
        RECT 396.275 -154.525 396.605 -154.195 ;
        RECT 396.275 -155.885 396.605 -155.555 ;
        RECT 396.275 -157.245 396.605 -156.915 ;
        RECT 396.275 -158.605 396.605 -158.275 ;
        RECT 396.275 -159.965 396.605 -159.635 ;
        RECT 396.275 -161.325 396.605 -160.995 ;
        RECT 396.275 -162.685 396.605 -162.355 ;
        RECT 396.275 -164.045 396.605 -163.715 ;
        RECT 396.275 -165.405 396.605 -165.075 ;
        RECT 396.275 -166.765 396.605 -166.435 ;
        RECT 396.275 -168.125 396.605 -167.795 ;
        RECT 396.275 -169.485 396.605 -169.155 ;
        RECT 396.275 -170.845 396.605 -170.515 ;
        RECT 396.275 -172.205 396.605 -171.875 ;
        RECT 396.275 -173.565 396.605 -173.235 ;
        RECT 396.275 -174.925 396.605 -174.595 ;
        RECT 396.275 -176.285 396.605 -175.955 ;
        RECT 396.275 -177.645 396.605 -177.315 ;
        RECT 396.275 -183.29 396.605 -182.16 ;
        RECT 396.28 -183.405 396.6 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 397.635 17.265 397.965 17.595 ;
        RECT 397.635 14.955 397.965 15.285 ;
        RECT 397.635 14.105 397.965 14.435 ;
        RECT 397.635 11.795 397.965 12.125 ;
        RECT 397.635 10.945 397.965 11.275 ;
        RECT 397.635 8.635 397.965 8.965 ;
        RECT 397.635 7.785 397.965 8.115 ;
        RECT 397.635 5.475 397.965 5.805 ;
        RECT 397.635 3.895 397.965 4.225 ;
        RECT 397.635 3.045 397.965 3.375 ;
        RECT 397.635 0.87 397.965 1.2 ;
        RECT 397.635 -0.845 397.965 -0.515 ;
        RECT 397.635 -2.205 397.965 -1.875 ;
        RECT 397.635 -3.565 397.965 -3.235 ;
        RECT 397.635 -4.925 397.965 -4.595 ;
        RECT 397.635 -6.285 397.965 -5.955 ;
        RECT 397.635 -7.645 397.965 -7.315 ;
        RECT 397.635 -9.005 397.965 -8.675 ;
        RECT 397.635 -10.365 397.965 -10.035 ;
        RECT 397.635 -11.725 397.965 -11.395 ;
        RECT 397.635 -13.085 397.965 -12.755 ;
        RECT 397.635 -14.445 397.965 -14.115 ;
        RECT 397.635 -15.805 397.965 -15.475 ;
        RECT 397.635 -17.165 397.965 -16.835 ;
        RECT 397.635 -18.525 397.965 -18.195 ;
        RECT 397.635 -19.885 397.965 -19.555 ;
        RECT 397.635 -21.245 397.965 -20.915 ;
        RECT 397.635 -22.605 397.965 -22.275 ;
        RECT 397.635 -23.965 397.965 -23.635 ;
        RECT 397.635 -25.325 397.965 -24.995 ;
        RECT 397.635 -26.685 397.965 -26.355 ;
        RECT 397.635 -28.045 397.965 -27.715 ;
        RECT 397.635 -29.405 397.965 -29.075 ;
        RECT 397.635 -30.765 397.965 -30.435 ;
        RECT 397.635 -32.125 397.965 -31.795 ;
        RECT 397.635 -33.485 397.965 -33.155 ;
        RECT 397.635 -34.845 397.965 -34.515 ;
        RECT 397.635 -36.205 397.965 -35.875 ;
        RECT 397.635 -37.565 397.965 -37.235 ;
        RECT 397.635 -38.925 397.965 -38.595 ;
        RECT 397.635 -40.285 397.965 -39.955 ;
        RECT 397.635 -41.645 397.965 -41.315 ;
        RECT 397.635 -43.005 397.965 -42.675 ;
        RECT 397.635 -44.365 397.965 -44.035 ;
        RECT 397.635 -45.725 397.965 -45.395 ;
        RECT 397.635 -47.085 397.965 -46.755 ;
        RECT 397.635 -48.445 397.965 -48.115 ;
        RECT 397.635 -49.805 397.965 -49.475 ;
        RECT 397.635 -51.165 397.965 -50.835 ;
        RECT 397.635 -52.525 397.965 -52.195 ;
        RECT 397.635 -53.885 397.965 -53.555 ;
        RECT 397.635 -55.245 397.965 -54.915 ;
        RECT 397.635 -56.605 397.965 -56.275 ;
        RECT 397.635 -57.965 397.965 -57.635 ;
        RECT 397.635 -59.325 397.965 -58.995 ;
        RECT 397.635 -60.685 397.965 -60.355 ;
        RECT 397.635 -62.045 397.965 -61.715 ;
        RECT 397.635 -63.405 397.965 -63.075 ;
        RECT 397.635 -64.765 397.965 -64.435 ;
        RECT 397.635 -66.125 397.965 -65.795 ;
        RECT 397.635 -67.485 397.965 -67.155 ;
        RECT 397.635 -68.845 397.965 -68.515 ;
        RECT 397.635 -70.205 397.965 -69.875 ;
        RECT 397.635 -71.565 397.965 -71.235 ;
        RECT 397.635 -72.925 397.965 -72.595 ;
        RECT 397.635 -74.285 397.965 -73.955 ;
        RECT 397.635 -75.645 397.965 -75.315 ;
        RECT 397.635 -77.005 397.965 -76.675 ;
        RECT 397.635 -78.365 397.965 -78.035 ;
        RECT 397.635 -79.725 397.965 -79.395 ;
        RECT 397.635 -81.085 397.965 -80.755 ;
        RECT 397.635 -82.445 397.965 -82.115 ;
        RECT 397.635 -83.805 397.965 -83.475 ;
        RECT 397.635 -85.165 397.965 -84.835 ;
        RECT 397.635 -86.525 397.965 -86.195 ;
        RECT 397.635 -87.885 397.965 -87.555 ;
        RECT 397.635 -89.245 397.965 -88.915 ;
        RECT 397.635 -90.605 397.965 -90.275 ;
        RECT 397.635 -91.965 397.965 -91.635 ;
        RECT 397.635 -93.325 397.965 -92.995 ;
        RECT 397.635 -94.685 397.965 -94.355 ;
        RECT 397.635 -96.045 397.965 -95.715 ;
        RECT 397.635 -97.405 397.965 -97.075 ;
        RECT 397.635 -98.765 397.965 -98.435 ;
        RECT 397.635 -100.125 397.965 -99.795 ;
        RECT 397.635 -101.485 397.965 -101.155 ;
        RECT 397.635 -102.845 397.965 -102.515 ;
        RECT 397.635 -104.205 397.965 -103.875 ;
        RECT 397.635 -105.565 397.965 -105.235 ;
        RECT 397.635 -106.925 397.965 -106.595 ;
        RECT 397.635 -108.285 397.965 -107.955 ;
        RECT 397.635 -109.645 397.965 -109.315 ;
        RECT 397.635 -111.005 397.965 -110.675 ;
        RECT 397.635 -112.365 397.965 -112.035 ;
        RECT 397.635 -113.725 397.965 -113.395 ;
        RECT 397.635 -115.085 397.965 -114.755 ;
        RECT 397.635 -116.445 397.965 -116.115 ;
        RECT 397.635 -117.805 397.965 -117.475 ;
        RECT 397.635 -119.165 397.965 -118.835 ;
        RECT 397.635 -120.525 397.965 -120.195 ;
        RECT 397.635 -121.885 397.965 -121.555 ;
        RECT 397.635 -123.245 397.965 -122.915 ;
        RECT 397.635 -124.605 397.965 -124.275 ;
        RECT 397.635 -125.965 397.965 -125.635 ;
        RECT 397.635 -127.325 397.965 -126.995 ;
        RECT 397.635 -128.685 397.965 -128.355 ;
        RECT 397.635 -130.045 397.965 -129.715 ;
        RECT 397.635 -131.405 397.965 -131.075 ;
        RECT 397.635 -132.765 397.965 -132.435 ;
        RECT 397.635 -134.125 397.965 -133.795 ;
        RECT 397.635 -135.485 397.965 -135.155 ;
        RECT 397.635 -136.845 397.965 -136.515 ;
        RECT 397.635 -138.205 397.965 -137.875 ;
        RECT 397.635 -139.565 397.965 -139.235 ;
        RECT 397.635 -140.925 397.965 -140.595 ;
        RECT 397.635 -142.285 397.965 -141.955 ;
        RECT 397.635 -143.645 397.965 -143.315 ;
        RECT 397.635 -145.005 397.965 -144.675 ;
        RECT 397.635 -146.365 397.965 -146.035 ;
        RECT 397.635 -147.725 397.965 -147.395 ;
        RECT 397.635 -149.085 397.965 -148.755 ;
        RECT 397.635 -150.445 397.965 -150.115 ;
        RECT 397.635 -151.805 397.965 -151.475 ;
        RECT 397.635 -153.165 397.965 -152.835 ;
        RECT 397.635 -154.525 397.965 -154.195 ;
        RECT 397.635 -155.885 397.965 -155.555 ;
        RECT 397.635 -157.245 397.965 -156.915 ;
        RECT 397.635 -158.605 397.965 -158.275 ;
        RECT 397.635 -159.965 397.965 -159.635 ;
        RECT 397.635 -161.325 397.965 -160.995 ;
        RECT 397.635 -162.685 397.965 -162.355 ;
        RECT 397.635 -164.045 397.965 -163.715 ;
        RECT 397.635 -165.405 397.965 -165.075 ;
        RECT 397.635 -166.765 397.965 -166.435 ;
        RECT 397.635 -168.125 397.965 -167.795 ;
        RECT 397.635 -169.485 397.965 -169.155 ;
        RECT 397.635 -170.845 397.965 -170.515 ;
        RECT 397.635 -172.205 397.965 -171.875 ;
        RECT 397.635 -173.565 397.965 -173.235 ;
        RECT 397.635 -174.925 397.965 -174.595 ;
        RECT 397.635 -176.285 397.965 -175.955 ;
        RECT 397.635 -177.645 397.965 -177.315 ;
        RECT 397.635 -183.29 397.965 -182.16 ;
        RECT 397.64 -183.405 397.96 245.285 ;
        RECT 397.635 244.04 397.965 245.17 ;
        RECT 397.635 239.875 397.965 240.205 ;
        RECT 397.635 238.515 397.965 238.845 ;
        RECT 397.635 237.155 397.965 237.485 ;
        RECT 397.635 235.17 397.965 235.5 ;
        RECT 397.635 232.995 397.965 233.325 ;
        RECT 397.635 231.415 397.965 231.745 ;
        RECT 397.635 230.565 397.965 230.895 ;
        RECT 397.635 228.255 397.965 228.585 ;
        RECT 397.635 227.405 397.965 227.735 ;
        RECT 397.635 225.095 397.965 225.425 ;
        RECT 397.635 224.245 397.965 224.575 ;
        RECT 397.635 221.935 397.965 222.265 ;
        RECT 397.635 221.085 397.965 221.415 ;
        RECT 397.635 218.775 397.965 219.105 ;
        RECT 397.635 217.195 397.965 217.525 ;
        RECT 397.635 216.345 397.965 216.675 ;
        RECT 397.635 214.035 397.965 214.365 ;
        RECT 397.635 213.185 397.965 213.515 ;
        RECT 397.635 210.875 397.965 211.205 ;
        RECT 397.635 210.025 397.965 210.355 ;
        RECT 397.635 207.715 397.965 208.045 ;
        RECT 397.635 206.865 397.965 207.195 ;
        RECT 397.635 204.555 397.965 204.885 ;
        RECT 397.635 202.975 397.965 203.305 ;
        RECT 397.635 202.125 397.965 202.455 ;
        RECT 397.635 199.815 397.965 200.145 ;
        RECT 397.635 198.965 397.965 199.295 ;
        RECT 397.635 196.655 397.965 196.985 ;
        RECT 397.635 195.805 397.965 196.135 ;
        RECT 397.635 193.495 397.965 193.825 ;
        RECT 397.635 192.645 397.965 192.975 ;
        RECT 397.635 190.335 397.965 190.665 ;
        RECT 397.635 188.755 397.965 189.085 ;
        RECT 397.635 187.905 397.965 188.235 ;
        RECT 397.635 185.595 397.965 185.925 ;
        RECT 397.635 184.745 397.965 185.075 ;
        RECT 397.635 182.435 397.965 182.765 ;
        RECT 397.635 181.585 397.965 181.915 ;
        RECT 397.635 179.275 397.965 179.605 ;
        RECT 397.635 178.425 397.965 178.755 ;
        RECT 397.635 176.115 397.965 176.445 ;
        RECT 397.635 174.535 397.965 174.865 ;
        RECT 397.635 173.685 397.965 174.015 ;
        RECT 397.635 171.375 397.965 171.705 ;
        RECT 397.635 170.525 397.965 170.855 ;
        RECT 397.635 168.215 397.965 168.545 ;
        RECT 397.635 167.365 397.965 167.695 ;
        RECT 397.635 165.055 397.965 165.385 ;
        RECT 397.635 164.205 397.965 164.535 ;
        RECT 397.635 161.895 397.965 162.225 ;
        RECT 397.635 160.315 397.965 160.645 ;
        RECT 397.635 159.465 397.965 159.795 ;
        RECT 397.635 157.155 397.965 157.485 ;
        RECT 397.635 156.305 397.965 156.635 ;
        RECT 397.635 153.995 397.965 154.325 ;
        RECT 397.635 153.145 397.965 153.475 ;
        RECT 397.635 150.835 397.965 151.165 ;
        RECT 397.635 149.985 397.965 150.315 ;
        RECT 397.635 147.675 397.965 148.005 ;
        RECT 397.635 146.095 397.965 146.425 ;
        RECT 397.635 145.245 397.965 145.575 ;
        RECT 397.635 142.935 397.965 143.265 ;
        RECT 397.635 142.085 397.965 142.415 ;
        RECT 397.635 139.775 397.965 140.105 ;
        RECT 397.635 138.925 397.965 139.255 ;
        RECT 397.635 136.615 397.965 136.945 ;
        RECT 397.635 135.765 397.965 136.095 ;
        RECT 397.635 133.455 397.965 133.785 ;
        RECT 397.635 131.875 397.965 132.205 ;
        RECT 397.635 131.025 397.965 131.355 ;
        RECT 397.635 128.715 397.965 129.045 ;
        RECT 397.635 127.865 397.965 128.195 ;
        RECT 397.635 125.555 397.965 125.885 ;
        RECT 397.635 124.705 397.965 125.035 ;
        RECT 397.635 122.395 397.965 122.725 ;
        RECT 397.635 121.545 397.965 121.875 ;
        RECT 397.635 119.235 397.965 119.565 ;
        RECT 397.635 117.655 397.965 117.985 ;
        RECT 397.635 116.805 397.965 117.135 ;
        RECT 397.635 114.495 397.965 114.825 ;
        RECT 397.635 113.645 397.965 113.975 ;
        RECT 397.635 111.335 397.965 111.665 ;
        RECT 397.635 110.485 397.965 110.815 ;
        RECT 397.635 108.175 397.965 108.505 ;
        RECT 397.635 107.325 397.965 107.655 ;
        RECT 397.635 105.015 397.965 105.345 ;
        RECT 397.635 103.435 397.965 103.765 ;
        RECT 397.635 102.585 397.965 102.915 ;
        RECT 397.635 100.275 397.965 100.605 ;
        RECT 397.635 99.425 397.965 99.755 ;
        RECT 397.635 97.115 397.965 97.445 ;
        RECT 397.635 96.265 397.965 96.595 ;
        RECT 397.635 93.955 397.965 94.285 ;
        RECT 397.635 93.105 397.965 93.435 ;
        RECT 397.635 90.795 397.965 91.125 ;
        RECT 397.635 89.215 397.965 89.545 ;
        RECT 397.635 88.365 397.965 88.695 ;
        RECT 397.635 86.055 397.965 86.385 ;
        RECT 397.635 85.205 397.965 85.535 ;
        RECT 397.635 82.895 397.965 83.225 ;
        RECT 397.635 82.045 397.965 82.375 ;
        RECT 397.635 79.735 397.965 80.065 ;
        RECT 397.635 78.885 397.965 79.215 ;
        RECT 397.635 76.575 397.965 76.905 ;
        RECT 397.635 74.995 397.965 75.325 ;
        RECT 397.635 74.145 397.965 74.475 ;
        RECT 397.635 71.835 397.965 72.165 ;
        RECT 397.635 70.985 397.965 71.315 ;
        RECT 397.635 68.675 397.965 69.005 ;
        RECT 397.635 67.825 397.965 68.155 ;
        RECT 397.635 65.515 397.965 65.845 ;
        RECT 397.635 64.665 397.965 64.995 ;
        RECT 397.635 62.355 397.965 62.685 ;
        RECT 397.635 60.775 397.965 61.105 ;
        RECT 397.635 59.925 397.965 60.255 ;
        RECT 397.635 57.615 397.965 57.945 ;
        RECT 397.635 56.765 397.965 57.095 ;
        RECT 397.635 54.455 397.965 54.785 ;
        RECT 397.635 53.605 397.965 53.935 ;
        RECT 397.635 51.295 397.965 51.625 ;
        RECT 397.635 50.445 397.965 50.775 ;
        RECT 397.635 48.135 397.965 48.465 ;
        RECT 397.635 46.555 397.965 46.885 ;
        RECT 397.635 45.705 397.965 46.035 ;
        RECT 397.635 43.395 397.965 43.725 ;
        RECT 397.635 42.545 397.965 42.875 ;
        RECT 397.635 40.235 397.965 40.565 ;
        RECT 397.635 39.385 397.965 39.715 ;
        RECT 397.635 37.075 397.965 37.405 ;
        RECT 397.635 36.225 397.965 36.555 ;
        RECT 397.635 33.915 397.965 34.245 ;
        RECT 397.635 32.335 397.965 32.665 ;
        RECT 397.635 31.485 397.965 31.815 ;
        RECT 397.635 29.175 397.965 29.505 ;
        RECT 397.635 28.325 397.965 28.655 ;
        RECT 397.635 26.015 397.965 26.345 ;
        RECT 397.635 25.165 397.965 25.495 ;
        RECT 397.635 22.855 397.965 23.185 ;
        RECT 397.635 22.005 397.965 22.335 ;
        RECT 397.635 19.695 397.965 20.025 ;
        RECT 397.635 18.115 397.965 18.445 ;
    END
    PORT
      LAYER met3 ;
        RECT 343.235 244.04 343.565 245.17 ;
        RECT 343.235 239.875 343.565 240.205 ;
        RECT 343.235 238.515 343.565 238.845 ;
        RECT 343.235 237.155 343.565 237.485 ;
        RECT 343.24 237.155 343.56 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 343.235 -0.845 343.565 -0.515 ;
        RECT 343.235 -2.205 343.565 -1.875 ;
        RECT 343.235 -3.565 343.565 -3.235 ;
        RECT 343.24 -3.565 343.56 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 343.235 -91.965 343.565 -91.635 ;
        RECT 343.235 -93.325 343.565 -92.995 ;
        RECT 343.235 -94.685 343.565 -94.355 ;
        RECT 343.235 -96.045 343.565 -95.715 ;
        RECT 343.235 -97.405 343.565 -97.075 ;
        RECT 343.235 -98.765 343.565 -98.435 ;
        RECT 343.235 -100.125 343.565 -99.795 ;
        RECT 343.235 -101.485 343.565 -101.155 ;
        RECT 343.235 -102.845 343.565 -102.515 ;
        RECT 343.235 -104.205 343.565 -103.875 ;
        RECT 343.235 -105.565 343.565 -105.235 ;
        RECT 343.235 -106.925 343.565 -106.595 ;
        RECT 343.235 -108.285 343.565 -107.955 ;
        RECT 343.235 -109.645 343.565 -109.315 ;
        RECT 343.235 -111.005 343.565 -110.675 ;
        RECT 343.235 -112.365 343.565 -112.035 ;
        RECT 343.235 -113.725 343.565 -113.395 ;
        RECT 343.235 -115.085 343.565 -114.755 ;
        RECT 343.235 -116.445 343.565 -116.115 ;
        RECT 343.235 -117.805 343.565 -117.475 ;
        RECT 343.235 -119.165 343.565 -118.835 ;
        RECT 343.235 -120.525 343.565 -120.195 ;
        RECT 343.235 -121.885 343.565 -121.555 ;
        RECT 343.235 -123.245 343.565 -122.915 ;
        RECT 343.235 -124.605 343.565 -124.275 ;
        RECT 343.235 -125.965 343.565 -125.635 ;
        RECT 343.235 -127.325 343.565 -126.995 ;
        RECT 343.235 -128.685 343.565 -128.355 ;
        RECT 343.235 -130.045 343.565 -129.715 ;
        RECT 343.235 -131.405 343.565 -131.075 ;
        RECT 343.235 -132.765 343.565 -132.435 ;
        RECT 343.235 -134.125 343.565 -133.795 ;
        RECT 343.235 -135.485 343.565 -135.155 ;
        RECT 343.235 -136.845 343.565 -136.515 ;
        RECT 343.235 -138.205 343.565 -137.875 ;
        RECT 343.235 -139.565 343.565 -139.235 ;
        RECT 343.235 -140.925 343.565 -140.595 ;
        RECT 343.235 -142.285 343.565 -141.955 ;
        RECT 343.235 -143.645 343.565 -143.315 ;
        RECT 343.235 -145.005 343.565 -144.675 ;
        RECT 343.235 -146.365 343.565 -146.035 ;
        RECT 343.235 -147.725 343.565 -147.395 ;
        RECT 343.235 -149.085 343.565 -148.755 ;
        RECT 343.235 -150.445 343.565 -150.115 ;
        RECT 343.235 -151.805 343.565 -151.475 ;
        RECT 343.235 -153.165 343.565 -152.835 ;
        RECT 343.235 -154.525 343.565 -154.195 ;
        RECT 343.235 -155.885 343.565 -155.555 ;
        RECT 343.235 -157.245 343.565 -156.915 ;
        RECT 343.235 -158.605 343.565 -158.275 ;
        RECT 343.235 -159.965 343.565 -159.635 ;
        RECT 343.235 -161.325 343.565 -160.995 ;
        RECT 343.235 -162.685 343.565 -162.355 ;
        RECT 343.235 -164.045 343.565 -163.715 ;
        RECT 343.235 -165.405 343.565 -165.075 ;
        RECT 343.235 -166.765 343.565 -166.435 ;
        RECT 343.235 -168.125 343.565 -167.795 ;
        RECT 343.235 -169.485 343.565 -169.155 ;
        RECT 343.235 -170.845 343.565 -170.515 ;
        RECT 343.235 -172.205 343.565 -171.875 ;
        RECT 343.235 -173.565 343.565 -173.235 ;
        RECT 343.235 -174.925 343.565 -174.595 ;
        RECT 343.235 -176.285 343.565 -175.955 ;
        RECT 343.235 -177.645 343.565 -177.315 ;
        RECT 343.235 -183.29 343.565 -182.16 ;
        RECT 343.24 -183.405 343.56 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 344.26 -94.075 344.59 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 344.595 244.04 344.925 245.17 ;
        RECT 344.595 239.875 344.925 240.205 ;
        RECT 344.595 238.515 344.925 238.845 ;
        RECT 344.595 237.155 344.925 237.485 ;
        RECT 344.6 237.155 344.92 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 344.595 -96.045 344.925 -95.715 ;
        RECT 344.595 -97.405 344.925 -97.075 ;
        RECT 344.595 -98.765 344.925 -98.435 ;
        RECT 344.595 -100.125 344.925 -99.795 ;
        RECT 344.595 -101.485 344.925 -101.155 ;
        RECT 344.595 -102.845 344.925 -102.515 ;
        RECT 344.595 -104.205 344.925 -103.875 ;
        RECT 344.595 -105.565 344.925 -105.235 ;
        RECT 344.595 -106.925 344.925 -106.595 ;
        RECT 344.595 -108.285 344.925 -107.955 ;
        RECT 344.595 -109.645 344.925 -109.315 ;
        RECT 344.595 -111.005 344.925 -110.675 ;
        RECT 344.595 -112.365 344.925 -112.035 ;
        RECT 344.595 -113.725 344.925 -113.395 ;
        RECT 344.595 -115.085 344.925 -114.755 ;
        RECT 344.595 -116.445 344.925 -116.115 ;
        RECT 344.595 -117.805 344.925 -117.475 ;
        RECT 344.595 -119.165 344.925 -118.835 ;
        RECT 344.595 -120.525 344.925 -120.195 ;
        RECT 344.595 -121.885 344.925 -121.555 ;
        RECT 344.595 -123.245 344.925 -122.915 ;
        RECT 344.595 -124.605 344.925 -124.275 ;
        RECT 344.595 -125.965 344.925 -125.635 ;
        RECT 344.595 -127.325 344.925 -126.995 ;
        RECT 344.595 -128.685 344.925 -128.355 ;
        RECT 344.595 -130.045 344.925 -129.715 ;
        RECT 344.595 -131.405 344.925 -131.075 ;
        RECT 344.595 -132.765 344.925 -132.435 ;
        RECT 344.595 -134.125 344.925 -133.795 ;
        RECT 344.595 -135.485 344.925 -135.155 ;
        RECT 344.595 -136.845 344.925 -136.515 ;
        RECT 344.595 -138.205 344.925 -137.875 ;
        RECT 344.595 -139.565 344.925 -139.235 ;
        RECT 344.595 -140.925 344.925 -140.595 ;
        RECT 344.595 -142.285 344.925 -141.955 ;
        RECT 344.595 -143.645 344.925 -143.315 ;
        RECT 344.595 -145.005 344.925 -144.675 ;
        RECT 344.595 -146.365 344.925 -146.035 ;
        RECT 344.595 -147.725 344.925 -147.395 ;
        RECT 344.595 -149.085 344.925 -148.755 ;
        RECT 344.595 -150.445 344.925 -150.115 ;
        RECT 344.595 -151.805 344.925 -151.475 ;
        RECT 344.595 -153.165 344.925 -152.835 ;
        RECT 344.595 -154.525 344.925 -154.195 ;
        RECT 344.595 -155.885 344.925 -155.555 ;
        RECT 344.595 -157.245 344.925 -156.915 ;
        RECT 344.595 -158.605 344.925 -158.275 ;
        RECT 344.595 -159.965 344.925 -159.635 ;
        RECT 344.595 -161.325 344.925 -160.995 ;
        RECT 344.595 -162.685 344.925 -162.355 ;
        RECT 344.595 -164.045 344.925 -163.715 ;
        RECT 344.595 -165.405 344.925 -165.075 ;
        RECT 344.595 -166.765 344.925 -166.435 ;
        RECT 344.595 -168.125 344.925 -167.795 ;
        RECT 344.595 -169.485 344.925 -169.155 ;
        RECT 344.595 -170.845 344.925 -170.515 ;
        RECT 344.595 -172.205 344.925 -171.875 ;
        RECT 344.595 -173.565 344.925 -173.235 ;
        RECT 344.595 -174.925 344.925 -174.595 ;
        RECT 344.595 -176.285 344.925 -175.955 ;
        RECT 344.595 -177.645 344.925 -177.315 ;
        RECT 344.595 -183.29 344.925 -182.16 ;
        RECT 344.6 -183.405 344.92 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 345.955 244.04 346.285 245.17 ;
        RECT 345.955 239.875 346.285 240.205 ;
        RECT 345.955 238.515 346.285 238.845 ;
        RECT 345.955 237.155 346.285 237.485 ;
        RECT 345.96 237.155 346.28 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 345.955 -0.845 346.285 -0.515 ;
        RECT 345.955 -2.205 346.285 -1.875 ;
        RECT 345.955 -3.565 346.285 -3.235 ;
        RECT 345.96 -3.565 346.28 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 347.315 244.04 347.645 245.17 ;
        RECT 347.315 239.875 347.645 240.205 ;
        RECT 347.315 238.515 347.645 238.845 ;
        RECT 347.315 237.155 347.645 237.485 ;
        RECT 347.32 237.155 347.64 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 347.315 -0.845 347.645 -0.515 ;
        RECT 347.315 -2.205 347.645 -1.875 ;
        RECT 347.315 -3.565 347.645 -3.235 ;
        RECT 347.32 -3.565 347.64 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 348.675 244.04 349.005 245.17 ;
        RECT 348.675 239.875 349.005 240.205 ;
        RECT 348.675 238.515 349.005 238.845 ;
        RECT 348.675 237.155 349.005 237.485 ;
        RECT 348.68 237.155 349 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 348.675 -0.845 349.005 -0.515 ;
        RECT 348.675 -2.205 349.005 -1.875 ;
        RECT 348.675 -3.565 349.005 -3.235 ;
        RECT 348.68 -3.565 349 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 350.035 244.04 350.365 245.17 ;
        RECT 350.035 239.875 350.365 240.205 ;
        RECT 350.035 238.515 350.365 238.845 ;
        RECT 350.035 237.155 350.365 237.485 ;
        RECT 350.04 237.155 350.36 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 350.035 -96.045 350.365 -95.715 ;
        RECT 350.035 -97.405 350.365 -97.075 ;
        RECT 350.035 -98.765 350.365 -98.435 ;
        RECT 350.035 -100.125 350.365 -99.795 ;
        RECT 350.035 -101.485 350.365 -101.155 ;
        RECT 350.035 -102.845 350.365 -102.515 ;
        RECT 350.035 -104.205 350.365 -103.875 ;
        RECT 350.035 -105.565 350.365 -105.235 ;
        RECT 350.035 -106.925 350.365 -106.595 ;
        RECT 350.035 -108.285 350.365 -107.955 ;
        RECT 350.035 -109.645 350.365 -109.315 ;
        RECT 350.035 -111.005 350.365 -110.675 ;
        RECT 350.035 -112.365 350.365 -112.035 ;
        RECT 350.035 -113.725 350.365 -113.395 ;
        RECT 350.035 -115.085 350.365 -114.755 ;
        RECT 350.035 -116.445 350.365 -116.115 ;
        RECT 350.035 -117.805 350.365 -117.475 ;
        RECT 350.035 -119.165 350.365 -118.835 ;
        RECT 350.035 -120.525 350.365 -120.195 ;
        RECT 350.035 -121.885 350.365 -121.555 ;
        RECT 350.035 -123.245 350.365 -122.915 ;
        RECT 350.035 -124.605 350.365 -124.275 ;
        RECT 350.035 -125.965 350.365 -125.635 ;
        RECT 350.035 -127.325 350.365 -126.995 ;
        RECT 350.035 -128.685 350.365 -128.355 ;
        RECT 350.035 -130.045 350.365 -129.715 ;
        RECT 350.035 -131.405 350.365 -131.075 ;
        RECT 350.035 -132.765 350.365 -132.435 ;
        RECT 350.035 -134.125 350.365 -133.795 ;
        RECT 350.035 -135.485 350.365 -135.155 ;
        RECT 350.035 -136.845 350.365 -136.515 ;
        RECT 350.035 -138.205 350.365 -137.875 ;
        RECT 350.035 -139.565 350.365 -139.235 ;
        RECT 350.035 -140.925 350.365 -140.595 ;
        RECT 350.035 -142.285 350.365 -141.955 ;
        RECT 350.035 -143.645 350.365 -143.315 ;
        RECT 350.035 -145.005 350.365 -144.675 ;
        RECT 350.035 -146.365 350.365 -146.035 ;
        RECT 350.035 -147.725 350.365 -147.395 ;
        RECT 350.035 -149.085 350.365 -148.755 ;
        RECT 350.035 -150.445 350.365 -150.115 ;
        RECT 350.035 -151.805 350.365 -151.475 ;
        RECT 350.035 -153.165 350.365 -152.835 ;
        RECT 350.035 -154.525 350.365 -154.195 ;
        RECT 350.035 -155.885 350.365 -155.555 ;
        RECT 350.035 -157.245 350.365 -156.915 ;
        RECT 350.035 -158.605 350.365 -158.275 ;
        RECT 350.035 -159.965 350.365 -159.635 ;
        RECT 350.035 -161.325 350.365 -160.995 ;
        RECT 350.035 -162.685 350.365 -162.355 ;
        RECT 350.035 -164.045 350.365 -163.715 ;
        RECT 350.035 -165.405 350.365 -165.075 ;
        RECT 350.035 -166.765 350.365 -166.435 ;
        RECT 350.035 -168.125 350.365 -167.795 ;
        RECT 350.035 -169.485 350.365 -169.155 ;
        RECT 350.035 -170.845 350.365 -170.515 ;
        RECT 350.035 -172.205 350.365 -171.875 ;
        RECT 350.035 -173.565 350.365 -173.235 ;
        RECT 350.035 -174.925 350.365 -174.595 ;
        RECT 350.035 -176.285 350.365 -175.955 ;
        RECT 350.035 -177.645 350.365 -177.315 ;
        RECT 350.035 -183.29 350.365 -182.16 ;
        RECT 350.04 -183.405 350.36 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 350.36 -94.075 350.69 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 351.395 244.04 351.725 245.17 ;
        RECT 351.395 239.875 351.725 240.205 ;
        RECT 351.395 238.515 351.725 238.845 ;
        RECT 351.395 237.155 351.725 237.485 ;
        RECT 351.4 237.155 351.72 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 352.755 244.04 353.085 245.17 ;
        RECT 352.755 239.875 353.085 240.205 ;
        RECT 352.755 238.515 353.085 238.845 ;
        RECT 352.755 237.155 353.085 237.485 ;
        RECT 352.76 237.155 353.08 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 352.755 -0.845 353.085 -0.515 ;
        RECT 352.755 -2.205 353.085 -1.875 ;
        RECT 352.755 -3.565 353.085 -3.235 ;
        RECT 352.76 -3.565 353.08 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 354.115 244.04 354.445 245.17 ;
        RECT 354.115 239.875 354.445 240.205 ;
        RECT 354.115 238.515 354.445 238.845 ;
        RECT 354.115 237.155 354.445 237.485 ;
        RECT 354.12 237.155 354.44 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 354.115 -0.845 354.445 -0.515 ;
        RECT 354.115 -2.205 354.445 -1.875 ;
        RECT 354.115 -3.565 354.445 -3.235 ;
        RECT 354.12 -3.565 354.44 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 354.115 -91.965 354.445 -91.635 ;
        RECT 354.115 -93.325 354.445 -92.995 ;
        RECT 354.115 -94.685 354.445 -94.355 ;
        RECT 354.115 -96.045 354.445 -95.715 ;
        RECT 354.115 -97.405 354.445 -97.075 ;
        RECT 354.115 -98.765 354.445 -98.435 ;
        RECT 354.115 -100.125 354.445 -99.795 ;
        RECT 354.115 -101.485 354.445 -101.155 ;
        RECT 354.115 -102.845 354.445 -102.515 ;
        RECT 354.115 -104.205 354.445 -103.875 ;
        RECT 354.115 -105.565 354.445 -105.235 ;
        RECT 354.115 -106.925 354.445 -106.595 ;
        RECT 354.115 -108.285 354.445 -107.955 ;
        RECT 354.115 -109.645 354.445 -109.315 ;
        RECT 354.115 -111.005 354.445 -110.675 ;
        RECT 354.115 -112.365 354.445 -112.035 ;
        RECT 354.115 -113.725 354.445 -113.395 ;
        RECT 354.115 -115.085 354.445 -114.755 ;
        RECT 354.115 -116.445 354.445 -116.115 ;
        RECT 354.115 -117.805 354.445 -117.475 ;
        RECT 354.115 -119.165 354.445 -118.835 ;
        RECT 354.115 -120.525 354.445 -120.195 ;
        RECT 354.115 -121.885 354.445 -121.555 ;
        RECT 354.115 -123.245 354.445 -122.915 ;
        RECT 354.115 -124.605 354.445 -124.275 ;
        RECT 354.115 -125.965 354.445 -125.635 ;
        RECT 354.115 -127.325 354.445 -126.995 ;
        RECT 354.115 -128.685 354.445 -128.355 ;
        RECT 354.115 -130.045 354.445 -129.715 ;
        RECT 354.115 -131.405 354.445 -131.075 ;
        RECT 354.115 -132.765 354.445 -132.435 ;
        RECT 354.115 -134.125 354.445 -133.795 ;
        RECT 354.115 -135.485 354.445 -135.155 ;
        RECT 354.115 -136.845 354.445 -136.515 ;
        RECT 354.115 -138.205 354.445 -137.875 ;
        RECT 354.115 -139.565 354.445 -139.235 ;
        RECT 354.115 -140.925 354.445 -140.595 ;
        RECT 354.115 -142.285 354.445 -141.955 ;
        RECT 354.115 -143.645 354.445 -143.315 ;
        RECT 354.115 -145.005 354.445 -144.675 ;
        RECT 354.115 -146.365 354.445 -146.035 ;
        RECT 354.115 -147.725 354.445 -147.395 ;
        RECT 354.115 -149.085 354.445 -148.755 ;
        RECT 354.115 -150.445 354.445 -150.115 ;
        RECT 354.115 -151.805 354.445 -151.475 ;
        RECT 354.115 -153.165 354.445 -152.835 ;
        RECT 354.115 -154.525 354.445 -154.195 ;
        RECT 354.115 -155.885 354.445 -155.555 ;
        RECT 354.115 -157.245 354.445 -156.915 ;
        RECT 354.115 -158.605 354.445 -158.275 ;
        RECT 354.115 -159.965 354.445 -159.635 ;
        RECT 354.115 -161.325 354.445 -160.995 ;
        RECT 354.115 -162.685 354.445 -162.355 ;
        RECT 354.115 -164.045 354.445 -163.715 ;
        RECT 354.115 -165.405 354.445 -165.075 ;
        RECT 354.115 -166.765 354.445 -166.435 ;
        RECT 354.115 -168.125 354.445 -167.795 ;
        RECT 354.115 -169.485 354.445 -169.155 ;
        RECT 354.115 -170.845 354.445 -170.515 ;
        RECT 354.115 -172.205 354.445 -171.875 ;
        RECT 354.115 -173.565 354.445 -173.235 ;
        RECT 354.115 -174.925 354.445 -174.595 ;
        RECT 354.115 -176.285 354.445 -175.955 ;
        RECT 354.115 -177.645 354.445 -177.315 ;
        RECT 354.115 -183.29 354.445 -182.16 ;
        RECT 354.12 -183.405 354.44 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 355.475 244.04 355.805 245.17 ;
        RECT 355.475 239.875 355.805 240.205 ;
        RECT 355.475 238.515 355.805 238.845 ;
        RECT 355.475 237.155 355.805 237.485 ;
        RECT 355.48 237.155 355.8 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 355.475 -0.845 355.805 -0.515 ;
        RECT 355.475 -2.205 355.805 -1.875 ;
        RECT 355.475 -3.565 355.805 -3.235 ;
        RECT 355.48 -3.565 355.8 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 355.475 -91.965 355.805 -91.635 ;
        RECT 355.475 -93.325 355.805 -92.995 ;
        RECT 355.475 -94.685 355.805 -94.355 ;
        RECT 355.475 -96.045 355.805 -95.715 ;
        RECT 355.475 -97.405 355.805 -97.075 ;
        RECT 355.475 -98.765 355.805 -98.435 ;
        RECT 355.475 -100.125 355.805 -99.795 ;
        RECT 355.475 -101.485 355.805 -101.155 ;
        RECT 355.475 -102.845 355.805 -102.515 ;
        RECT 355.475 -104.205 355.805 -103.875 ;
        RECT 355.475 -105.565 355.805 -105.235 ;
        RECT 355.475 -106.925 355.805 -106.595 ;
        RECT 355.475 -108.285 355.805 -107.955 ;
        RECT 355.475 -109.645 355.805 -109.315 ;
        RECT 355.475 -111.005 355.805 -110.675 ;
        RECT 355.475 -112.365 355.805 -112.035 ;
        RECT 355.475 -113.725 355.805 -113.395 ;
        RECT 355.475 -115.085 355.805 -114.755 ;
        RECT 355.475 -116.445 355.805 -116.115 ;
        RECT 355.475 -117.805 355.805 -117.475 ;
        RECT 355.475 -119.165 355.805 -118.835 ;
        RECT 355.475 -120.525 355.805 -120.195 ;
        RECT 355.475 -121.885 355.805 -121.555 ;
        RECT 355.475 -123.245 355.805 -122.915 ;
        RECT 355.475 -124.605 355.805 -124.275 ;
        RECT 355.475 -125.965 355.805 -125.635 ;
        RECT 355.475 -127.325 355.805 -126.995 ;
        RECT 355.475 -128.685 355.805 -128.355 ;
        RECT 355.475 -130.045 355.805 -129.715 ;
        RECT 355.475 -131.405 355.805 -131.075 ;
        RECT 355.475 -132.765 355.805 -132.435 ;
        RECT 355.475 -134.125 355.805 -133.795 ;
        RECT 355.475 -135.485 355.805 -135.155 ;
        RECT 355.475 -136.845 355.805 -136.515 ;
        RECT 355.475 -138.205 355.805 -137.875 ;
        RECT 355.475 -139.565 355.805 -139.235 ;
        RECT 355.475 -140.925 355.805 -140.595 ;
        RECT 355.475 -142.285 355.805 -141.955 ;
        RECT 355.475 -143.645 355.805 -143.315 ;
        RECT 355.475 -145.005 355.805 -144.675 ;
        RECT 355.475 -146.365 355.805 -146.035 ;
        RECT 355.475 -147.725 355.805 -147.395 ;
        RECT 355.475 -149.085 355.805 -148.755 ;
        RECT 355.475 -150.445 355.805 -150.115 ;
        RECT 355.475 -151.805 355.805 -151.475 ;
        RECT 355.475 -153.165 355.805 -152.835 ;
        RECT 355.475 -154.525 355.805 -154.195 ;
        RECT 355.475 -155.885 355.805 -155.555 ;
        RECT 355.475 -157.245 355.805 -156.915 ;
        RECT 355.475 -158.605 355.805 -158.275 ;
        RECT 355.475 -159.965 355.805 -159.635 ;
        RECT 355.475 -161.325 355.805 -160.995 ;
        RECT 355.475 -162.685 355.805 -162.355 ;
        RECT 355.475 -164.045 355.805 -163.715 ;
        RECT 355.475 -165.405 355.805 -165.075 ;
        RECT 355.475 -166.765 355.805 -166.435 ;
        RECT 355.475 -168.125 355.805 -167.795 ;
        RECT 355.475 -169.485 355.805 -169.155 ;
        RECT 355.475 -170.845 355.805 -170.515 ;
        RECT 355.475 -172.205 355.805 -171.875 ;
        RECT 355.475 -173.565 355.805 -173.235 ;
        RECT 355.475 -174.925 355.805 -174.595 ;
        RECT 355.475 -176.285 355.805 -175.955 ;
        RECT 355.475 -177.645 355.805 -177.315 ;
        RECT 355.475 -183.29 355.805 -182.16 ;
        RECT 355.48 -183.405 355.8 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 356.46 -94.075 356.79 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 356.835 244.04 357.165 245.17 ;
        RECT 356.835 239.875 357.165 240.205 ;
        RECT 356.835 238.515 357.165 238.845 ;
        RECT 356.835 237.155 357.165 237.485 ;
        RECT 356.84 237.155 357.16 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 356.835 -96.045 357.165 -95.715 ;
        RECT 356.835 -97.405 357.165 -97.075 ;
        RECT 356.835 -98.765 357.165 -98.435 ;
        RECT 356.835 -100.125 357.165 -99.795 ;
        RECT 356.835 -101.485 357.165 -101.155 ;
        RECT 356.835 -102.845 357.165 -102.515 ;
        RECT 356.835 -104.205 357.165 -103.875 ;
        RECT 356.835 -105.565 357.165 -105.235 ;
        RECT 356.835 -106.925 357.165 -106.595 ;
        RECT 356.835 -108.285 357.165 -107.955 ;
        RECT 356.835 -109.645 357.165 -109.315 ;
        RECT 356.835 -111.005 357.165 -110.675 ;
        RECT 356.835 -112.365 357.165 -112.035 ;
        RECT 356.835 -113.725 357.165 -113.395 ;
        RECT 356.835 -115.085 357.165 -114.755 ;
        RECT 356.835 -116.445 357.165 -116.115 ;
        RECT 356.835 -117.805 357.165 -117.475 ;
        RECT 356.835 -119.165 357.165 -118.835 ;
        RECT 356.835 -120.525 357.165 -120.195 ;
        RECT 356.835 -121.885 357.165 -121.555 ;
        RECT 356.835 -123.245 357.165 -122.915 ;
        RECT 356.835 -124.605 357.165 -124.275 ;
        RECT 356.835 -125.965 357.165 -125.635 ;
        RECT 356.835 -127.325 357.165 -126.995 ;
        RECT 356.835 -128.685 357.165 -128.355 ;
        RECT 356.835 -130.045 357.165 -129.715 ;
        RECT 356.835 -131.405 357.165 -131.075 ;
        RECT 356.835 -132.765 357.165 -132.435 ;
        RECT 356.835 -134.125 357.165 -133.795 ;
        RECT 356.835 -135.485 357.165 -135.155 ;
        RECT 356.835 -136.845 357.165 -136.515 ;
        RECT 356.835 -138.205 357.165 -137.875 ;
        RECT 356.835 -139.565 357.165 -139.235 ;
        RECT 356.835 -140.925 357.165 -140.595 ;
        RECT 356.835 -142.285 357.165 -141.955 ;
        RECT 356.835 -143.645 357.165 -143.315 ;
        RECT 356.835 -145.005 357.165 -144.675 ;
        RECT 356.835 -146.365 357.165 -146.035 ;
        RECT 356.835 -147.725 357.165 -147.395 ;
        RECT 356.835 -149.085 357.165 -148.755 ;
        RECT 356.835 -150.445 357.165 -150.115 ;
        RECT 356.835 -151.805 357.165 -151.475 ;
        RECT 356.835 -153.165 357.165 -152.835 ;
        RECT 356.835 -154.525 357.165 -154.195 ;
        RECT 356.835 -155.885 357.165 -155.555 ;
        RECT 356.835 -157.245 357.165 -156.915 ;
        RECT 356.835 -158.605 357.165 -158.275 ;
        RECT 356.835 -159.965 357.165 -159.635 ;
        RECT 356.835 -161.325 357.165 -160.995 ;
        RECT 356.835 -162.685 357.165 -162.355 ;
        RECT 356.835 -164.045 357.165 -163.715 ;
        RECT 356.835 -165.405 357.165 -165.075 ;
        RECT 356.835 -166.765 357.165 -166.435 ;
        RECT 356.835 -168.125 357.165 -167.795 ;
        RECT 356.835 -169.485 357.165 -169.155 ;
        RECT 356.835 -170.845 357.165 -170.515 ;
        RECT 356.835 -172.205 357.165 -171.875 ;
        RECT 356.835 -173.565 357.165 -173.235 ;
        RECT 356.835 -174.925 357.165 -174.595 ;
        RECT 356.835 -176.285 357.165 -175.955 ;
        RECT 356.835 -177.645 357.165 -177.315 ;
        RECT 356.835 -183.29 357.165 -182.16 ;
        RECT 356.84 -183.405 357.16 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 358.195 244.04 358.525 245.17 ;
        RECT 358.195 239.875 358.525 240.205 ;
        RECT 358.195 238.515 358.525 238.845 ;
        RECT 358.195 237.155 358.525 237.485 ;
        RECT 358.2 237.155 358.52 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 358.195 -0.845 358.525 -0.515 ;
        RECT 358.195 -2.205 358.525 -1.875 ;
        RECT 358.195 -3.565 358.525 -3.235 ;
        RECT 358.2 -3.565 358.52 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 359.555 244.04 359.885 245.17 ;
        RECT 359.555 239.875 359.885 240.205 ;
        RECT 359.555 238.515 359.885 238.845 ;
        RECT 359.555 237.155 359.885 237.485 ;
        RECT 359.56 237.155 359.88 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 359.555 -0.845 359.885 -0.515 ;
        RECT 359.555 -2.205 359.885 -1.875 ;
        RECT 359.555 -3.565 359.885 -3.235 ;
        RECT 359.56 -3.565 359.88 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 360.915 244.04 361.245 245.17 ;
        RECT 360.915 239.875 361.245 240.205 ;
        RECT 360.915 238.515 361.245 238.845 ;
        RECT 360.915 237.155 361.245 237.485 ;
        RECT 360.92 237.155 361.24 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 360.915 -0.845 361.245 -0.515 ;
        RECT 360.915 -2.205 361.245 -1.875 ;
        RECT 360.915 -3.565 361.245 -3.235 ;
        RECT 360.92 -3.565 361.24 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 360.915 -91.965 361.245 -91.635 ;
        RECT 360.915 -93.325 361.245 -92.995 ;
        RECT 360.915 -94.685 361.245 -94.355 ;
        RECT 360.915 -96.045 361.245 -95.715 ;
        RECT 360.915 -97.405 361.245 -97.075 ;
        RECT 360.915 -98.765 361.245 -98.435 ;
        RECT 360.915 -100.125 361.245 -99.795 ;
        RECT 360.915 -101.485 361.245 -101.155 ;
        RECT 360.915 -102.845 361.245 -102.515 ;
        RECT 360.915 -104.205 361.245 -103.875 ;
        RECT 360.915 -105.565 361.245 -105.235 ;
        RECT 360.915 -106.925 361.245 -106.595 ;
        RECT 360.915 -108.285 361.245 -107.955 ;
        RECT 360.915 -109.645 361.245 -109.315 ;
        RECT 360.915 -111.005 361.245 -110.675 ;
        RECT 360.915 -112.365 361.245 -112.035 ;
        RECT 360.915 -113.725 361.245 -113.395 ;
        RECT 360.915 -115.085 361.245 -114.755 ;
        RECT 360.915 -116.445 361.245 -116.115 ;
        RECT 360.915 -117.805 361.245 -117.475 ;
        RECT 360.915 -119.165 361.245 -118.835 ;
        RECT 360.915 -120.525 361.245 -120.195 ;
        RECT 360.915 -121.885 361.245 -121.555 ;
        RECT 360.915 -123.245 361.245 -122.915 ;
        RECT 360.915 -124.605 361.245 -124.275 ;
        RECT 360.915 -125.965 361.245 -125.635 ;
        RECT 360.915 -127.325 361.245 -126.995 ;
        RECT 360.915 -128.685 361.245 -128.355 ;
        RECT 360.915 -130.045 361.245 -129.715 ;
        RECT 360.915 -131.405 361.245 -131.075 ;
        RECT 360.915 -132.765 361.245 -132.435 ;
        RECT 360.915 -134.125 361.245 -133.795 ;
        RECT 360.915 -135.485 361.245 -135.155 ;
        RECT 360.915 -136.845 361.245 -136.515 ;
        RECT 360.915 -138.205 361.245 -137.875 ;
        RECT 360.915 -139.565 361.245 -139.235 ;
        RECT 360.915 -140.925 361.245 -140.595 ;
        RECT 360.915 -142.285 361.245 -141.955 ;
        RECT 360.915 -143.645 361.245 -143.315 ;
        RECT 360.915 -145.005 361.245 -144.675 ;
        RECT 360.915 -146.365 361.245 -146.035 ;
        RECT 360.915 -147.725 361.245 -147.395 ;
        RECT 360.915 -149.085 361.245 -148.755 ;
        RECT 360.915 -150.445 361.245 -150.115 ;
        RECT 360.915 -151.805 361.245 -151.475 ;
        RECT 360.915 -153.165 361.245 -152.835 ;
        RECT 360.915 -154.525 361.245 -154.195 ;
        RECT 360.915 -155.885 361.245 -155.555 ;
        RECT 360.915 -157.245 361.245 -156.915 ;
        RECT 360.915 -158.605 361.245 -158.275 ;
        RECT 360.915 -159.965 361.245 -159.635 ;
        RECT 360.915 -161.325 361.245 -160.995 ;
        RECT 360.915 -162.685 361.245 -162.355 ;
        RECT 360.915 -164.045 361.245 -163.715 ;
        RECT 360.915 -165.405 361.245 -165.075 ;
        RECT 360.915 -166.765 361.245 -166.435 ;
        RECT 360.915 -168.125 361.245 -167.795 ;
        RECT 360.915 -169.485 361.245 -169.155 ;
        RECT 360.915 -170.845 361.245 -170.515 ;
        RECT 360.915 -172.205 361.245 -171.875 ;
        RECT 360.915 -173.565 361.245 -173.235 ;
        RECT 360.915 -174.925 361.245 -174.595 ;
        RECT 360.915 -176.285 361.245 -175.955 ;
        RECT 360.915 -177.645 361.245 -177.315 ;
        RECT 360.915 -183.29 361.245 -182.16 ;
        RECT 360.92 -183.405 361.24 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 362.275 244.04 362.605 245.17 ;
        RECT 362.275 239.875 362.605 240.205 ;
        RECT 362.275 238.515 362.605 238.845 ;
        RECT 362.275 237.155 362.605 237.485 ;
        RECT 362.28 237.155 362.6 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 362.275 -96.045 362.605 -95.715 ;
        RECT 362.275 -97.405 362.605 -97.075 ;
        RECT 362.275 -98.765 362.605 -98.435 ;
        RECT 362.275 -100.125 362.605 -99.795 ;
        RECT 362.275 -101.485 362.605 -101.155 ;
        RECT 362.275 -102.845 362.605 -102.515 ;
        RECT 362.275 -104.205 362.605 -103.875 ;
        RECT 362.275 -105.565 362.605 -105.235 ;
        RECT 362.275 -106.925 362.605 -106.595 ;
        RECT 362.275 -108.285 362.605 -107.955 ;
        RECT 362.275 -109.645 362.605 -109.315 ;
        RECT 362.275 -111.005 362.605 -110.675 ;
        RECT 362.275 -112.365 362.605 -112.035 ;
        RECT 362.275 -113.725 362.605 -113.395 ;
        RECT 362.275 -115.085 362.605 -114.755 ;
        RECT 362.275 -116.445 362.605 -116.115 ;
        RECT 362.275 -117.805 362.605 -117.475 ;
        RECT 362.275 -119.165 362.605 -118.835 ;
        RECT 362.275 -120.525 362.605 -120.195 ;
        RECT 362.275 -121.885 362.605 -121.555 ;
        RECT 362.275 -123.245 362.605 -122.915 ;
        RECT 362.275 -124.605 362.605 -124.275 ;
        RECT 362.275 -125.965 362.605 -125.635 ;
        RECT 362.275 -127.325 362.605 -126.995 ;
        RECT 362.275 -128.685 362.605 -128.355 ;
        RECT 362.275 -130.045 362.605 -129.715 ;
        RECT 362.275 -131.405 362.605 -131.075 ;
        RECT 362.275 -132.765 362.605 -132.435 ;
        RECT 362.275 -134.125 362.605 -133.795 ;
        RECT 362.275 -135.485 362.605 -135.155 ;
        RECT 362.275 -136.845 362.605 -136.515 ;
        RECT 362.275 -138.205 362.605 -137.875 ;
        RECT 362.275 -139.565 362.605 -139.235 ;
        RECT 362.275 -140.925 362.605 -140.595 ;
        RECT 362.275 -142.285 362.605 -141.955 ;
        RECT 362.275 -143.645 362.605 -143.315 ;
        RECT 362.275 -145.005 362.605 -144.675 ;
        RECT 362.275 -146.365 362.605 -146.035 ;
        RECT 362.275 -147.725 362.605 -147.395 ;
        RECT 362.275 -149.085 362.605 -148.755 ;
        RECT 362.275 -150.445 362.605 -150.115 ;
        RECT 362.275 -151.805 362.605 -151.475 ;
        RECT 362.275 -153.165 362.605 -152.835 ;
        RECT 362.275 -154.525 362.605 -154.195 ;
        RECT 362.275 -155.885 362.605 -155.555 ;
        RECT 362.275 -157.245 362.605 -156.915 ;
        RECT 362.275 -158.605 362.605 -158.275 ;
        RECT 362.275 -159.965 362.605 -159.635 ;
        RECT 362.275 -161.325 362.605 -160.995 ;
        RECT 362.275 -162.685 362.605 -162.355 ;
        RECT 362.275 -164.045 362.605 -163.715 ;
        RECT 362.275 -165.405 362.605 -165.075 ;
        RECT 362.275 -166.765 362.605 -166.435 ;
        RECT 362.275 -168.125 362.605 -167.795 ;
        RECT 362.275 -169.485 362.605 -169.155 ;
        RECT 362.275 -170.845 362.605 -170.515 ;
        RECT 362.275 -172.205 362.605 -171.875 ;
        RECT 362.275 -173.565 362.605 -173.235 ;
        RECT 362.275 -174.925 362.605 -174.595 ;
        RECT 362.275 -176.285 362.605 -175.955 ;
        RECT 362.275 -177.645 362.605 -177.315 ;
        RECT 362.275 -183.29 362.605 -182.16 ;
        RECT 362.28 -183.405 362.6 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 362.56 -94.075 362.89 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 363.635 244.04 363.965 245.17 ;
        RECT 363.635 239.875 363.965 240.205 ;
        RECT 363.635 238.515 363.965 238.845 ;
        RECT 363.635 237.155 363.965 237.485 ;
        RECT 363.64 237.155 363.96 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 364.995 244.04 365.325 245.17 ;
        RECT 364.995 239.875 365.325 240.205 ;
        RECT 364.995 238.515 365.325 238.845 ;
        RECT 364.995 237.155 365.325 237.485 ;
        RECT 365 237.155 365.32 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 364.995 -0.845 365.325 -0.515 ;
        RECT 364.995 -2.205 365.325 -1.875 ;
        RECT 364.995 -3.565 365.325 -3.235 ;
        RECT 365 -3.565 365.32 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 366.355 244.04 366.685 245.17 ;
        RECT 366.355 239.875 366.685 240.205 ;
        RECT 366.355 238.515 366.685 238.845 ;
        RECT 366.355 237.155 366.685 237.485 ;
        RECT 366.36 237.155 366.68 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 366.355 -0.845 366.685 -0.515 ;
        RECT 366.355 -2.205 366.685 -1.875 ;
        RECT 366.355 -3.565 366.685 -3.235 ;
        RECT 366.36 -3.565 366.68 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 366.355 -91.965 366.685 -91.635 ;
        RECT 366.355 -93.325 366.685 -92.995 ;
        RECT 366.355 -94.685 366.685 -94.355 ;
        RECT 366.355 -96.045 366.685 -95.715 ;
        RECT 366.355 -97.405 366.685 -97.075 ;
        RECT 366.355 -98.765 366.685 -98.435 ;
        RECT 366.355 -100.125 366.685 -99.795 ;
        RECT 366.355 -101.485 366.685 -101.155 ;
        RECT 366.355 -102.845 366.685 -102.515 ;
        RECT 366.355 -104.205 366.685 -103.875 ;
        RECT 366.355 -105.565 366.685 -105.235 ;
        RECT 366.355 -106.925 366.685 -106.595 ;
        RECT 366.355 -108.285 366.685 -107.955 ;
        RECT 366.355 -109.645 366.685 -109.315 ;
        RECT 366.355 -111.005 366.685 -110.675 ;
        RECT 366.355 -112.365 366.685 -112.035 ;
        RECT 366.355 -113.725 366.685 -113.395 ;
        RECT 366.355 -115.085 366.685 -114.755 ;
        RECT 366.355 -116.445 366.685 -116.115 ;
        RECT 366.355 -117.805 366.685 -117.475 ;
        RECT 366.355 -119.165 366.685 -118.835 ;
        RECT 366.355 -120.525 366.685 -120.195 ;
        RECT 366.355 -121.885 366.685 -121.555 ;
        RECT 366.355 -123.245 366.685 -122.915 ;
        RECT 366.355 -124.605 366.685 -124.275 ;
        RECT 366.355 -125.965 366.685 -125.635 ;
        RECT 366.355 -127.325 366.685 -126.995 ;
        RECT 366.355 -128.685 366.685 -128.355 ;
        RECT 366.355 -130.045 366.685 -129.715 ;
        RECT 366.355 -131.405 366.685 -131.075 ;
        RECT 366.355 -132.765 366.685 -132.435 ;
        RECT 366.355 -134.125 366.685 -133.795 ;
        RECT 366.355 -135.485 366.685 -135.155 ;
        RECT 366.355 -136.845 366.685 -136.515 ;
        RECT 366.355 -138.205 366.685 -137.875 ;
        RECT 366.355 -139.565 366.685 -139.235 ;
        RECT 366.355 -140.925 366.685 -140.595 ;
        RECT 366.355 -142.285 366.685 -141.955 ;
        RECT 366.355 -143.645 366.685 -143.315 ;
        RECT 366.355 -145.005 366.685 -144.675 ;
        RECT 366.355 -146.365 366.685 -146.035 ;
        RECT 366.355 -147.725 366.685 -147.395 ;
        RECT 366.355 -149.085 366.685 -148.755 ;
        RECT 366.355 -150.445 366.685 -150.115 ;
        RECT 366.355 -151.805 366.685 -151.475 ;
        RECT 366.355 -153.165 366.685 -152.835 ;
        RECT 366.355 -154.525 366.685 -154.195 ;
        RECT 366.355 -155.885 366.685 -155.555 ;
        RECT 366.355 -157.245 366.685 -156.915 ;
        RECT 366.355 -158.605 366.685 -158.275 ;
        RECT 366.355 -159.965 366.685 -159.635 ;
        RECT 366.355 -161.325 366.685 -160.995 ;
        RECT 366.355 -162.685 366.685 -162.355 ;
        RECT 366.355 -164.045 366.685 -163.715 ;
        RECT 366.355 -165.405 366.685 -165.075 ;
        RECT 366.355 -166.765 366.685 -166.435 ;
        RECT 366.355 -168.125 366.685 -167.795 ;
        RECT 366.355 -169.485 366.685 -169.155 ;
        RECT 366.355 -170.845 366.685 -170.515 ;
        RECT 366.355 -172.205 366.685 -171.875 ;
        RECT 366.355 -173.565 366.685 -173.235 ;
        RECT 366.355 -174.925 366.685 -174.595 ;
        RECT 366.355 -176.285 366.685 -175.955 ;
        RECT 366.355 -177.645 366.685 -177.315 ;
        RECT 366.355 -183.29 366.685 -182.16 ;
        RECT 366.36 -183.405 366.68 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 367.715 244.04 368.045 245.17 ;
        RECT 367.715 239.875 368.045 240.205 ;
        RECT 367.715 238.515 368.045 238.845 ;
        RECT 367.715 237.155 368.045 237.485 ;
        RECT 367.72 237.155 368.04 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 367.715 -0.845 368.045 -0.515 ;
        RECT 367.715 -2.205 368.045 -1.875 ;
        RECT 367.715 -3.565 368.045 -3.235 ;
        RECT 367.72 -3.565 368.04 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 367.715 -91.965 368.045 -91.635 ;
        RECT 367.715 -93.325 368.045 -92.995 ;
        RECT 367.715 -94.685 368.045 -94.355 ;
        RECT 367.715 -96.045 368.045 -95.715 ;
        RECT 367.715 -97.405 368.045 -97.075 ;
        RECT 367.715 -98.765 368.045 -98.435 ;
        RECT 367.715 -100.125 368.045 -99.795 ;
        RECT 367.715 -101.485 368.045 -101.155 ;
        RECT 367.715 -102.845 368.045 -102.515 ;
        RECT 367.715 -104.205 368.045 -103.875 ;
        RECT 367.715 -105.565 368.045 -105.235 ;
        RECT 367.715 -106.925 368.045 -106.595 ;
        RECT 367.715 -108.285 368.045 -107.955 ;
        RECT 367.715 -109.645 368.045 -109.315 ;
        RECT 367.715 -111.005 368.045 -110.675 ;
        RECT 367.715 -112.365 368.045 -112.035 ;
        RECT 367.715 -113.725 368.045 -113.395 ;
        RECT 367.715 -115.085 368.045 -114.755 ;
        RECT 367.715 -116.445 368.045 -116.115 ;
        RECT 367.715 -117.805 368.045 -117.475 ;
        RECT 367.715 -119.165 368.045 -118.835 ;
        RECT 367.715 -120.525 368.045 -120.195 ;
        RECT 367.715 -121.885 368.045 -121.555 ;
        RECT 367.715 -123.245 368.045 -122.915 ;
        RECT 367.715 -124.605 368.045 -124.275 ;
        RECT 367.715 -125.965 368.045 -125.635 ;
        RECT 367.715 -127.325 368.045 -126.995 ;
        RECT 367.715 -128.685 368.045 -128.355 ;
        RECT 367.715 -130.045 368.045 -129.715 ;
        RECT 367.715 -131.405 368.045 -131.075 ;
        RECT 367.715 -132.765 368.045 -132.435 ;
        RECT 367.715 -134.125 368.045 -133.795 ;
        RECT 367.715 -135.485 368.045 -135.155 ;
        RECT 367.715 -136.845 368.045 -136.515 ;
        RECT 367.715 -138.205 368.045 -137.875 ;
        RECT 367.715 -139.565 368.045 -139.235 ;
        RECT 367.715 -140.925 368.045 -140.595 ;
        RECT 367.715 -142.285 368.045 -141.955 ;
        RECT 367.715 -143.645 368.045 -143.315 ;
        RECT 367.715 -145.005 368.045 -144.675 ;
        RECT 367.715 -146.365 368.045 -146.035 ;
        RECT 367.715 -147.725 368.045 -147.395 ;
        RECT 367.715 -149.085 368.045 -148.755 ;
        RECT 367.715 -150.445 368.045 -150.115 ;
        RECT 367.715 -151.805 368.045 -151.475 ;
        RECT 367.715 -153.165 368.045 -152.835 ;
        RECT 367.715 -154.525 368.045 -154.195 ;
        RECT 367.715 -155.885 368.045 -155.555 ;
        RECT 367.715 -157.245 368.045 -156.915 ;
        RECT 367.715 -158.605 368.045 -158.275 ;
        RECT 367.715 -159.965 368.045 -159.635 ;
        RECT 367.715 -161.325 368.045 -160.995 ;
        RECT 367.715 -162.685 368.045 -162.355 ;
        RECT 367.715 -164.045 368.045 -163.715 ;
        RECT 367.715 -165.405 368.045 -165.075 ;
        RECT 367.715 -166.765 368.045 -166.435 ;
        RECT 367.715 -168.125 368.045 -167.795 ;
        RECT 367.715 -169.485 368.045 -169.155 ;
        RECT 367.715 -170.845 368.045 -170.515 ;
        RECT 367.715 -172.205 368.045 -171.875 ;
        RECT 367.715 -173.565 368.045 -173.235 ;
        RECT 367.715 -174.925 368.045 -174.595 ;
        RECT 367.715 -176.285 368.045 -175.955 ;
        RECT 367.715 -177.645 368.045 -177.315 ;
        RECT 367.715 -183.29 368.045 -182.16 ;
        RECT 367.72 -183.405 368.04 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 368.66 -94.075 368.99 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 369.075 244.04 369.405 245.17 ;
        RECT 369.075 239.875 369.405 240.205 ;
        RECT 369.075 238.515 369.405 238.845 ;
        RECT 369.075 237.155 369.405 237.485 ;
        RECT 369.08 237.155 369.4 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 369.075 -96.045 369.405 -95.715 ;
        RECT 369.075 -97.405 369.405 -97.075 ;
        RECT 369.075 -98.765 369.405 -98.435 ;
        RECT 369.075 -100.125 369.405 -99.795 ;
        RECT 369.075 -101.485 369.405 -101.155 ;
        RECT 369.075 -102.845 369.405 -102.515 ;
        RECT 369.075 -104.205 369.405 -103.875 ;
        RECT 369.075 -105.565 369.405 -105.235 ;
        RECT 369.075 -106.925 369.405 -106.595 ;
        RECT 369.075 -108.285 369.405 -107.955 ;
        RECT 369.075 -109.645 369.405 -109.315 ;
        RECT 369.075 -111.005 369.405 -110.675 ;
        RECT 369.075 -112.365 369.405 -112.035 ;
        RECT 369.075 -113.725 369.405 -113.395 ;
        RECT 369.075 -115.085 369.405 -114.755 ;
        RECT 369.075 -116.445 369.405 -116.115 ;
        RECT 369.075 -117.805 369.405 -117.475 ;
        RECT 369.075 -119.165 369.405 -118.835 ;
        RECT 369.075 -120.525 369.405 -120.195 ;
        RECT 369.075 -121.885 369.405 -121.555 ;
        RECT 369.075 -123.245 369.405 -122.915 ;
        RECT 369.075 -124.605 369.405 -124.275 ;
        RECT 369.075 -125.965 369.405 -125.635 ;
        RECT 369.075 -127.325 369.405 -126.995 ;
        RECT 369.075 -128.685 369.405 -128.355 ;
        RECT 369.075 -130.045 369.405 -129.715 ;
        RECT 369.075 -131.405 369.405 -131.075 ;
        RECT 369.075 -132.765 369.405 -132.435 ;
        RECT 369.075 -134.125 369.405 -133.795 ;
        RECT 369.075 -135.485 369.405 -135.155 ;
        RECT 369.075 -136.845 369.405 -136.515 ;
        RECT 369.075 -138.205 369.405 -137.875 ;
        RECT 369.075 -139.565 369.405 -139.235 ;
        RECT 369.075 -140.925 369.405 -140.595 ;
        RECT 369.075 -142.285 369.405 -141.955 ;
        RECT 369.075 -143.645 369.405 -143.315 ;
        RECT 369.075 -145.005 369.405 -144.675 ;
        RECT 369.075 -146.365 369.405 -146.035 ;
        RECT 369.075 -147.725 369.405 -147.395 ;
        RECT 369.075 -149.085 369.405 -148.755 ;
        RECT 369.075 -150.445 369.405 -150.115 ;
        RECT 369.075 -151.805 369.405 -151.475 ;
        RECT 369.075 -153.165 369.405 -152.835 ;
        RECT 369.075 -154.525 369.405 -154.195 ;
        RECT 369.075 -155.885 369.405 -155.555 ;
        RECT 369.075 -157.245 369.405 -156.915 ;
        RECT 369.075 -158.605 369.405 -158.275 ;
        RECT 369.075 -159.965 369.405 -159.635 ;
        RECT 369.075 -161.325 369.405 -160.995 ;
        RECT 369.075 -162.685 369.405 -162.355 ;
        RECT 369.075 -164.045 369.405 -163.715 ;
        RECT 369.075 -165.405 369.405 -165.075 ;
        RECT 369.075 -166.765 369.405 -166.435 ;
        RECT 369.075 -168.125 369.405 -167.795 ;
        RECT 369.075 -169.485 369.405 -169.155 ;
        RECT 369.075 -170.845 369.405 -170.515 ;
        RECT 369.075 -172.205 369.405 -171.875 ;
        RECT 369.075 -173.565 369.405 -173.235 ;
        RECT 369.075 -174.925 369.405 -174.595 ;
        RECT 369.075 -176.285 369.405 -175.955 ;
        RECT 369.075 -177.645 369.405 -177.315 ;
        RECT 369.075 -183.29 369.405 -182.16 ;
        RECT 369.08 -183.405 369.4 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 370.435 244.04 370.765 245.17 ;
        RECT 370.435 239.875 370.765 240.205 ;
        RECT 370.435 238.515 370.765 238.845 ;
        RECT 370.435 237.155 370.765 237.485 ;
        RECT 370.44 237.155 370.76 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 370.435 -0.845 370.765 -0.515 ;
        RECT 370.435 -2.205 370.765 -1.875 ;
        RECT 370.435 -3.565 370.765 -3.235 ;
        RECT 370.44 -3.565 370.76 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 371.795 244.04 372.125 245.17 ;
        RECT 371.795 239.875 372.125 240.205 ;
        RECT 371.795 238.515 372.125 238.845 ;
        RECT 371.795 237.155 372.125 237.485 ;
        RECT 371.8 237.155 372.12 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 371.795 -0.845 372.125 -0.515 ;
        RECT 371.795 -2.205 372.125 -1.875 ;
        RECT 371.795 -3.565 372.125 -3.235 ;
        RECT 371.8 -3.565 372.12 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 373.155 244.04 373.485 245.17 ;
        RECT 373.155 239.875 373.485 240.205 ;
        RECT 373.155 238.515 373.485 238.845 ;
        RECT 373.155 237.155 373.485 237.485 ;
        RECT 373.16 237.155 373.48 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 373.155 -0.845 373.485 -0.515 ;
        RECT 373.155 -2.205 373.485 -1.875 ;
        RECT 373.155 -3.565 373.485 -3.235 ;
        RECT 373.16 -3.565 373.48 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 373.155 -104.205 373.485 -103.875 ;
        RECT 373.155 -105.565 373.485 -105.235 ;
        RECT 373.155 -106.925 373.485 -106.595 ;
        RECT 373.155 -108.285 373.485 -107.955 ;
        RECT 373.155 -109.645 373.485 -109.315 ;
        RECT 373.155 -111.005 373.485 -110.675 ;
        RECT 373.155 -112.365 373.485 -112.035 ;
        RECT 373.155 -113.725 373.485 -113.395 ;
        RECT 373.155 -115.085 373.485 -114.755 ;
        RECT 373.155 -116.445 373.485 -116.115 ;
        RECT 373.155 -117.805 373.485 -117.475 ;
        RECT 373.155 -119.165 373.485 -118.835 ;
        RECT 373.155 -120.525 373.485 -120.195 ;
        RECT 373.155 -121.885 373.485 -121.555 ;
        RECT 373.155 -123.245 373.485 -122.915 ;
        RECT 373.155 -124.605 373.485 -124.275 ;
        RECT 373.155 -125.965 373.485 -125.635 ;
        RECT 373.155 -127.325 373.485 -126.995 ;
        RECT 373.155 -128.685 373.485 -128.355 ;
        RECT 373.155 -130.045 373.485 -129.715 ;
        RECT 373.155 -131.405 373.485 -131.075 ;
        RECT 373.155 -132.765 373.485 -132.435 ;
        RECT 373.155 -134.125 373.485 -133.795 ;
        RECT 373.155 -135.485 373.485 -135.155 ;
        RECT 373.155 -136.845 373.485 -136.515 ;
        RECT 373.155 -138.205 373.485 -137.875 ;
        RECT 373.155 -139.565 373.485 -139.235 ;
        RECT 373.155 -140.925 373.485 -140.595 ;
        RECT 373.155 -142.285 373.485 -141.955 ;
        RECT 373.155 -143.645 373.485 -143.315 ;
        RECT 373.155 -145.005 373.485 -144.675 ;
        RECT 373.155 -146.365 373.485 -146.035 ;
        RECT 373.155 -147.725 373.485 -147.395 ;
        RECT 373.155 -149.085 373.485 -148.755 ;
        RECT 373.155 -150.445 373.485 -150.115 ;
        RECT 373.155 -151.805 373.485 -151.475 ;
        RECT 373.155 -153.165 373.485 -152.835 ;
        RECT 373.155 -154.525 373.485 -154.195 ;
        RECT 373.155 -155.885 373.485 -155.555 ;
        RECT 373.155 -157.245 373.485 -156.915 ;
        RECT 373.155 -158.605 373.485 -158.275 ;
        RECT 373.155 -159.965 373.485 -159.635 ;
        RECT 373.155 -161.325 373.485 -160.995 ;
        RECT 373.155 -162.685 373.485 -162.355 ;
        RECT 373.155 -164.045 373.485 -163.715 ;
        RECT 373.155 -165.405 373.485 -165.075 ;
        RECT 373.155 -166.765 373.485 -166.435 ;
        RECT 373.155 -168.125 373.485 -167.795 ;
        RECT 373.155 -169.485 373.485 -169.155 ;
        RECT 373.155 -170.845 373.485 -170.515 ;
        RECT 373.155 -172.205 373.485 -171.875 ;
        RECT 373.155 -173.565 373.485 -173.235 ;
        RECT 373.155 -174.925 373.485 -174.595 ;
        RECT 373.155 -176.285 373.485 -175.955 ;
        RECT 373.155 -177.645 373.485 -177.315 ;
        RECT 373.155 -183.29 373.485 -182.16 ;
        RECT 373.16 -183.405 373.48 -90.96 ;
        RECT 373.155 -91.965 373.485 -91.635 ;
        RECT 373.155 -93.325 373.485 -92.995 ;
        RECT 373.155 -94.685 373.485 -94.355 ;
        RECT 373.155 -96.045 373.485 -95.715 ;
        RECT 373.155 -97.405 373.485 -97.075 ;
        RECT 373.155 -98.765 373.485 -98.435 ;
        RECT 373.155 -100.125 373.485 -99.795 ;
        RECT 373.155 -101.485 373.485 -101.155 ;
        RECT 373.155 -102.845 373.485 -102.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 306.515 -0.845 306.845 -0.515 ;
        RECT 306.515 -2.205 306.845 -1.875 ;
        RECT 306.515 -3.565 306.845 -3.235 ;
        RECT 306.52 -3.565 306.84 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 306.515 -91.965 306.845 -91.635 ;
        RECT 306.515 -93.325 306.845 -92.995 ;
        RECT 306.515 -94.685 306.845 -94.355 ;
        RECT 306.515 -96.045 306.845 -95.715 ;
        RECT 306.515 -97.405 306.845 -97.075 ;
        RECT 306.515 -98.765 306.845 -98.435 ;
        RECT 306.515 -100.125 306.845 -99.795 ;
        RECT 306.515 -101.485 306.845 -101.155 ;
        RECT 306.515 -102.845 306.845 -102.515 ;
        RECT 306.515 -104.205 306.845 -103.875 ;
        RECT 306.515 -105.565 306.845 -105.235 ;
        RECT 306.515 -106.925 306.845 -106.595 ;
        RECT 306.515 -108.285 306.845 -107.955 ;
        RECT 306.515 -109.645 306.845 -109.315 ;
        RECT 306.515 -111.005 306.845 -110.675 ;
        RECT 306.515 -112.365 306.845 -112.035 ;
        RECT 306.515 -113.725 306.845 -113.395 ;
        RECT 306.515 -115.085 306.845 -114.755 ;
        RECT 306.515 -116.445 306.845 -116.115 ;
        RECT 306.515 -117.805 306.845 -117.475 ;
        RECT 306.515 -119.165 306.845 -118.835 ;
        RECT 306.515 -120.525 306.845 -120.195 ;
        RECT 306.515 -121.885 306.845 -121.555 ;
        RECT 306.515 -123.245 306.845 -122.915 ;
        RECT 306.515 -124.605 306.845 -124.275 ;
        RECT 306.515 -125.965 306.845 -125.635 ;
        RECT 306.515 -127.325 306.845 -126.995 ;
        RECT 306.515 -128.685 306.845 -128.355 ;
        RECT 306.515 -130.045 306.845 -129.715 ;
        RECT 306.515 -131.405 306.845 -131.075 ;
        RECT 306.515 -132.765 306.845 -132.435 ;
        RECT 306.515 -134.125 306.845 -133.795 ;
        RECT 306.515 -135.485 306.845 -135.155 ;
        RECT 306.515 -136.845 306.845 -136.515 ;
        RECT 306.515 -138.205 306.845 -137.875 ;
        RECT 306.515 -139.565 306.845 -139.235 ;
        RECT 306.515 -140.925 306.845 -140.595 ;
        RECT 306.515 -142.285 306.845 -141.955 ;
        RECT 306.515 -143.645 306.845 -143.315 ;
        RECT 306.515 -145.005 306.845 -144.675 ;
        RECT 306.515 -146.365 306.845 -146.035 ;
        RECT 306.515 -147.725 306.845 -147.395 ;
        RECT 306.515 -149.085 306.845 -148.755 ;
        RECT 306.515 -150.445 306.845 -150.115 ;
        RECT 306.515 -151.805 306.845 -151.475 ;
        RECT 306.515 -153.165 306.845 -152.835 ;
        RECT 306.515 -154.525 306.845 -154.195 ;
        RECT 306.515 -155.885 306.845 -155.555 ;
        RECT 306.515 -157.245 306.845 -156.915 ;
        RECT 306.515 -158.605 306.845 -158.275 ;
        RECT 306.515 -159.965 306.845 -159.635 ;
        RECT 306.515 -161.325 306.845 -160.995 ;
        RECT 306.515 -162.685 306.845 -162.355 ;
        RECT 306.515 -164.045 306.845 -163.715 ;
        RECT 306.515 -165.405 306.845 -165.075 ;
        RECT 306.515 -166.765 306.845 -166.435 ;
        RECT 306.515 -168.125 306.845 -167.795 ;
        RECT 306.515 -169.485 306.845 -169.155 ;
        RECT 306.515 -170.845 306.845 -170.515 ;
        RECT 306.515 -172.205 306.845 -171.875 ;
        RECT 306.515 -173.565 306.845 -173.235 ;
        RECT 306.515 -174.925 306.845 -174.595 ;
        RECT 306.515 -176.285 306.845 -175.955 ;
        RECT 306.515 -177.645 306.845 -177.315 ;
        RECT 306.515 -183.29 306.845 -182.16 ;
        RECT 306.52 -183.405 306.84 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 307.66 -94.075 307.99 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 307.875 244.04 308.205 245.17 ;
        RECT 307.875 239.875 308.205 240.205 ;
        RECT 307.875 238.515 308.205 238.845 ;
        RECT 307.875 237.155 308.205 237.485 ;
        RECT 307.88 237.155 308.2 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 307.875 -96.045 308.205 -95.715 ;
        RECT 307.875 -97.405 308.205 -97.075 ;
        RECT 307.875 -98.765 308.205 -98.435 ;
        RECT 307.875 -100.125 308.205 -99.795 ;
        RECT 307.875 -101.485 308.205 -101.155 ;
        RECT 307.875 -102.845 308.205 -102.515 ;
        RECT 307.875 -104.205 308.205 -103.875 ;
        RECT 307.875 -105.565 308.205 -105.235 ;
        RECT 307.875 -106.925 308.205 -106.595 ;
        RECT 307.875 -108.285 308.205 -107.955 ;
        RECT 307.875 -109.645 308.205 -109.315 ;
        RECT 307.875 -111.005 308.205 -110.675 ;
        RECT 307.875 -112.365 308.205 -112.035 ;
        RECT 307.875 -113.725 308.205 -113.395 ;
        RECT 307.875 -115.085 308.205 -114.755 ;
        RECT 307.875 -116.445 308.205 -116.115 ;
        RECT 307.875 -117.805 308.205 -117.475 ;
        RECT 307.875 -119.165 308.205 -118.835 ;
        RECT 307.875 -120.525 308.205 -120.195 ;
        RECT 307.875 -121.885 308.205 -121.555 ;
        RECT 307.875 -123.245 308.205 -122.915 ;
        RECT 307.875 -124.605 308.205 -124.275 ;
        RECT 307.875 -125.965 308.205 -125.635 ;
        RECT 307.875 -127.325 308.205 -126.995 ;
        RECT 307.875 -128.685 308.205 -128.355 ;
        RECT 307.875 -130.045 308.205 -129.715 ;
        RECT 307.875 -131.405 308.205 -131.075 ;
        RECT 307.875 -132.765 308.205 -132.435 ;
        RECT 307.875 -134.125 308.205 -133.795 ;
        RECT 307.875 -135.485 308.205 -135.155 ;
        RECT 307.875 -136.845 308.205 -136.515 ;
        RECT 307.875 -138.205 308.205 -137.875 ;
        RECT 307.875 -139.565 308.205 -139.235 ;
        RECT 307.875 -140.925 308.205 -140.595 ;
        RECT 307.875 -142.285 308.205 -141.955 ;
        RECT 307.875 -143.645 308.205 -143.315 ;
        RECT 307.875 -145.005 308.205 -144.675 ;
        RECT 307.875 -146.365 308.205 -146.035 ;
        RECT 307.875 -147.725 308.205 -147.395 ;
        RECT 307.875 -149.085 308.205 -148.755 ;
        RECT 307.875 -150.445 308.205 -150.115 ;
        RECT 307.875 -151.805 308.205 -151.475 ;
        RECT 307.875 -153.165 308.205 -152.835 ;
        RECT 307.875 -154.525 308.205 -154.195 ;
        RECT 307.875 -155.885 308.205 -155.555 ;
        RECT 307.875 -157.245 308.205 -156.915 ;
        RECT 307.875 -158.605 308.205 -158.275 ;
        RECT 307.875 -159.965 308.205 -159.635 ;
        RECT 307.875 -161.325 308.205 -160.995 ;
        RECT 307.875 -162.685 308.205 -162.355 ;
        RECT 307.875 -164.045 308.205 -163.715 ;
        RECT 307.875 -165.405 308.205 -165.075 ;
        RECT 307.875 -166.765 308.205 -166.435 ;
        RECT 307.875 -168.125 308.205 -167.795 ;
        RECT 307.875 -169.485 308.205 -169.155 ;
        RECT 307.875 -170.845 308.205 -170.515 ;
        RECT 307.875 -172.205 308.205 -171.875 ;
        RECT 307.875 -173.565 308.205 -173.235 ;
        RECT 307.875 -174.925 308.205 -174.595 ;
        RECT 307.875 -176.285 308.205 -175.955 ;
        RECT 307.875 -177.645 308.205 -177.315 ;
        RECT 307.875 -183.29 308.205 -182.16 ;
        RECT 307.88 -183.405 308.2 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 309.235 244.04 309.565 245.17 ;
        RECT 309.235 239.875 309.565 240.205 ;
        RECT 309.235 238.515 309.565 238.845 ;
        RECT 309.235 237.155 309.565 237.485 ;
        RECT 309.24 237.155 309.56 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 309.235 -0.845 309.565 -0.515 ;
        RECT 309.235 -2.205 309.565 -1.875 ;
        RECT 309.235 -3.565 309.565 -3.235 ;
        RECT 309.24 -3.565 309.56 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 310.595 244.04 310.925 245.17 ;
        RECT 310.595 239.875 310.925 240.205 ;
        RECT 310.595 238.515 310.925 238.845 ;
        RECT 310.595 237.155 310.925 237.485 ;
        RECT 310.6 237.155 310.92 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 310.595 -0.845 310.925 -0.515 ;
        RECT 310.595 -2.205 310.925 -1.875 ;
        RECT 310.595 -3.565 310.925 -3.235 ;
        RECT 310.6 -3.565 310.92 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 311.955 244.04 312.285 245.17 ;
        RECT 311.955 239.875 312.285 240.205 ;
        RECT 311.955 238.515 312.285 238.845 ;
        RECT 311.955 237.155 312.285 237.485 ;
        RECT 311.96 237.155 312.28 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 311.955 -0.845 312.285 -0.515 ;
        RECT 311.955 -2.205 312.285 -1.875 ;
        RECT 311.955 -3.565 312.285 -3.235 ;
        RECT 311.96 -3.565 312.28 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 311.955 -91.965 312.285 -91.635 ;
        RECT 311.955 -93.325 312.285 -92.995 ;
        RECT 311.955 -94.685 312.285 -94.355 ;
        RECT 311.955 -96.045 312.285 -95.715 ;
        RECT 311.955 -97.405 312.285 -97.075 ;
        RECT 311.955 -98.765 312.285 -98.435 ;
        RECT 311.955 -100.125 312.285 -99.795 ;
        RECT 311.955 -101.485 312.285 -101.155 ;
        RECT 311.955 -102.845 312.285 -102.515 ;
        RECT 311.955 -104.205 312.285 -103.875 ;
        RECT 311.955 -105.565 312.285 -105.235 ;
        RECT 311.955 -106.925 312.285 -106.595 ;
        RECT 311.955 -108.285 312.285 -107.955 ;
        RECT 311.955 -109.645 312.285 -109.315 ;
        RECT 311.955 -111.005 312.285 -110.675 ;
        RECT 311.955 -112.365 312.285 -112.035 ;
        RECT 311.955 -113.725 312.285 -113.395 ;
        RECT 311.955 -115.085 312.285 -114.755 ;
        RECT 311.955 -116.445 312.285 -116.115 ;
        RECT 311.955 -117.805 312.285 -117.475 ;
        RECT 311.955 -119.165 312.285 -118.835 ;
        RECT 311.955 -120.525 312.285 -120.195 ;
        RECT 311.955 -121.885 312.285 -121.555 ;
        RECT 311.955 -123.245 312.285 -122.915 ;
        RECT 311.955 -124.605 312.285 -124.275 ;
        RECT 311.955 -125.965 312.285 -125.635 ;
        RECT 311.955 -127.325 312.285 -126.995 ;
        RECT 311.955 -128.685 312.285 -128.355 ;
        RECT 311.955 -130.045 312.285 -129.715 ;
        RECT 311.955 -131.405 312.285 -131.075 ;
        RECT 311.955 -132.765 312.285 -132.435 ;
        RECT 311.955 -134.125 312.285 -133.795 ;
        RECT 311.955 -135.485 312.285 -135.155 ;
        RECT 311.955 -136.845 312.285 -136.515 ;
        RECT 311.955 -138.205 312.285 -137.875 ;
        RECT 311.955 -139.565 312.285 -139.235 ;
        RECT 311.955 -140.925 312.285 -140.595 ;
        RECT 311.955 -142.285 312.285 -141.955 ;
        RECT 311.955 -143.645 312.285 -143.315 ;
        RECT 311.955 -145.005 312.285 -144.675 ;
        RECT 311.955 -146.365 312.285 -146.035 ;
        RECT 311.955 -147.725 312.285 -147.395 ;
        RECT 311.955 -149.085 312.285 -148.755 ;
        RECT 311.955 -150.445 312.285 -150.115 ;
        RECT 311.955 -151.805 312.285 -151.475 ;
        RECT 311.955 -153.165 312.285 -152.835 ;
        RECT 311.955 -154.525 312.285 -154.195 ;
        RECT 311.955 -155.885 312.285 -155.555 ;
        RECT 311.955 -157.245 312.285 -156.915 ;
        RECT 311.955 -158.605 312.285 -158.275 ;
        RECT 311.955 -159.965 312.285 -159.635 ;
        RECT 311.955 -161.325 312.285 -160.995 ;
        RECT 311.955 -162.685 312.285 -162.355 ;
        RECT 311.955 -164.045 312.285 -163.715 ;
        RECT 311.955 -165.405 312.285 -165.075 ;
        RECT 311.955 -166.765 312.285 -166.435 ;
        RECT 311.955 -168.125 312.285 -167.795 ;
        RECT 311.955 -169.485 312.285 -169.155 ;
        RECT 311.955 -170.845 312.285 -170.515 ;
        RECT 311.955 -172.205 312.285 -171.875 ;
        RECT 311.955 -173.565 312.285 -173.235 ;
        RECT 311.955 -174.925 312.285 -174.595 ;
        RECT 311.955 -176.285 312.285 -175.955 ;
        RECT 311.955 -177.645 312.285 -177.315 ;
        RECT 311.955 -183.29 312.285 -182.16 ;
        RECT 311.96 -183.405 312.28 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 313.315 244.04 313.645 245.17 ;
        RECT 313.315 239.875 313.645 240.205 ;
        RECT 313.315 238.515 313.645 238.845 ;
        RECT 313.315 237.155 313.645 237.485 ;
        RECT 313.32 237.155 313.64 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 313.315 -96.045 313.645 -95.715 ;
        RECT 313.315 -97.405 313.645 -97.075 ;
        RECT 313.315 -98.765 313.645 -98.435 ;
        RECT 313.315 -100.125 313.645 -99.795 ;
        RECT 313.315 -101.485 313.645 -101.155 ;
        RECT 313.315 -102.845 313.645 -102.515 ;
        RECT 313.315 -104.205 313.645 -103.875 ;
        RECT 313.315 -105.565 313.645 -105.235 ;
        RECT 313.315 -106.925 313.645 -106.595 ;
        RECT 313.315 -108.285 313.645 -107.955 ;
        RECT 313.315 -109.645 313.645 -109.315 ;
        RECT 313.315 -111.005 313.645 -110.675 ;
        RECT 313.315 -112.365 313.645 -112.035 ;
        RECT 313.315 -113.725 313.645 -113.395 ;
        RECT 313.315 -115.085 313.645 -114.755 ;
        RECT 313.315 -116.445 313.645 -116.115 ;
        RECT 313.315 -117.805 313.645 -117.475 ;
        RECT 313.315 -119.165 313.645 -118.835 ;
        RECT 313.315 -120.525 313.645 -120.195 ;
        RECT 313.315 -121.885 313.645 -121.555 ;
        RECT 313.315 -123.245 313.645 -122.915 ;
        RECT 313.315 -124.605 313.645 -124.275 ;
        RECT 313.315 -125.965 313.645 -125.635 ;
        RECT 313.315 -127.325 313.645 -126.995 ;
        RECT 313.315 -128.685 313.645 -128.355 ;
        RECT 313.315 -130.045 313.645 -129.715 ;
        RECT 313.315 -131.405 313.645 -131.075 ;
        RECT 313.315 -132.765 313.645 -132.435 ;
        RECT 313.315 -134.125 313.645 -133.795 ;
        RECT 313.315 -135.485 313.645 -135.155 ;
        RECT 313.315 -136.845 313.645 -136.515 ;
        RECT 313.315 -138.205 313.645 -137.875 ;
        RECT 313.315 -139.565 313.645 -139.235 ;
        RECT 313.315 -140.925 313.645 -140.595 ;
        RECT 313.315 -142.285 313.645 -141.955 ;
        RECT 313.315 -143.645 313.645 -143.315 ;
        RECT 313.315 -145.005 313.645 -144.675 ;
        RECT 313.315 -146.365 313.645 -146.035 ;
        RECT 313.315 -147.725 313.645 -147.395 ;
        RECT 313.315 -149.085 313.645 -148.755 ;
        RECT 313.315 -150.445 313.645 -150.115 ;
        RECT 313.315 -151.805 313.645 -151.475 ;
        RECT 313.315 -153.165 313.645 -152.835 ;
        RECT 313.315 -154.525 313.645 -154.195 ;
        RECT 313.315 -155.885 313.645 -155.555 ;
        RECT 313.315 -157.245 313.645 -156.915 ;
        RECT 313.315 -158.605 313.645 -158.275 ;
        RECT 313.315 -159.965 313.645 -159.635 ;
        RECT 313.315 -161.325 313.645 -160.995 ;
        RECT 313.315 -162.685 313.645 -162.355 ;
        RECT 313.315 -164.045 313.645 -163.715 ;
        RECT 313.315 -165.405 313.645 -165.075 ;
        RECT 313.315 -166.765 313.645 -166.435 ;
        RECT 313.315 -168.125 313.645 -167.795 ;
        RECT 313.315 -169.485 313.645 -169.155 ;
        RECT 313.315 -170.845 313.645 -170.515 ;
        RECT 313.315 -172.205 313.645 -171.875 ;
        RECT 313.315 -173.565 313.645 -173.235 ;
        RECT 313.315 -174.925 313.645 -174.595 ;
        RECT 313.315 -176.285 313.645 -175.955 ;
        RECT 313.315 -177.645 313.645 -177.315 ;
        RECT 313.315 -183.29 313.645 -182.16 ;
        RECT 313.32 -183.405 313.64 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 313.76 -94.075 314.09 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 314.675 244.04 315.005 245.17 ;
        RECT 314.675 239.875 315.005 240.205 ;
        RECT 314.675 238.515 315.005 238.845 ;
        RECT 314.675 237.155 315.005 237.485 ;
        RECT 314.68 237.155 315 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 316.035 244.04 316.365 245.17 ;
        RECT 316.035 239.875 316.365 240.205 ;
        RECT 316.035 238.515 316.365 238.845 ;
        RECT 316.035 237.155 316.365 237.485 ;
        RECT 316.04 237.155 316.36 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 316.035 -0.845 316.365 -0.515 ;
        RECT 316.035 -2.205 316.365 -1.875 ;
        RECT 316.035 -3.565 316.365 -3.235 ;
        RECT 316.04 -3.565 316.36 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 317.395 244.04 317.725 245.17 ;
        RECT 317.395 239.875 317.725 240.205 ;
        RECT 317.395 238.515 317.725 238.845 ;
        RECT 317.395 237.155 317.725 237.485 ;
        RECT 317.4 237.155 317.72 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 317.395 -0.845 317.725 -0.515 ;
        RECT 317.395 -2.205 317.725 -1.875 ;
        RECT 317.395 -3.565 317.725 -3.235 ;
        RECT 317.4 -3.565 317.72 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 318.755 244.04 319.085 245.17 ;
        RECT 318.755 239.875 319.085 240.205 ;
        RECT 318.755 238.515 319.085 238.845 ;
        RECT 318.755 237.155 319.085 237.485 ;
        RECT 318.76 237.155 319.08 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 318.755 -0.845 319.085 -0.515 ;
        RECT 318.755 -2.205 319.085 -1.875 ;
        RECT 318.755 -3.565 319.085 -3.235 ;
        RECT 318.76 -3.565 319.08 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 318.755 -91.965 319.085 -91.635 ;
        RECT 318.755 -93.325 319.085 -92.995 ;
        RECT 318.755 -94.685 319.085 -94.355 ;
        RECT 318.755 -96.045 319.085 -95.715 ;
        RECT 318.755 -97.405 319.085 -97.075 ;
        RECT 318.755 -98.765 319.085 -98.435 ;
        RECT 318.755 -100.125 319.085 -99.795 ;
        RECT 318.755 -101.485 319.085 -101.155 ;
        RECT 318.755 -102.845 319.085 -102.515 ;
        RECT 318.755 -104.205 319.085 -103.875 ;
        RECT 318.755 -105.565 319.085 -105.235 ;
        RECT 318.755 -106.925 319.085 -106.595 ;
        RECT 318.755 -108.285 319.085 -107.955 ;
        RECT 318.755 -109.645 319.085 -109.315 ;
        RECT 318.755 -111.005 319.085 -110.675 ;
        RECT 318.755 -112.365 319.085 -112.035 ;
        RECT 318.755 -113.725 319.085 -113.395 ;
        RECT 318.755 -115.085 319.085 -114.755 ;
        RECT 318.755 -116.445 319.085 -116.115 ;
        RECT 318.755 -117.805 319.085 -117.475 ;
        RECT 318.755 -119.165 319.085 -118.835 ;
        RECT 318.755 -120.525 319.085 -120.195 ;
        RECT 318.755 -121.885 319.085 -121.555 ;
        RECT 318.755 -123.245 319.085 -122.915 ;
        RECT 318.755 -124.605 319.085 -124.275 ;
        RECT 318.755 -125.965 319.085 -125.635 ;
        RECT 318.755 -127.325 319.085 -126.995 ;
        RECT 318.755 -128.685 319.085 -128.355 ;
        RECT 318.755 -130.045 319.085 -129.715 ;
        RECT 318.755 -131.405 319.085 -131.075 ;
        RECT 318.755 -132.765 319.085 -132.435 ;
        RECT 318.755 -134.125 319.085 -133.795 ;
        RECT 318.755 -135.485 319.085 -135.155 ;
        RECT 318.755 -136.845 319.085 -136.515 ;
        RECT 318.755 -138.205 319.085 -137.875 ;
        RECT 318.755 -139.565 319.085 -139.235 ;
        RECT 318.755 -140.925 319.085 -140.595 ;
        RECT 318.755 -142.285 319.085 -141.955 ;
        RECT 318.755 -143.645 319.085 -143.315 ;
        RECT 318.755 -145.005 319.085 -144.675 ;
        RECT 318.755 -146.365 319.085 -146.035 ;
        RECT 318.755 -147.725 319.085 -147.395 ;
        RECT 318.755 -149.085 319.085 -148.755 ;
        RECT 318.755 -150.445 319.085 -150.115 ;
        RECT 318.755 -151.805 319.085 -151.475 ;
        RECT 318.755 -153.165 319.085 -152.835 ;
        RECT 318.755 -154.525 319.085 -154.195 ;
        RECT 318.755 -155.885 319.085 -155.555 ;
        RECT 318.755 -157.245 319.085 -156.915 ;
        RECT 318.755 -158.605 319.085 -158.275 ;
        RECT 318.755 -159.965 319.085 -159.635 ;
        RECT 318.755 -161.325 319.085 -160.995 ;
        RECT 318.755 -162.685 319.085 -162.355 ;
        RECT 318.755 -164.045 319.085 -163.715 ;
        RECT 318.755 -165.405 319.085 -165.075 ;
        RECT 318.755 -166.765 319.085 -166.435 ;
        RECT 318.755 -168.125 319.085 -167.795 ;
        RECT 318.755 -169.485 319.085 -169.155 ;
        RECT 318.755 -170.845 319.085 -170.515 ;
        RECT 318.755 -172.205 319.085 -171.875 ;
        RECT 318.755 -173.565 319.085 -173.235 ;
        RECT 318.755 -174.925 319.085 -174.595 ;
        RECT 318.755 -176.285 319.085 -175.955 ;
        RECT 318.755 -177.645 319.085 -177.315 ;
        RECT 318.755 -183.29 319.085 -182.16 ;
        RECT 318.76 -183.405 319.08 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 319.86 -94.075 320.19 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 320.115 244.04 320.445 245.17 ;
        RECT 320.115 239.875 320.445 240.205 ;
        RECT 320.115 238.515 320.445 238.845 ;
        RECT 320.115 237.155 320.445 237.485 ;
        RECT 320.12 237.155 320.44 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 320.115 -96.045 320.445 -95.715 ;
        RECT 320.115 -97.405 320.445 -97.075 ;
        RECT 320.115 -98.765 320.445 -98.435 ;
        RECT 320.115 -100.125 320.445 -99.795 ;
        RECT 320.115 -101.485 320.445 -101.155 ;
        RECT 320.115 -102.845 320.445 -102.515 ;
        RECT 320.115 -104.205 320.445 -103.875 ;
        RECT 320.115 -105.565 320.445 -105.235 ;
        RECT 320.115 -106.925 320.445 -106.595 ;
        RECT 320.115 -108.285 320.445 -107.955 ;
        RECT 320.115 -109.645 320.445 -109.315 ;
        RECT 320.115 -111.005 320.445 -110.675 ;
        RECT 320.115 -112.365 320.445 -112.035 ;
        RECT 320.115 -113.725 320.445 -113.395 ;
        RECT 320.115 -115.085 320.445 -114.755 ;
        RECT 320.115 -116.445 320.445 -116.115 ;
        RECT 320.115 -117.805 320.445 -117.475 ;
        RECT 320.115 -119.165 320.445 -118.835 ;
        RECT 320.115 -120.525 320.445 -120.195 ;
        RECT 320.115 -121.885 320.445 -121.555 ;
        RECT 320.115 -123.245 320.445 -122.915 ;
        RECT 320.115 -124.605 320.445 -124.275 ;
        RECT 320.115 -125.965 320.445 -125.635 ;
        RECT 320.115 -127.325 320.445 -126.995 ;
        RECT 320.115 -128.685 320.445 -128.355 ;
        RECT 320.115 -130.045 320.445 -129.715 ;
        RECT 320.115 -131.405 320.445 -131.075 ;
        RECT 320.115 -132.765 320.445 -132.435 ;
        RECT 320.115 -134.125 320.445 -133.795 ;
        RECT 320.115 -135.485 320.445 -135.155 ;
        RECT 320.115 -136.845 320.445 -136.515 ;
        RECT 320.115 -138.205 320.445 -137.875 ;
        RECT 320.115 -139.565 320.445 -139.235 ;
        RECT 320.115 -140.925 320.445 -140.595 ;
        RECT 320.115 -142.285 320.445 -141.955 ;
        RECT 320.115 -143.645 320.445 -143.315 ;
        RECT 320.115 -145.005 320.445 -144.675 ;
        RECT 320.115 -146.365 320.445 -146.035 ;
        RECT 320.115 -147.725 320.445 -147.395 ;
        RECT 320.115 -149.085 320.445 -148.755 ;
        RECT 320.115 -150.445 320.445 -150.115 ;
        RECT 320.115 -151.805 320.445 -151.475 ;
        RECT 320.115 -153.165 320.445 -152.835 ;
        RECT 320.115 -154.525 320.445 -154.195 ;
        RECT 320.115 -155.885 320.445 -155.555 ;
        RECT 320.115 -157.245 320.445 -156.915 ;
        RECT 320.115 -158.605 320.445 -158.275 ;
        RECT 320.115 -159.965 320.445 -159.635 ;
        RECT 320.115 -161.325 320.445 -160.995 ;
        RECT 320.115 -162.685 320.445 -162.355 ;
        RECT 320.115 -164.045 320.445 -163.715 ;
        RECT 320.115 -165.405 320.445 -165.075 ;
        RECT 320.115 -166.765 320.445 -166.435 ;
        RECT 320.115 -168.125 320.445 -167.795 ;
        RECT 320.115 -169.485 320.445 -169.155 ;
        RECT 320.115 -170.845 320.445 -170.515 ;
        RECT 320.115 -172.205 320.445 -171.875 ;
        RECT 320.115 -173.565 320.445 -173.235 ;
        RECT 320.115 -174.925 320.445 -174.595 ;
        RECT 320.115 -176.285 320.445 -175.955 ;
        RECT 320.115 -177.645 320.445 -177.315 ;
        RECT 320.115 -183.29 320.445 -182.16 ;
        RECT 320.12 -183.405 320.44 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 321.475 244.04 321.805 245.17 ;
        RECT 321.475 239.875 321.805 240.205 ;
        RECT 321.475 238.515 321.805 238.845 ;
        RECT 321.475 237.155 321.805 237.485 ;
        RECT 321.48 237.155 321.8 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 321.475 -0.845 321.805 -0.515 ;
        RECT 321.475 -2.205 321.805 -1.875 ;
        RECT 321.475 -3.565 321.805 -3.235 ;
        RECT 321.48 -3.565 321.8 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 322.835 244.04 323.165 245.17 ;
        RECT 322.835 239.875 323.165 240.205 ;
        RECT 322.835 238.515 323.165 238.845 ;
        RECT 322.835 237.155 323.165 237.485 ;
        RECT 322.84 237.155 323.16 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 322.835 -0.845 323.165 -0.515 ;
        RECT 322.835 -2.205 323.165 -1.875 ;
        RECT 322.835 -3.565 323.165 -3.235 ;
        RECT 322.84 -3.565 323.16 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 324.195 244.04 324.525 245.17 ;
        RECT 324.195 239.875 324.525 240.205 ;
        RECT 324.195 238.515 324.525 238.845 ;
        RECT 324.195 237.155 324.525 237.485 ;
        RECT 324.2 237.155 324.52 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 324.195 -0.845 324.525 -0.515 ;
        RECT 324.195 -2.205 324.525 -1.875 ;
        RECT 324.195 -3.565 324.525 -3.235 ;
        RECT 324.2 -3.565 324.52 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 324.195 -91.965 324.525 -91.635 ;
        RECT 324.195 -93.325 324.525 -92.995 ;
        RECT 324.195 -94.685 324.525 -94.355 ;
        RECT 324.195 -96.045 324.525 -95.715 ;
        RECT 324.195 -97.405 324.525 -97.075 ;
        RECT 324.195 -98.765 324.525 -98.435 ;
        RECT 324.195 -100.125 324.525 -99.795 ;
        RECT 324.195 -101.485 324.525 -101.155 ;
        RECT 324.195 -102.845 324.525 -102.515 ;
        RECT 324.195 -104.205 324.525 -103.875 ;
        RECT 324.195 -105.565 324.525 -105.235 ;
        RECT 324.195 -106.925 324.525 -106.595 ;
        RECT 324.195 -108.285 324.525 -107.955 ;
        RECT 324.195 -109.645 324.525 -109.315 ;
        RECT 324.195 -111.005 324.525 -110.675 ;
        RECT 324.195 -112.365 324.525 -112.035 ;
        RECT 324.195 -113.725 324.525 -113.395 ;
        RECT 324.195 -115.085 324.525 -114.755 ;
        RECT 324.195 -116.445 324.525 -116.115 ;
        RECT 324.195 -117.805 324.525 -117.475 ;
        RECT 324.195 -119.165 324.525 -118.835 ;
        RECT 324.195 -120.525 324.525 -120.195 ;
        RECT 324.195 -121.885 324.525 -121.555 ;
        RECT 324.195 -123.245 324.525 -122.915 ;
        RECT 324.195 -124.605 324.525 -124.275 ;
        RECT 324.195 -125.965 324.525 -125.635 ;
        RECT 324.195 -127.325 324.525 -126.995 ;
        RECT 324.195 -128.685 324.525 -128.355 ;
        RECT 324.195 -130.045 324.525 -129.715 ;
        RECT 324.195 -131.405 324.525 -131.075 ;
        RECT 324.195 -132.765 324.525 -132.435 ;
        RECT 324.195 -134.125 324.525 -133.795 ;
        RECT 324.195 -135.485 324.525 -135.155 ;
        RECT 324.195 -136.845 324.525 -136.515 ;
        RECT 324.195 -138.205 324.525 -137.875 ;
        RECT 324.195 -139.565 324.525 -139.235 ;
        RECT 324.195 -140.925 324.525 -140.595 ;
        RECT 324.195 -142.285 324.525 -141.955 ;
        RECT 324.195 -143.645 324.525 -143.315 ;
        RECT 324.195 -145.005 324.525 -144.675 ;
        RECT 324.195 -146.365 324.525 -146.035 ;
        RECT 324.195 -147.725 324.525 -147.395 ;
        RECT 324.195 -149.085 324.525 -148.755 ;
        RECT 324.195 -150.445 324.525 -150.115 ;
        RECT 324.195 -151.805 324.525 -151.475 ;
        RECT 324.195 -153.165 324.525 -152.835 ;
        RECT 324.195 -154.525 324.525 -154.195 ;
        RECT 324.195 -155.885 324.525 -155.555 ;
        RECT 324.195 -157.245 324.525 -156.915 ;
        RECT 324.195 -158.605 324.525 -158.275 ;
        RECT 324.195 -159.965 324.525 -159.635 ;
        RECT 324.195 -161.325 324.525 -160.995 ;
        RECT 324.195 -162.685 324.525 -162.355 ;
        RECT 324.195 -164.045 324.525 -163.715 ;
        RECT 324.195 -165.405 324.525 -165.075 ;
        RECT 324.195 -166.765 324.525 -166.435 ;
        RECT 324.195 -168.125 324.525 -167.795 ;
        RECT 324.195 -169.485 324.525 -169.155 ;
        RECT 324.195 -170.845 324.525 -170.515 ;
        RECT 324.195 -172.205 324.525 -171.875 ;
        RECT 324.195 -173.565 324.525 -173.235 ;
        RECT 324.195 -174.925 324.525 -174.595 ;
        RECT 324.195 -176.285 324.525 -175.955 ;
        RECT 324.195 -177.645 324.525 -177.315 ;
        RECT 324.195 -183.29 324.525 -182.16 ;
        RECT 324.2 -183.405 324.52 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 325.555 244.04 325.885 245.17 ;
        RECT 325.555 239.875 325.885 240.205 ;
        RECT 325.555 238.515 325.885 238.845 ;
        RECT 325.555 237.155 325.885 237.485 ;
        RECT 325.56 237.155 325.88 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 325.555 -96.045 325.885 -95.715 ;
        RECT 325.555 -97.405 325.885 -97.075 ;
        RECT 325.555 -98.765 325.885 -98.435 ;
        RECT 325.555 -100.125 325.885 -99.795 ;
        RECT 325.555 -101.485 325.885 -101.155 ;
        RECT 325.555 -102.845 325.885 -102.515 ;
        RECT 325.555 -104.205 325.885 -103.875 ;
        RECT 325.555 -105.565 325.885 -105.235 ;
        RECT 325.555 -106.925 325.885 -106.595 ;
        RECT 325.555 -108.285 325.885 -107.955 ;
        RECT 325.555 -109.645 325.885 -109.315 ;
        RECT 325.555 -111.005 325.885 -110.675 ;
        RECT 325.555 -112.365 325.885 -112.035 ;
        RECT 325.555 -113.725 325.885 -113.395 ;
        RECT 325.555 -115.085 325.885 -114.755 ;
        RECT 325.555 -116.445 325.885 -116.115 ;
        RECT 325.555 -117.805 325.885 -117.475 ;
        RECT 325.555 -119.165 325.885 -118.835 ;
        RECT 325.555 -120.525 325.885 -120.195 ;
        RECT 325.555 -121.885 325.885 -121.555 ;
        RECT 325.555 -123.245 325.885 -122.915 ;
        RECT 325.555 -124.605 325.885 -124.275 ;
        RECT 325.555 -125.965 325.885 -125.635 ;
        RECT 325.555 -127.325 325.885 -126.995 ;
        RECT 325.555 -128.685 325.885 -128.355 ;
        RECT 325.555 -130.045 325.885 -129.715 ;
        RECT 325.555 -131.405 325.885 -131.075 ;
        RECT 325.555 -132.765 325.885 -132.435 ;
        RECT 325.555 -134.125 325.885 -133.795 ;
        RECT 325.555 -135.485 325.885 -135.155 ;
        RECT 325.555 -136.845 325.885 -136.515 ;
        RECT 325.555 -138.205 325.885 -137.875 ;
        RECT 325.555 -139.565 325.885 -139.235 ;
        RECT 325.555 -140.925 325.885 -140.595 ;
        RECT 325.555 -142.285 325.885 -141.955 ;
        RECT 325.555 -143.645 325.885 -143.315 ;
        RECT 325.555 -145.005 325.885 -144.675 ;
        RECT 325.555 -146.365 325.885 -146.035 ;
        RECT 325.555 -147.725 325.885 -147.395 ;
        RECT 325.555 -149.085 325.885 -148.755 ;
        RECT 325.555 -150.445 325.885 -150.115 ;
        RECT 325.555 -151.805 325.885 -151.475 ;
        RECT 325.555 -153.165 325.885 -152.835 ;
        RECT 325.555 -154.525 325.885 -154.195 ;
        RECT 325.555 -155.885 325.885 -155.555 ;
        RECT 325.555 -157.245 325.885 -156.915 ;
        RECT 325.555 -158.605 325.885 -158.275 ;
        RECT 325.555 -159.965 325.885 -159.635 ;
        RECT 325.555 -161.325 325.885 -160.995 ;
        RECT 325.555 -162.685 325.885 -162.355 ;
        RECT 325.555 -164.045 325.885 -163.715 ;
        RECT 325.555 -165.405 325.885 -165.075 ;
        RECT 325.555 -166.765 325.885 -166.435 ;
        RECT 325.555 -168.125 325.885 -167.795 ;
        RECT 325.555 -169.485 325.885 -169.155 ;
        RECT 325.555 -170.845 325.885 -170.515 ;
        RECT 325.555 -172.205 325.885 -171.875 ;
        RECT 325.555 -173.565 325.885 -173.235 ;
        RECT 325.555 -174.925 325.885 -174.595 ;
        RECT 325.555 -176.285 325.885 -175.955 ;
        RECT 325.555 -177.645 325.885 -177.315 ;
        RECT 325.555 -183.29 325.885 -182.16 ;
        RECT 325.56 -183.405 325.88 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 325.96 -94.075 326.29 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 326.915 244.04 327.245 245.17 ;
        RECT 326.915 239.875 327.245 240.205 ;
        RECT 326.915 238.515 327.245 238.845 ;
        RECT 326.915 237.155 327.245 237.485 ;
        RECT 326.92 237.155 327.24 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 328.275 244.04 328.605 245.17 ;
        RECT 328.275 239.875 328.605 240.205 ;
        RECT 328.275 238.515 328.605 238.845 ;
        RECT 328.275 237.155 328.605 237.485 ;
        RECT 328.28 237.155 328.6 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 328.275 -0.845 328.605 -0.515 ;
        RECT 328.275 -2.205 328.605 -1.875 ;
        RECT 328.275 -3.565 328.605 -3.235 ;
        RECT 328.28 -3.565 328.6 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 329.635 244.04 329.965 245.17 ;
        RECT 329.635 239.875 329.965 240.205 ;
        RECT 329.635 238.515 329.965 238.845 ;
        RECT 329.635 237.155 329.965 237.485 ;
        RECT 329.64 237.155 329.96 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 329.635 -0.845 329.965 -0.515 ;
        RECT 329.635 -2.205 329.965 -1.875 ;
        RECT 329.635 -3.565 329.965 -3.235 ;
        RECT 329.64 -3.565 329.96 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 330.995 244.04 331.325 245.17 ;
        RECT 330.995 239.875 331.325 240.205 ;
        RECT 330.995 238.515 331.325 238.845 ;
        RECT 330.995 237.155 331.325 237.485 ;
        RECT 331 237.155 331.32 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 330.995 -0.845 331.325 -0.515 ;
        RECT 330.995 -2.205 331.325 -1.875 ;
        RECT 330.995 -3.565 331.325 -3.235 ;
        RECT 331 -3.565 331.32 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 330.995 -91.965 331.325 -91.635 ;
        RECT 330.995 -93.325 331.325 -92.995 ;
        RECT 330.995 -94.685 331.325 -94.355 ;
        RECT 330.995 -96.045 331.325 -95.715 ;
        RECT 330.995 -97.405 331.325 -97.075 ;
        RECT 330.995 -98.765 331.325 -98.435 ;
        RECT 330.995 -100.125 331.325 -99.795 ;
        RECT 330.995 -101.485 331.325 -101.155 ;
        RECT 330.995 -102.845 331.325 -102.515 ;
        RECT 330.995 -104.205 331.325 -103.875 ;
        RECT 330.995 -105.565 331.325 -105.235 ;
        RECT 330.995 -106.925 331.325 -106.595 ;
        RECT 330.995 -108.285 331.325 -107.955 ;
        RECT 330.995 -109.645 331.325 -109.315 ;
        RECT 330.995 -111.005 331.325 -110.675 ;
        RECT 330.995 -112.365 331.325 -112.035 ;
        RECT 330.995 -113.725 331.325 -113.395 ;
        RECT 330.995 -115.085 331.325 -114.755 ;
        RECT 330.995 -116.445 331.325 -116.115 ;
        RECT 330.995 -117.805 331.325 -117.475 ;
        RECT 330.995 -119.165 331.325 -118.835 ;
        RECT 330.995 -120.525 331.325 -120.195 ;
        RECT 330.995 -121.885 331.325 -121.555 ;
        RECT 330.995 -123.245 331.325 -122.915 ;
        RECT 330.995 -124.605 331.325 -124.275 ;
        RECT 330.995 -125.965 331.325 -125.635 ;
        RECT 330.995 -127.325 331.325 -126.995 ;
        RECT 330.995 -128.685 331.325 -128.355 ;
        RECT 330.995 -130.045 331.325 -129.715 ;
        RECT 330.995 -131.405 331.325 -131.075 ;
        RECT 330.995 -132.765 331.325 -132.435 ;
        RECT 330.995 -134.125 331.325 -133.795 ;
        RECT 330.995 -135.485 331.325 -135.155 ;
        RECT 330.995 -136.845 331.325 -136.515 ;
        RECT 330.995 -138.205 331.325 -137.875 ;
        RECT 330.995 -139.565 331.325 -139.235 ;
        RECT 330.995 -140.925 331.325 -140.595 ;
        RECT 330.995 -142.285 331.325 -141.955 ;
        RECT 330.995 -143.645 331.325 -143.315 ;
        RECT 330.995 -145.005 331.325 -144.675 ;
        RECT 330.995 -146.365 331.325 -146.035 ;
        RECT 330.995 -147.725 331.325 -147.395 ;
        RECT 330.995 -149.085 331.325 -148.755 ;
        RECT 330.995 -150.445 331.325 -150.115 ;
        RECT 330.995 -151.805 331.325 -151.475 ;
        RECT 330.995 -153.165 331.325 -152.835 ;
        RECT 330.995 -154.525 331.325 -154.195 ;
        RECT 330.995 -155.885 331.325 -155.555 ;
        RECT 330.995 -157.245 331.325 -156.915 ;
        RECT 330.995 -158.605 331.325 -158.275 ;
        RECT 330.995 -159.965 331.325 -159.635 ;
        RECT 330.995 -161.325 331.325 -160.995 ;
        RECT 330.995 -162.685 331.325 -162.355 ;
        RECT 330.995 -164.045 331.325 -163.715 ;
        RECT 330.995 -165.405 331.325 -165.075 ;
        RECT 330.995 -166.765 331.325 -166.435 ;
        RECT 330.995 -168.125 331.325 -167.795 ;
        RECT 330.995 -169.485 331.325 -169.155 ;
        RECT 330.995 -170.845 331.325 -170.515 ;
        RECT 330.995 -172.205 331.325 -171.875 ;
        RECT 330.995 -173.565 331.325 -173.235 ;
        RECT 330.995 -174.925 331.325 -174.595 ;
        RECT 330.995 -176.285 331.325 -175.955 ;
        RECT 330.995 -177.645 331.325 -177.315 ;
        RECT 330.995 -183.29 331.325 -182.16 ;
        RECT 331 -183.405 331.32 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 332.06 -94.075 332.39 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 332.355 244.04 332.685 245.17 ;
        RECT 332.355 239.875 332.685 240.205 ;
        RECT 332.355 238.515 332.685 238.845 ;
        RECT 332.355 237.155 332.685 237.485 ;
        RECT 332.36 237.155 332.68 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 332.355 -96.045 332.685 -95.715 ;
        RECT 332.355 -97.405 332.685 -97.075 ;
        RECT 332.355 -98.765 332.685 -98.435 ;
        RECT 332.355 -100.125 332.685 -99.795 ;
        RECT 332.355 -101.485 332.685 -101.155 ;
        RECT 332.355 -102.845 332.685 -102.515 ;
        RECT 332.355 -104.205 332.685 -103.875 ;
        RECT 332.355 -105.565 332.685 -105.235 ;
        RECT 332.355 -106.925 332.685 -106.595 ;
        RECT 332.355 -108.285 332.685 -107.955 ;
        RECT 332.355 -109.645 332.685 -109.315 ;
        RECT 332.355 -111.005 332.685 -110.675 ;
        RECT 332.355 -112.365 332.685 -112.035 ;
        RECT 332.355 -113.725 332.685 -113.395 ;
        RECT 332.355 -115.085 332.685 -114.755 ;
        RECT 332.355 -116.445 332.685 -116.115 ;
        RECT 332.355 -117.805 332.685 -117.475 ;
        RECT 332.355 -119.165 332.685 -118.835 ;
        RECT 332.355 -120.525 332.685 -120.195 ;
        RECT 332.355 -121.885 332.685 -121.555 ;
        RECT 332.355 -123.245 332.685 -122.915 ;
        RECT 332.355 -124.605 332.685 -124.275 ;
        RECT 332.355 -125.965 332.685 -125.635 ;
        RECT 332.355 -127.325 332.685 -126.995 ;
        RECT 332.355 -128.685 332.685 -128.355 ;
        RECT 332.355 -130.045 332.685 -129.715 ;
        RECT 332.355 -131.405 332.685 -131.075 ;
        RECT 332.355 -132.765 332.685 -132.435 ;
        RECT 332.355 -134.125 332.685 -133.795 ;
        RECT 332.355 -135.485 332.685 -135.155 ;
        RECT 332.355 -136.845 332.685 -136.515 ;
        RECT 332.355 -138.205 332.685 -137.875 ;
        RECT 332.355 -139.565 332.685 -139.235 ;
        RECT 332.355 -140.925 332.685 -140.595 ;
        RECT 332.355 -142.285 332.685 -141.955 ;
        RECT 332.355 -143.645 332.685 -143.315 ;
        RECT 332.355 -145.005 332.685 -144.675 ;
        RECT 332.355 -146.365 332.685 -146.035 ;
        RECT 332.355 -147.725 332.685 -147.395 ;
        RECT 332.355 -149.085 332.685 -148.755 ;
        RECT 332.355 -150.445 332.685 -150.115 ;
        RECT 332.355 -151.805 332.685 -151.475 ;
        RECT 332.355 -153.165 332.685 -152.835 ;
        RECT 332.355 -154.525 332.685 -154.195 ;
        RECT 332.355 -155.885 332.685 -155.555 ;
        RECT 332.355 -157.245 332.685 -156.915 ;
        RECT 332.355 -158.605 332.685 -158.275 ;
        RECT 332.355 -159.965 332.685 -159.635 ;
        RECT 332.355 -161.325 332.685 -160.995 ;
        RECT 332.355 -162.685 332.685 -162.355 ;
        RECT 332.355 -164.045 332.685 -163.715 ;
        RECT 332.355 -165.405 332.685 -165.075 ;
        RECT 332.355 -166.765 332.685 -166.435 ;
        RECT 332.355 -168.125 332.685 -167.795 ;
        RECT 332.355 -169.485 332.685 -169.155 ;
        RECT 332.355 -170.845 332.685 -170.515 ;
        RECT 332.355 -172.205 332.685 -171.875 ;
        RECT 332.355 -173.565 332.685 -173.235 ;
        RECT 332.355 -174.925 332.685 -174.595 ;
        RECT 332.355 -176.285 332.685 -175.955 ;
        RECT 332.355 -177.645 332.685 -177.315 ;
        RECT 332.355 -183.29 332.685 -182.16 ;
        RECT 332.36 -183.405 332.68 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 333.715 244.04 334.045 245.17 ;
        RECT 333.715 239.875 334.045 240.205 ;
        RECT 333.715 238.515 334.045 238.845 ;
        RECT 333.715 237.155 334.045 237.485 ;
        RECT 333.72 237.155 334.04 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 333.715 -0.845 334.045 -0.515 ;
        RECT 333.715 -2.205 334.045 -1.875 ;
        RECT 333.715 -3.565 334.045 -3.235 ;
        RECT 333.72 -3.565 334.04 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 335.075 244.04 335.405 245.17 ;
        RECT 335.075 239.875 335.405 240.205 ;
        RECT 335.075 238.515 335.405 238.845 ;
        RECT 335.075 237.155 335.405 237.485 ;
        RECT 335.08 237.155 335.4 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 335.075 -0.845 335.405 -0.515 ;
        RECT 335.075 -2.205 335.405 -1.875 ;
        RECT 335.075 -3.565 335.405 -3.235 ;
        RECT 335.08 -3.565 335.4 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 336.435 244.04 336.765 245.17 ;
        RECT 336.435 239.875 336.765 240.205 ;
        RECT 336.435 238.515 336.765 238.845 ;
        RECT 336.435 237.155 336.765 237.485 ;
        RECT 336.44 237.155 336.76 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 336.435 -0.845 336.765 -0.515 ;
        RECT 336.435 -2.205 336.765 -1.875 ;
        RECT 336.435 -3.565 336.765 -3.235 ;
        RECT 336.44 -3.565 336.76 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 336.435 -91.965 336.765 -91.635 ;
        RECT 336.435 -93.325 336.765 -92.995 ;
        RECT 336.435 -94.685 336.765 -94.355 ;
        RECT 336.435 -96.045 336.765 -95.715 ;
        RECT 336.435 -97.405 336.765 -97.075 ;
        RECT 336.435 -98.765 336.765 -98.435 ;
        RECT 336.435 -100.125 336.765 -99.795 ;
        RECT 336.435 -101.485 336.765 -101.155 ;
        RECT 336.435 -102.845 336.765 -102.515 ;
        RECT 336.435 -104.205 336.765 -103.875 ;
        RECT 336.435 -105.565 336.765 -105.235 ;
        RECT 336.435 -106.925 336.765 -106.595 ;
        RECT 336.435 -108.285 336.765 -107.955 ;
        RECT 336.435 -109.645 336.765 -109.315 ;
        RECT 336.435 -111.005 336.765 -110.675 ;
        RECT 336.435 -112.365 336.765 -112.035 ;
        RECT 336.435 -113.725 336.765 -113.395 ;
        RECT 336.435 -115.085 336.765 -114.755 ;
        RECT 336.435 -116.445 336.765 -116.115 ;
        RECT 336.435 -117.805 336.765 -117.475 ;
        RECT 336.435 -119.165 336.765 -118.835 ;
        RECT 336.435 -120.525 336.765 -120.195 ;
        RECT 336.435 -121.885 336.765 -121.555 ;
        RECT 336.435 -123.245 336.765 -122.915 ;
        RECT 336.435 -124.605 336.765 -124.275 ;
        RECT 336.435 -125.965 336.765 -125.635 ;
        RECT 336.435 -127.325 336.765 -126.995 ;
        RECT 336.435 -128.685 336.765 -128.355 ;
        RECT 336.435 -130.045 336.765 -129.715 ;
        RECT 336.435 -131.405 336.765 -131.075 ;
        RECT 336.435 -132.765 336.765 -132.435 ;
        RECT 336.435 -134.125 336.765 -133.795 ;
        RECT 336.435 -135.485 336.765 -135.155 ;
        RECT 336.435 -136.845 336.765 -136.515 ;
        RECT 336.435 -138.205 336.765 -137.875 ;
        RECT 336.435 -139.565 336.765 -139.235 ;
        RECT 336.435 -140.925 336.765 -140.595 ;
        RECT 336.435 -142.285 336.765 -141.955 ;
        RECT 336.435 -143.645 336.765 -143.315 ;
        RECT 336.435 -145.005 336.765 -144.675 ;
        RECT 336.435 -146.365 336.765 -146.035 ;
        RECT 336.435 -147.725 336.765 -147.395 ;
        RECT 336.435 -149.085 336.765 -148.755 ;
        RECT 336.435 -150.445 336.765 -150.115 ;
        RECT 336.435 -151.805 336.765 -151.475 ;
        RECT 336.435 -153.165 336.765 -152.835 ;
        RECT 336.435 -154.525 336.765 -154.195 ;
        RECT 336.435 -155.885 336.765 -155.555 ;
        RECT 336.435 -157.245 336.765 -156.915 ;
        RECT 336.435 -158.605 336.765 -158.275 ;
        RECT 336.435 -159.965 336.765 -159.635 ;
        RECT 336.435 -161.325 336.765 -160.995 ;
        RECT 336.435 -162.685 336.765 -162.355 ;
        RECT 336.435 -164.045 336.765 -163.715 ;
        RECT 336.435 -165.405 336.765 -165.075 ;
        RECT 336.435 -166.765 336.765 -166.435 ;
        RECT 336.435 -168.125 336.765 -167.795 ;
        RECT 336.435 -169.485 336.765 -169.155 ;
        RECT 336.435 -170.845 336.765 -170.515 ;
        RECT 336.435 -172.205 336.765 -171.875 ;
        RECT 336.435 -173.565 336.765 -173.235 ;
        RECT 336.435 -174.925 336.765 -174.595 ;
        RECT 336.435 -176.285 336.765 -175.955 ;
        RECT 336.435 -177.645 336.765 -177.315 ;
        RECT 336.435 -183.29 336.765 -182.16 ;
        RECT 336.44 -183.405 336.76 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 337.795 244.04 338.125 245.17 ;
        RECT 337.795 239.875 338.125 240.205 ;
        RECT 337.795 238.515 338.125 238.845 ;
        RECT 337.795 237.155 338.125 237.485 ;
        RECT 337.8 237.155 338.12 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 337.795 -96.045 338.125 -95.715 ;
        RECT 337.795 -97.405 338.125 -97.075 ;
        RECT 337.795 -98.765 338.125 -98.435 ;
        RECT 337.795 -100.125 338.125 -99.795 ;
        RECT 337.795 -101.485 338.125 -101.155 ;
        RECT 337.795 -102.845 338.125 -102.515 ;
        RECT 337.795 -104.205 338.125 -103.875 ;
        RECT 337.795 -105.565 338.125 -105.235 ;
        RECT 337.795 -106.925 338.125 -106.595 ;
        RECT 337.795 -108.285 338.125 -107.955 ;
        RECT 337.795 -109.645 338.125 -109.315 ;
        RECT 337.795 -111.005 338.125 -110.675 ;
        RECT 337.795 -112.365 338.125 -112.035 ;
        RECT 337.795 -113.725 338.125 -113.395 ;
        RECT 337.795 -115.085 338.125 -114.755 ;
        RECT 337.795 -116.445 338.125 -116.115 ;
        RECT 337.795 -117.805 338.125 -117.475 ;
        RECT 337.795 -119.165 338.125 -118.835 ;
        RECT 337.795 -120.525 338.125 -120.195 ;
        RECT 337.795 -121.885 338.125 -121.555 ;
        RECT 337.795 -123.245 338.125 -122.915 ;
        RECT 337.795 -124.605 338.125 -124.275 ;
        RECT 337.795 -125.965 338.125 -125.635 ;
        RECT 337.795 -127.325 338.125 -126.995 ;
        RECT 337.795 -128.685 338.125 -128.355 ;
        RECT 337.795 -130.045 338.125 -129.715 ;
        RECT 337.795 -131.405 338.125 -131.075 ;
        RECT 337.795 -132.765 338.125 -132.435 ;
        RECT 337.795 -134.125 338.125 -133.795 ;
        RECT 337.795 -135.485 338.125 -135.155 ;
        RECT 337.795 -136.845 338.125 -136.515 ;
        RECT 337.795 -138.205 338.125 -137.875 ;
        RECT 337.795 -139.565 338.125 -139.235 ;
        RECT 337.795 -140.925 338.125 -140.595 ;
        RECT 337.795 -142.285 338.125 -141.955 ;
        RECT 337.795 -143.645 338.125 -143.315 ;
        RECT 337.795 -145.005 338.125 -144.675 ;
        RECT 337.795 -146.365 338.125 -146.035 ;
        RECT 337.795 -147.725 338.125 -147.395 ;
        RECT 337.795 -149.085 338.125 -148.755 ;
        RECT 337.795 -150.445 338.125 -150.115 ;
        RECT 337.795 -151.805 338.125 -151.475 ;
        RECT 337.795 -153.165 338.125 -152.835 ;
        RECT 337.795 -154.525 338.125 -154.195 ;
        RECT 337.795 -155.885 338.125 -155.555 ;
        RECT 337.795 -157.245 338.125 -156.915 ;
        RECT 337.795 -158.605 338.125 -158.275 ;
        RECT 337.795 -159.965 338.125 -159.635 ;
        RECT 337.795 -161.325 338.125 -160.995 ;
        RECT 337.795 -162.685 338.125 -162.355 ;
        RECT 337.795 -164.045 338.125 -163.715 ;
        RECT 337.795 -165.405 338.125 -165.075 ;
        RECT 337.795 -166.765 338.125 -166.435 ;
        RECT 337.795 -168.125 338.125 -167.795 ;
        RECT 337.795 -169.485 338.125 -169.155 ;
        RECT 337.795 -170.845 338.125 -170.515 ;
        RECT 337.795 -172.205 338.125 -171.875 ;
        RECT 337.795 -173.565 338.125 -173.235 ;
        RECT 337.795 -174.925 338.125 -174.595 ;
        RECT 337.795 -176.285 338.125 -175.955 ;
        RECT 337.795 -177.645 338.125 -177.315 ;
        RECT 337.795 -183.29 338.125 -182.16 ;
        RECT 337.8 -183.405 338.12 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 338.16 -94.075 338.49 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 339.155 244.04 339.485 245.17 ;
        RECT 339.155 239.875 339.485 240.205 ;
        RECT 339.155 238.515 339.485 238.845 ;
        RECT 339.155 237.155 339.485 237.485 ;
        RECT 339.16 237.155 339.48 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 340.515 244.04 340.845 245.17 ;
        RECT 340.515 239.875 340.845 240.205 ;
        RECT 340.515 238.515 340.845 238.845 ;
        RECT 340.515 237.155 340.845 237.485 ;
        RECT 340.52 237.155 340.84 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 340.515 -0.845 340.845 -0.515 ;
        RECT 340.515 -2.205 340.845 -1.875 ;
        RECT 340.515 -3.565 340.845 -3.235 ;
        RECT 340.52 -3.565 340.84 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 341.875 244.04 342.205 245.17 ;
        RECT 341.875 239.875 342.205 240.205 ;
        RECT 341.875 238.515 342.205 238.845 ;
        RECT 341.875 237.155 342.205 237.485 ;
        RECT 341.88 237.155 342.2 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 341.875 -0.845 342.205 -0.515 ;
        RECT 341.875 -2.205 342.205 -1.875 ;
        RECT 341.875 -3.565 342.205 -3.235 ;
        RECT 341.88 -3.565 342.2 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 341.875 -157.245 342.205 -156.915 ;
        RECT 341.875 -158.605 342.205 -158.275 ;
        RECT 341.875 -159.965 342.205 -159.635 ;
        RECT 341.875 -161.325 342.205 -160.995 ;
        RECT 341.875 -162.685 342.205 -162.355 ;
        RECT 341.875 -164.045 342.205 -163.715 ;
        RECT 341.875 -165.405 342.205 -165.075 ;
        RECT 341.875 -166.765 342.205 -166.435 ;
        RECT 341.875 -168.125 342.205 -167.795 ;
        RECT 341.875 -169.485 342.205 -169.155 ;
        RECT 341.875 -170.845 342.205 -170.515 ;
        RECT 341.875 -172.205 342.205 -171.875 ;
        RECT 341.875 -173.565 342.205 -173.235 ;
        RECT 341.875 -174.925 342.205 -174.595 ;
        RECT 341.875 -176.285 342.205 -175.955 ;
        RECT 341.875 -177.645 342.205 -177.315 ;
        RECT 341.875 -183.29 342.205 -182.16 ;
        RECT 341.88 -183.405 342.2 -90.96 ;
        RECT 341.875 -91.965 342.205 -91.635 ;
        RECT 341.875 -93.325 342.205 -92.995 ;
        RECT 341.875 -94.685 342.205 -94.355 ;
        RECT 341.875 -96.045 342.205 -95.715 ;
        RECT 341.875 -97.405 342.205 -97.075 ;
        RECT 341.875 -98.765 342.205 -98.435 ;
        RECT 341.875 -100.125 342.205 -99.795 ;
        RECT 341.875 -101.485 342.205 -101.155 ;
        RECT 341.875 -102.845 342.205 -102.515 ;
        RECT 341.875 -104.205 342.205 -103.875 ;
        RECT 341.875 -105.565 342.205 -105.235 ;
        RECT 341.875 -106.925 342.205 -106.595 ;
        RECT 341.875 -108.285 342.205 -107.955 ;
        RECT 341.875 -109.645 342.205 -109.315 ;
        RECT 341.875 -111.005 342.205 -110.675 ;
        RECT 341.875 -112.365 342.205 -112.035 ;
        RECT 341.875 -113.725 342.205 -113.395 ;
        RECT 341.875 -115.085 342.205 -114.755 ;
        RECT 341.875 -116.445 342.205 -116.115 ;
        RECT 341.875 -117.805 342.205 -117.475 ;
        RECT 341.875 -119.165 342.205 -118.835 ;
        RECT 341.875 -120.525 342.205 -120.195 ;
        RECT 341.875 -121.885 342.205 -121.555 ;
        RECT 341.875 -123.245 342.205 -122.915 ;
        RECT 341.875 -124.605 342.205 -124.275 ;
        RECT 341.875 -125.965 342.205 -125.635 ;
        RECT 341.875 -127.325 342.205 -126.995 ;
        RECT 341.875 -128.685 342.205 -128.355 ;
        RECT 341.875 -130.045 342.205 -129.715 ;
        RECT 341.875 -131.405 342.205 -131.075 ;
        RECT 341.875 -132.765 342.205 -132.435 ;
        RECT 341.875 -134.125 342.205 -133.795 ;
        RECT 341.875 -135.485 342.205 -135.155 ;
        RECT 341.875 -136.845 342.205 -136.515 ;
        RECT 341.875 -138.205 342.205 -137.875 ;
        RECT 341.875 -139.565 342.205 -139.235 ;
        RECT 341.875 -140.925 342.205 -140.595 ;
        RECT 341.875 -142.285 342.205 -141.955 ;
        RECT 341.875 -143.645 342.205 -143.315 ;
        RECT 341.875 -145.005 342.205 -144.675 ;
        RECT 341.875 -146.365 342.205 -146.035 ;
        RECT 341.875 -147.725 342.205 -147.395 ;
        RECT 341.875 -149.085 342.205 -148.755 ;
        RECT 341.875 -150.445 342.205 -150.115 ;
        RECT 341.875 -151.805 342.205 -151.475 ;
        RECT 341.875 -153.165 342.205 -152.835 ;
        RECT 341.875 -154.525 342.205 -154.195 ;
        RECT 341.875 -155.885 342.205 -155.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 272.515 244.04 272.845 245.17 ;
        RECT 272.515 239.875 272.845 240.205 ;
        RECT 272.515 238.515 272.845 238.845 ;
        RECT 272.515 237.155 272.845 237.485 ;
        RECT 272.52 237.155 272.84 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 272.515 -0.845 272.845 -0.515 ;
        RECT 272.515 -2.205 272.845 -1.875 ;
        RECT 272.515 -3.565 272.845 -3.235 ;
        RECT 272.52 -3.565 272.84 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 273.875 244.04 274.205 245.17 ;
        RECT 273.875 239.875 274.205 240.205 ;
        RECT 273.875 238.515 274.205 238.845 ;
        RECT 273.875 237.155 274.205 237.485 ;
        RECT 273.88 237.155 274.2 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 273.875 -0.845 274.205 -0.515 ;
        RECT 273.875 -2.205 274.205 -1.875 ;
        RECT 273.875 -3.565 274.205 -3.235 ;
        RECT 273.88 -3.565 274.2 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 275.235 244.04 275.565 245.17 ;
        RECT 275.235 239.875 275.565 240.205 ;
        RECT 275.235 238.515 275.565 238.845 ;
        RECT 275.235 237.155 275.565 237.485 ;
        RECT 275.24 237.155 275.56 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 275.235 -0.845 275.565 -0.515 ;
        RECT 275.235 -2.205 275.565 -1.875 ;
        RECT 275.235 -3.565 275.565 -3.235 ;
        RECT 275.24 -3.565 275.56 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 275.235 -91.965 275.565 -91.635 ;
        RECT 275.235 -93.325 275.565 -92.995 ;
        RECT 275.235 -94.685 275.565 -94.355 ;
        RECT 275.235 -96.045 275.565 -95.715 ;
        RECT 275.235 -97.405 275.565 -97.075 ;
        RECT 275.235 -98.765 275.565 -98.435 ;
        RECT 275.235 -100.125 275.565 -99.795 ;
        RECT 275.235 -101.485 275.565 -101.155 ;
        RECT 275.235 -102.845 275.565 -102.515 ;
        RECT 275.235 -104.205 275.565 -103.875 ;
        RECT 275.235 -105.565 275.565 -105.235 ;
        RECT 275.235 -106.925 275.565 -106.595 ;
        RECT 275.235 -108.285 275.565 -107.955 ;
        RECT 275.235 -109.645 275.565 -109.315 ;
        RECT 275.235 -111.005 275.565 -110.675 ;
        RECT 275.235 -112.365 275.565 -112.035 ;
        RECT 275.235 -113.725 275.565 -113.395 ;
        RECT 275.235 -115.085 275.565 -114.755 ;
        RECT 275.235 -116.445 275.565 -116.115 ;
        RECT 275.235 -117.805 275.565 -117.475 ;
        RECT 275.235 -119.165 275.565 -118.835 ;
        RECT 275.235 -120.525 275.565 -120.195 ;
        RECT 275.235 -121.885 275.565 -121.555 ;
        RECT 275.235 -123.245 275.565 -122.915 ;
        RECT 275.235 -124.605 275.565 -124.275 ;
        RECT 275.235 -125.965 275.565 -125.635 ;
        RECT 275.235 -127.325 275.565 -126.995 ;
        RECT 275.235 -128.685 275.565 -128.355 ;
        RECT 275.235 -130.045 275.565 -129.715 ;
        RECT 275.235 -131.405 275.565 -131.075 ;
        RECT 275.235 -132.765 275.565 -132.435 ;
        RECT 275.235 -134.125 275.565 -133.795 ;
        RECT 275.235 -135.485 275.565 -135.155 ;
        RECT 275.235 -136.845 275.565 -136.515 ;
        RECT 275.235 -138.205 275.565 -137.875 ;
        RECT 275.235 -139.565 275.565 -139.235 ;
        RECT 275.235 -140.925 275.565 -140.595 ;
        RECT 275.235 -142.285 275.565 -141.955 ;
        RECT 275.235 -143.645 275.565 -143.315 ;
        RECT 275.235 -145.005 275.565 -144.675 ;
        RECT 275.235 -146.365 275.565 -146.035 ;
        RECT 275.235 -147.725 275.565 -147.395 ;
        RECT 275.235 -149.085 275.565 -148.755 ;
        RECT 275.235 -150.445 275.565 -150.115 ;
        RECT 275.235 -151.805 275.565 -151.475 ;
        RECT 275.235 -153.165 275.565 -152.835 ;
        RECT 275.235 -154.525 275.565 -154.195 ;
        RECT 275.235 -155.885 275.565 -155.555 ;
        RECT 275.235 -157.245 275.565 -156.915 ;
        RECT 275.235 -158.605 275.565 -158.275 ;
        RECT 275.235 -159.965 275.565 -159.635 ;
        RECT 275.235 -161.325 275.565 -160.995 ;
        RECT 275.235 -162.685 275.565 -162.355 ;
        RECT 275.235 -164.045 275.565 -163.715 ;
        RECT 275.235 -165.405 275.565 -165.075 ;
        RECT 275.235 -166.765 275.565 -166.435 ;
        RECT 275.235 -168.125 275.565 -167.795 ;
        RECT 275.235 -169.485 275.565 -169.155 ;
        RECT 275.235 -170.845 275.565 -170.515 ;
        RECT 275.235 -172.205 275.565 -171.875 ;
        RECT 275.235 -173.565 275.565 -173.235 ;
        RECT 275.235 -174.925 275.565 -174.595 ;
        RECT 275.235 -176.285 275.565 -175.955 ;
        RECT 275.235 -177.645 275.565 -177.315 ;
        RECT 275.235 -183.29 275.565 -182.16 ;
        RECT 275.24 -183.405 275.56 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 276.595 244.04 276.925 245.17 ;
        RECT 276.595 239.875 276.925 240.205 ;
        RECT 276.595 238.515 276.925 238.845 ;
        RECT 276.595 237.155 276.925 237.485 ;
        RECT 276.6 237.155 276.92 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 276.595 -96.045 276.925 -95.715 ;
        RECT 276.595 -97.405 276.925 -97.075 ;
        RECT 276.595 -98.765 276.925 -98.435 ;
        RECT 276.595 -100.125 276.925 -99.795 ;
        RECT 276.595 -101.485 276.925 -101.155 ;
        RECT 276.595 -102.845 276.925 -102.515 ;
        RECT 276.595 -104.205 276.925 -103.875 ;
        RECT 276.595 -105.565 276.925 -105.235 ;
        RECT 276.595 -106.925 276.925 -106.595 ;
        RECT 276.595 -108.285 276.925 -107.955 ;
        RECT 276.595 -109.645 276.925 -109.315 ;
        RECT 276.595 -111.005 276.925 -110.675 ;
        RECT 276.595 -112.365 276.925 -112.035 ;
        RECT 276.595 -113.725 276.925 -113.395 ;
        RECT 276.595 -115.085 276.925 -114.755 ;
        RECT 276.595 -116.445 276.925 -116.115 ;
        RECT 276.595 -117.805 276.925 -117.475 ;
        RECT 276.595 -119.165 276.925 -118.835 ;
        RECT 276.595 -120.525 276.925 -120.195 ;
        RECT 276.595 -121.885 276.925 -121.555 ;
        RECT 276.595 -123.245 276.925 -122.915 ;
        RECT 276.595 -124.605 276.925 -124.275 ;
        RECT 276.595 -125.965 276.925 -125.635 ;
        RECT 276.595 -127.325 276.925 -126.995 ;
        RECT 276.595 -128.685 276.925 -128.355 ;
        RECT 276.595 -130.045 276.925 -129.715 ;
        RECT 276.595 -131.405 276.925 -131.075 ;
        RECT 276.595 -132.765 276.925 -132.435 ;
        RECT 276.595 -134.125 276.925 -133.795 ;
        RECT 276.595 -135.485 276.925 -135.155 ;
        RECT 276.595 -136.845 276.925 -136.515 ;
        RECT 276.595 -138.205 276.925 -137.875 ;
        RECT 276.595 -139.565 276.925 -139.235 ;
        RECT 276.595 -140.925 276.925 -140.595 ;
        RECT 276.595 -142.285 276.925 -141.955 ;
        RECT 276.595 -143.645 276.925 -143.315 ;
        RECT 276.595 -145.005 276.925 -144.675 ;
        RECT 276.595 -146.365 276.925 -146.035 ;
        RECT 276.595 -147.725 276.925 -147.395 ;
        RECT 276.595 -149.085 276.925 -148.755 ;
        RECT 276.595 -150.445 276.925 -150.115 ;
        RECT 276.595 -151.805 276.925 -151.475 ;
        RECT 276.595 -153.165 276.925 -152.835 ;
        RECT 276.595 -154.525 276.925 -154.195 ;
        RECT 276.595 -155.885 276.925 -155.555 ;
        RECT 276.595 -157.245 276.925 -156.915 ;
        RECT 276.595 -158.605 276.925 -158.275 ;
        RECT 276.595 -159.965 276.925 -159.635 ;
        RECT 276.595 -161.325 276.925 -160.995 ;
        RECT 276.595 -162.685 276.925 -162.355 ;
        RECT 276.595 -164.045 276.925 -163.715 ;
        RECT 276.595 -165.405 276.925 -165.075 ;
        RECT 276.595 -166.765 276.925 -166.435 ;
        RECT 276.595 -168.125 276.925 -167.795 ;
        RECT 276.595 -169.485 276.925 -169.155 ;
        RECT 276.595 -170.845 276.925 -170.515 ;
        RECT 276.595 -172.205 276.925 -171.875 ;
        RECT 276.595 -173.565 276.925 -173.235 ;
        RECT 276.595 -174.925 276.925 -174.595 ;
        RECT 276.595 -176.285 276.925 -175.955 ;
        RECT 276.595 -177.645 276.925 -177.315 ;
        RECT 276.595 -183.29 276.925 -182.16 ;
        RECT 276.6 -183.405 276.92 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 277.16 -94.075 277.49 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 277.955 244.04 278.285 245.17 ;
        RECT 277.955 239.875 278.285 240.205 ;
        RECT 277.955 238.515 278.285 238.845 ;
        RECT 277.955 237.155 278.285 237.485 ;
        RECT 277.96 237.155 278.28 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 279.315 244.04 279.645 245.17 ;
        RECT 279.315 239.875 279.645 240.205 ;
        RECT 279.315 238.515 279.645 238.845 ;
        RECT 279.315 237.155 279.645 237.485 ;
        RECT 279.32 237.155 279.64 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 279.315 -0.845 279.645 -0.515 ;
        RECT 279.315 -2.205 279.645 -1.875 ;
        RECT 279.315 -3.565 279.645 -3.235 ;
        RECT 279.32 -3.565 279.64 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 279.315 -91.965 279.645 -91.635 ;
        RECT 279.315 -93.325 279.645 -92.995 ;
        RECT 279.315 -94.685 279.645 -94.355 ;
        RECT 279.315 -96.045 279.645 -95.715 ;
        RECT 279.315 -97.405 279.645 -97.075 ;
        RECT 279.315 -98.765 279.645 -98.435 ;
        RECT 279.315 -100.125 279.645 -99.795 ;
        RECT 279.315 -101.485 279.645 -101.155 ;
        RECT 279.315 -102.845 279.645 -102.515 ;
        RECT 279.315 -104.205 279.645 -103.875 ;
        RECT 279.315 -105.565 279.645 -105.235 ;
        RECT 279.315 -106.925 279.645 -106.595 ;
        RECT 279.315 -108.285 279.645 -107.955 ;
        RECT 279.315 -109.645 279.645 -109.315 ;
        RECT 279.315 -111.005 279.645 -110.675 ;
        RECT 279.315 -112.365 279.645 -112.035 ;
        RECT 279.315 -113.725 279.645 -113.395 ;
        RECT 279.315 -115.085 279.645 -114.755 ;
        RECT 279.315 -116.445 279.645 -116.115 ;
        RECT 279.315 -117.805 279.645 -117.475 ;
        RECT 279.315 -119.165 279.645 -118.835 ;
        RECT 279.315 -120.525 279.645 -120.195 ;
        RECT 279.315 -121.885 279.645 -121.555 ;
        RECT 279.315 -123.245 279.645 -122.915 ;
        RECT 279.315 -124.605 279.645 -124.275 ;
        RECT 279.315 -125.965 279.645 -125.635 ;
        RECT 279.315 -127.325 279.645 -126.995 ;
        RECT 279.315 -128.685 279.645 -128.355 ;
        RECT 279.315 -130.045 279.645 -129.715 ;
        RECT 279.315 -131.405 279.645 -131.075 ;
        RECT 279.315 -132.765 279.645 -132.435 ;
        RECT 279.315 -134.125 279.645 -133.795 ;
        RECT 279.315 -135.485 279.645 -135.155 ;
        RECT 279.315 -136.845 279.645 -136.515 ;
        RECT 279.315 -138.205 279.645 -137.875 ;
        RECT 279.315 -139.565 279.645 -139.235 ;
        RECT 279.315 -140.925 279.645 -140.595 ;
        RECT 279.315 -142.285 279.645 -141.955 ;
        RECT 279.315 -143.645 279.645 -143.315 ;
        RECT 279.315 -145.005 279.645 -144.675 ;
        RECT 279.315 -146.365 279.645 -146.035 ;
        RECT 279.315 -147.725 279.645 -147.395 ;
        RECT 279.315 -149.085 279.645 -148.755 ;
        RECT 279.315 -150.445 279.645 -150.115 ;
        RECT 279.315 -151.805 279.645 -151.475 ;
        RECT 279.315 -153.165 279.645 -152.835 ;
        RECT 279.315 -154.525 279.645 -154.195 ;
        RECT 279.315 -155.885 279.645 -155.555 ;
        RECT 279.315 -157.245 279.645 -156.915 ;
        RECT 279.315 -158.605 279.645 -158.275 ;
        RECT 279.315 -159.965 279.645 -159.635 ;
        RECT 279.315 -161.325 279.645 -160.995 ;
        RECT 279.315 -162.685 279.645 -162.355 ;
        RECT 279.315 -164.045 279.645 -163.715 ;
        RECT 279.315 -165.405 279.645 -165.075 ;
        RECT 279.315 -166.765 279.645 -166.435 ;
        RECT 279.315 -168.125 279.645 -167.795 ;
        RECT 279.315 -169.485 279.645 -169.155 ;
        RECT 279.315 -170.845 279.645 -170.515 ;
        RECT 279.315 -172.205 279.645 -171.875 ;
        RECT 279.315 -173.565 279.645 -173.235 ;
        RECT 279.315 -174.925 279.645 -174.595 ;
        RECT 279.315 -176.285 279.645 -175.955 ;
        RECT 279.315 -177.645 279.645 -177.315 ;
        RECT 279.315 -183.29 279.645 -182.16 ;
        RECT 279.32 -183.405 279.64 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 280.675 244.04 281.005 245.17 ;
        RECT 280.675 239.875 281.005 240.205 ;
        RECT 280.675 238.515 281.005 238.845 ;
        RECT 280.675 237.155 281.005 237.485 ;
        RECT 280.68 237.155 281 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 280.675 -0.845 281.005 -0.515 ;
        RECT 280.675 -2.205 281.005 -1.875 ;
        RECT 280.675 -3.565 281.005 -3.235 ;
        RECT 280.68 -3.565 281 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 282.035 244.04 282.365 245.17 ;
        RECT 282.035 239.875 282.365 240.205 ;
        RECT 282.035 238.515 282.365 238.845 ;
        RECT 282.035 237.155 282.365 237.485 ;
        RECT 282.04 237.155 282.36 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 282.035 -0.845 282.365 -0.515 ;
        RECT 282.035 -2.205 282.365 -1.875 ;
        RECT 282.035 -3.565 282.365 -3.235 ;
        RECT 282.04 -3.565 282.36 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 282.035 -91.965 282.365 -91.635 ;
        RECT 282.035 -93.325 282.365 -92.995 ;
        RECT 282.035 -94.685 282.365 -94.355 ;
        RECT 282.035 -96.045 282.365 -95.715 ;
        RECT 282.035 -97.405 282.365 -97.075 ;
        RECT 282.035 -98.765 282.365 -98.435 ;
        RECT 282.035 -100.125 282.365 -99.795 ;
        RECT 282.035 -101.485 282.365 -101.155 ;
        RECT 282.035 -102.845 282.365 -102.515 ;
        RECT 282.035 -104.205 282.365 -103.875 ;
        RECT 282.035 -105.565 282.365 -105.235 ;
        RECT 282.035 -106.925 282.365 -106.595 ;
        RECT 282.035 -108.285 282.365 -107.955 ;
        RECT 282.035 -109.645 282.365 -109.315 ;
        RECT 282.035 -111.005 282.365 -110.675 ;
        RECT 282.035 -112.365 282.365 -112.035 ;
        RECT 282.035 -113.725 282.365 -113.395 ;
        RECT 282.035 -115.085 282.365 -114.755 ;
        RECT 282.035 -116.445 282.365 -116.115 ;
        RECT 282.035 -117.805 282.365 -117.475 ;
        RECT 282.035 -119.165 282.365 -118.835 ;
        RECT 282.035 -120.525 282.365 -120.195 ;
        RECT 282.035 -121.885 282.365 -121.555 ;
        RECT 282.035 -123.245 282.365 -122.915 ;
        RECT 282.035 -124.605 282.365 -124.275 ;
        RECT 282.035 -125.965 282.365 -125.635 ;
        RECT 282.035 -127.325 282.365 -126.995 ;
        RECT 282.035 -128.685 282.365 -128.355 ;
        RECT 282.035 -130.045 282.365 -129.715 ;
        RECT 282.035 -131.405 282.365 -131.075 ;
        RECT 282.035 -132.765 282.365 -132.435 ;
        RECT 282.035 -134.125 282.365 -133.795 ;
        RECT 282.035 -135.485 282.365 -135.155 ;
        RECT 282.035 -136.845 282.365 -136.515 ;
        RECT 282.035 -138.205 282.365 -137.875 ;
        RECT 282.035 -139.565 282.365 -139.235 ;
        RECT 282.035 -140.925 282.365 -140.595 ;
        RECT 282.035 -142.285 282.365 -141.955 ;
        RECT 282.035 -143.645 282.365 -143.315 ;
        RECT 282.035 -145.005 282.365 -144.675 ;
        RECT 282.035 -146.365 282.365 -146.035 ;
        RECT 282.035 -147.725 282.365 -147.395 ;
        RECT 282.035 -149.085 282.365 -148.755 ;
        RECT 282.035 -150.445 282.365 -150.115 ;
        RECT 282.035 -151.805 282.365 -151.475 ;
        RECT 282.035 -153.165 282.365 -152.835 ;
        RECT 282.035 -154.525 282.365 -154.195 ;
        RECT 282.035 -155.885 282.365 -155.555 ;
        RECT 282.035 -157.245 282.365 -156.915 ;
        RECT 282.035 -158.605 282.365 -158.275 ;
        RECT 282.035 -159.965 282.365 -159.635 ;
        RECT 282.035 -161.325 282.365 -160.995 ;
        RECT 282.035 -162.685 282.365 -162.355 ;
        RECT 282.035 -164.045 282.365 -163.715 ;
        RECT 282.035 -165.405 282.365 -165.075 ;
        RECT 282.035 -166.765 282.365 -166.435 ;
        RECT 282.035 -168.125 282.365 -167.795 ;
        RECT 282.035 -169.485 282.365 -169.155 ;
        RECT 282.035 -170.845 282.365 -170.515 ;
        RECT 282.035 -172.205 282.365 -171.875 ;
        RECT 282.035 -173.565 282.365 -173.235 ;
        RECT 282.035 -174.925 282.365 -174.595 ;
        RECT 282.035 -176.285 282.365 -175.955 ;
        RECT 282.035 -177.645 282.365 -177.315 ;
        RECT 282.035 -183.29 282.365 -182.16 ;
        RECT 282.04 -183.405 282.36 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 283.26 -94.075 283.59 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 283.395 244.04 283.725 245.17 ;
        RECT 283.395 239.875 283.725 240.205 ;
        RECT 283.395 238.515 283.725 238.845 ;
        RECT 283.395 237.155 283.725 237.485 ;
        RECT 283.4 237.155 283.72 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 283.395 -96.045 283.725 -95.715 ;
        RECT 283.395 -97.405 283.725 -97.075 ;
        RECT 283.395 -98.765 283.725 -98.435 ;
        RECT 283.395 -100.125 283.725 -99.795 ;
        RECT 283.395 -101.485 283.725 -101.155 ;
        RECT 283.395 -102.845 283.725 -102.515 ;
        RECT 283.395 -104.205 283.725 -103.875 ;
        RECT 283.395 -105.565 283.725 -105.235 ;
        RECT 283.395 -106.925 283.725 -106.595 ;
        RECT 283.395 -108.285 283.725 -107.955 ;
        RECT 283.395 -109.645 283.725 -109.315 ;
        RECT 283.395 -111.005 283.725 -110.675 ;
        RECT 283.395 -112.365 283.725 -112.035 ;
        RECT 283.395 -113.725 283.725 -113.395 ;
        RECT 283.395 -115.085 283.725 -114.755 ;
        RECT 283.395 -116.445 283.725 -116.115 ;
        RECT 283.395 -117.805 283.725 -117.475 ;
        RECT 283.395 -119.165 283.725 -118.835 ;
        RECT 283.395 -120.525 283.725 -120.195 ;
        RECT 283.395 -121.885 283.725 -121.555 ;
        RECT 283.395 -123.245 283.725 -122.915 ;
        RECT 283.395 -124.605 283.725 -124.275 ;
        RECT 283.395 -125.965 283.725 -125.635 ;
        RECT 283.395 -127.325 283.725 -126.995 ;
        RECT 283.395 -128.685 283.725 -128.355 ;
        RECT 283.395 -130.045 283.725 -129.715 ;
        RECT 283.395 -131.405 283.725 -131.075 ;
        RECT 283.395 -132.765 283.725 -132.435 ;
        RECT 283.395 -134.125 283.725 -133.795 ;
        RECT 283.395 -135.485 283.725 -135.155 ;
        RECT 283.395 -136.845 283.725 -136.515 ;
        RECT 283.395 -138.205 283.725 -137.875 ;
        RECT 283.395 -139.565 283.725 -139.235 ;
        RECT 283.395 -140.925 283.725 -140.595 ;
        RECT 283.395 -142.285 283.725 -141.955 ;
        RECT 283.395 -143.645 283.725 -143.315 ;
        RECT 283.395 -145.005 283.725 -144.675 ;
        RECT 283.395 -146.365 283.725 -146.035 ;
        RECT 283.395 -147.725 283.725 -147.395 ;
        RECT 283.395 -149.085 283.725 -148.755 ;
        RECT 283.395 -150.445 283.725 -150.115 ;
        RECT 283.395 -151.805 283.725 -151.475 ;
        RECT 283.395 -153.165 283.725 -152.835 ;
        RECT 283.395 -154.525 283.725 -154.195 ;
        RECT 283.395 -155.885 283.725 -155.555 ;
        RECT 283.395 -157.245 283.725 -156.915 ;
        RECT 283.395 -158.605 283.725 -158.275 ;
        RECT 283.395 -159.965 283.725 -159.635 ;
        RECT 283.395 -161.325 283.725 -160.995 ;
        RECT 283.395 -162.685 283.725 -162.355 ;
        RECT 283.395 -164.045 283.725 -163.715 ;
        RECT 283.395 -165.405 283.725 -165.075 ;
        RECT 283.395 -166.765 283.725 -166.435 ;
        RECT 283.395 -168.125 283.725 -167.795 ;
        RECT 283.395 -169.485 283.725 -169.155 ;
        RECT 283.395 -170.845 283.725 -170.515 ;
        RECT 283.395 -172.205 283.725 -171.875 ;
        RECT 283.395 -173.565 283.725 -173.235 ;
        RECT 283.395 -174.925 283.725 -174.595 ;
        RECT 283.395 -176.285 283.725 -175.955 ;
        RECT 283.395 -177.645 283.725 -177.315 ;
        RECT 283.395 -183.29 283.725 -182.16 ;
        RECT 283.4 -183.405 283.72 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 284.755 244.04 285.085 245.17 ;
        RECT 284.755 239.875 285.085 240.205 ;
        RECT 284.755 238.515 285.085 238.845 ;
        RECT 284.755 237.155 285.085 237.485 ;
        RECT 284.76 237.155 285.08 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 284.755 -0.845 285.085 -0.515 ;
        RECT 284.755 -2.205 285.085 -1.875 ;
        RECT 284.755 -3.565 285.085 -3.235 ;
        RECT 284.76 -3.565 285.08 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 286.115 244.04 286.445 245.17 ;
        RECT 286.115 239.875 286.445 240.205 ;
        RECT 286.115 238.515 286.445 238.845 ;
        RECT 286.115 237.155 286.445 237.485 ;
        RECT 286.12 237.155 286.44 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 286.115 -0.845 286.445 -0.515 ;
        RECT 286.115 -2.205 286.445 -1.875 ;
        RECT 286.115 -3.565 286.445 -3.235 ;
        RECT 286.12 -3.565 286.44 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 287.475 244.04 287.805 245.17 ;
        RECT 287.475 239.875 287.805 240.205 ;
        RECT 287.475 238.515 287.805 238.845 ;
        RECT 287.475 237.155 287.805 237.485 ;
        RECT 287.48 237.155 287.8 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 287.475 -0.845 287.805 -0.515 ;
        RECT 287.475 -2.205 287.805 -1.875 ;
        RECT 287.475 -3.565 287.805 -3.235 ;
        RECT 287.48 -3.565 287.8 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 287.475 -91.965 287.805 -91.635 ;
        RECT 287.475 -93.325 287.805 -92.995 ;
        RECT 287.475 -94.685 287.805 -94.355 ;
        RECT 287.475 -96.045 287.805 -95.715 ;
        RECT 287.475 -97.405 287.805 -97.075 ;
        RECT 287.475 -98.765 287.805 -98.435 ;
        RECT 287.475 -100.125 287.805 -99.795 ;
        RECT 287.475 -101.485 287.805 -101.155 ;
        RECT 287.475 -102.845 287.805 -102.515 ;
        RECT 287.475 -104.205 287.805 -103.875 ;
        RECT 287.475 -105.565 287.805 -105.235 ;
        RECT 287.475 -106.925 287.805 -106.595 ;
        RECT 287.475 -108.285 287.805 -107.955 ;
        RECT 287.475 -109.645 287.805 -109.315 ;
        RECT 287.475 -111.005 287.805 -110.675 ;
        RECT 287.475 -112.365 287.805 -112.035 ;
        RECT 287.475 -113.725 287.805 -113.395 ;
        RECT 287.475 -115.085 287.805 -114.755 ;
        RECT 287.475 -116.445 287.805 -116.115 ;
        RECT 287.475 -117.805 287.805 -117.475 ;
        RECT 287.475 -119.165 287.805 -118.835 ;
        RECT 287.475 -120.525 287.805 -120.195 ;
        RECT 287.475 -121.885 287.805 -121.555 ;
        RECT 287.475 -123.245 287.805 -122.915 ;
        RECT 287.475 -124.605 287.805 -124.275 ;
        RECT 287.475 -125.965 287.805 -125.635 ;
        RECT 287.475 -127.325 287.805 -126.995 ;
        RECT 287.475 -128.685 287.805 -128.355 ;
        RECT 287.475 -130.045 287.805 -129.715 ;
        RECT 287.475 -131.405 287.805 -131.075 ;
        RECT 287.475 -132.765 287.805 -132.435 ;
        RECT 287.475 -134.125 287.805 -133.795 ;
        RECT 287.475 -135.485 287.805 -135.155 ;
        RECT 287.475 -136.845 287.805 -136.515 ;
        RECT 287.475 -138.205 287.805 -137.875 ;
        RECT 287.475 -139.565 287.805 -139.235 ;
        RECT 287.475 -140.925 287.805 -140.595 ;
        RECT 287.475 -142.285 287.805 -141.955 ;
        RECT 287.475 -143.645 287.805 -143.315 ;
        RECT 287.475 -145.005 287.805 -144.675 ;
        RECT 287.475 -146.365 287.805 -146.035 ;
        RECT 287.475 -147.725 287.805 -147.395 ;
        RECT 287.475 -149.085 287.805 -148.755 ;
        RECT 287.475 -150.445 287.805 -150.115 ;
        RECT 287.475 -151.805 287.805 -151.475 ;
        RECT 287.475 -153.165 287.805 -152.835 ;
        RECT 287.475 -154.525 287.805 -154.195 ;
        RECT 287.475 -155.885 287.805 -155.555 ;
        RECT 287.475 -157.245 287.805 -156.915 ;
        RECT 287.475 -158.605 287.805 -158.275 ;
        RECT 287.475 -159.965 287.805 -159.635 ;
        RECT 287.475 -161.325 287.805 -160.995 ;
        RECT 287.475 -162.685 287.805 -162.355 ;
        RECT 287.475 -164.045 287.805 -163.715 ;
        RECT 287.475 -165.405 287.805 -165.075 ;
        RECT 287.475 -166.765 287.805 -166.435 ;
        RECT 287.475 -168.125 287.805 -167.795 ;
        RECT 287.475 -169.485 287.805 -169.155 ;
        RECT 287.475 -170.845 287.805 -170.515 ;
        RECT 287.475 -172.205 287.805 -171.875 ;
        RECT 287.475 -173.565 287.805 -173.235 ;
        RECT 287.475 -174.925 287.805 -174.595 ;
        RECT 287.475 -176.285 287.805 -175.955 ;
        RECT 287.475 -177.645 287.805 -177.315 ;
        RECT 287.475 -183.29 287.805 -182.16 ;
        RECT 287.48 -183.405 287.8 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 288.835 244.04 289.165 245.17 ;
        RECT 288.835 239.875 289.165 240.205 ;
        RECT 288.835 238.515 289.165 238.845 ;
        RECT 288.835 237.155 289.165 237.485 ;
        RECT 288.84 237.155 289.16 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 288.835 -96.045 289.165 -95.715 ;
        RECT 288.835 -97.405 289.165 -97.075 ;
        RECT 288.835 -98.765 289.165 -98.435 ;
        RECT 288.835 -100.125 289.165 -99.795 ;
        RECT 288.835 -101.485 289.165 -101.155 ;
        RECT 288.835 -102.845 289.165 -102.515 ;
        RECT 288.835 -104.205 289.165 -103.875 ;
        RECT 288.835 -105.565 289.165 -105.235 ;
        RECT 288.835 -106.925 289.165 -106.595 ;
        RECT 288.835 -108.285 289.165 -107.955 ;
        RECT 288.835 -109.645 289.165 -109.315 ;
        RECT 288.835 -111.005 289.165 -110.675 ;
        RECT 288.835 -112.365 289.165 -112.035 ;
        RECT 288.835 -113.725 289.165 -113.395 ;
        RECT 288.835 -115.085 289.165 -114.755 ;
        RECT 288.835 -116.445 289.165 -116.115 ;
        RECT 288.835 -117.805 289.165 -117.475 ;
        RECT 288.835 -119.165 289.165 -118.835 ;
        RECT 288.835 -120.525 289.165 -120.195 ;
        RECT 288.835 -121.885 289.165 -121.555 ;
        RECT 288.835 -123.245 289.165 -122.915 ;
        RECT 288.835 -124.605 289.165 -124.275 ;
        RECT 288.835 -125.965 289.165 -125.635 ;
        RECT 288.835 -127.325 289.165 -126.995 ;
        RECT 288.835 -128.685 289.165 -128.355 ;
        RECT 288.835 -130.045 289.165 -129.715 ;
        RECT 288.835 -131.405 289.165 -131.075 ;
        RECT 288.835 -132.765 289.165 -132.435 ;
        RECT 288.835 -134.125 289.165 -133.795 ;
        RECT 288.835 -135.485 289.165 -135.155 ;
        RECT 288.835 -136.845 289.165 -136.515 ;
        RECT 288.835 -138.205 289.165 -137.875 ;
        RECT 288.835 -139.565 289.165 -139.235 ;
        RECT 288.835 -140.925 289.165 -140.595 ;
        RECT 288.835 -142.285 289.165 -141.955 ;
        RECT 288.835 -143.645 289.165 -143.315 ;
        RECT 288.835 -145.005 289.165 -144.675 ;
        RECT 288.835 -146.365 289.165 -146.035 ;
        RECT 288.835 -147.725 289.165 -147.395 ;
        RECT 288.835 -149.085 289.165 -148.755 ;
        RECT 288.835 -150.445 289.165 -150.115 ;
        RECT 288.835 -151.805 289.165 -151.475 ;
        RECT 288.835 -153.165 289.165 -152.835 ;
        RECT 288.835 -154.525 289.165 -154.195 ;
        RECT 288.835 -155.885 289.165 -155.555 ;
        RECT 288.835 -157.245 289.165 -156.915 ;
        RECT 288.835 -158.605 289.165 -158.275 ;
        RECT 288.835 -159.965 289.165 -159.635 ;
        RECT 288.835 -161.325 289.165 -160.995 ;
        RECT 288.835 -162.685 289.165 -162.355 ;
        RECT 288.835 -164.045 289.165 -163.715 ;
        RECT 288.835 -165.405 289.165 -165.075 ;
        RECT 288.835 -166.765 289.165 -166.435 ;
        RECT 288.835 -168.125 289.165 -167.795 ;
        RECT 288.835 -169.485 289.165 -169.155 ;
        RECT 288.835 -170.845 289.165 -170.515 ;
        RECT 288.835 -172.205 289.165 -171.875 ;
        RECT 288.835 -173.565 289.165 -173.235 ;
        RECT 288.835 -174.925 289.165 -174.595 ;
        RECT 288.835 -176.285 289.165 -175.955 ;
        RECT 288.835 -177.645 289.165 -177.315 ;
        RECT 288.835 -183.29 289.165 -182.16 ;
        RECT 288.84 -183.405 289.16 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 289.36 -94.075 289.69 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 290.195 244.04 290.525 245.17 ;
        RECT 290.195 239.875 290.525 240.205 ;
        RECT 290.195 238.515 290.525 238.845 ;
        RECT 290.195 237.155 290.525 237.485 ;
        RECT 290.2 237.155 290.52 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 291.555 244.04 291.885 245.17 ;
        RECT 291.555 239.875 291.885 240.205 ;
        RECT 291.555 238.515 291.885 238.845 ;
        RECT 291.555 237.155 291.885 237.485 ;
        RECT 291.56 237.155 291.88 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 291.555 -0.845 291.885 -0.515 ;
        RECT 291.555 -2.205 291.885 -1.875 ;
        RECT 291.555 -3.565 291.885 -3.235 ;
        RECT 291.56 -3.565 291.88 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 291.555 -91.965 291.885 -91.635 ;
        RECT 291.555 -93.325 291.885 -92.995 ;
        RECT 291.555 -94.685 291.885 -94.355 ;
        RECT 291.555 -96.045 291.885 -95.715 ;
        RECT 291.555 -97.405 291.885 -97.075 ;
        RECT 291.555 -98.765 291.885 -98.435 ;
        RECT 291.555 -100.125 291.885 -99.795 ;
        RECT 291.555 -101.485 291.885 -101.155 ;
        RECT 291.555 -102.845 291.885 -102.515 ;
        RECT 291.555 -104.205 291.885 -103.875 ;
        RECT 291.555 -105.565 291.885 -105.235 ;
        RECT 291.555 -106.925 291.885 -106.595 ;
        RECT 291.555 -108.285 291.885 -107.955 ;
        RECT 291.555 -109.645 291.885 -109.315 ;
        RECT 291.555 -111.005 291.885 -110.675 ;
        RECT 291.555 -112.365 291.885 -112.035 ;
        RECT 291.555 -113.725 291.885 -113.395 ;
        RECT 291.555 -115.085 291.885 -114.755 ;
        RECT 291.555 -116.445 291.885 -116.115 ;
        RECT 291.555 -117.805 291.885 -117.475 ;
        RECT 291.555 -119.165 291.885 -118.835 ;
        RECT 291.555 -120.525 291.885 -120.195 ;
        RECT 291.555 -121.885 291.885 -121.555 ;
        RECT 291.555 -123.245 291.885 -122.915 ;
        RECT 291.555 -124.605 291.885 -124.275 ;
        RECT 291.555 -125.965 291.885 -125.635 ;
        RECT 291.555 -127.325 291.885 -126.995 ;
        RECT 291.555 -128.685 291.885 -128.355 ;
        RECT 291.555 -130.045 291.885 -129.715 ;
        RECT 291.555 -131.405 291.885 -131.075 ;
        RECT 291.555 -132.765 291.885 -132.435 ;
        RECT 291.555 -134.125 291.885 -133.795 ;
        RECT 291.555 -135.485 291.885 -135.155 ;
        RECT 291.555 -136.845 291.885 -136.515 ;
        RECT 291.555 -138.205 291.885 -137.875 ;
        RECT 291.555 -139.565 291.885 -139.235 ;
        RECT 291.555 -140.925 291.885 -140.595 ;
        RECT 291.555 -142.285 291.885 -141.955 ;
        RECT 291.555 -143.645 291.885 -143.315 ;
        RECT 291.555 -145.005 291.885 -144.675 ;
        RECT 291.555 -146.365 291.885 -146.035 ;
        RECT 291.555 -147.725 291.885 -147.395 ;
        RECT 291.555 -149.085 291.885 -148.755 ;
        RECT 291.555 -150.445 291.885 -150.115 ;
        RECT 291.555 -151.805 291.885 -151.475 ;
        RECT 291.555 -153.165 291.885 -152.835 ;
        RECT 291.555 -154.525 291.885 -154.195 ;
        RECT 291.555 -155.885 291.885 -155.555 ;
        RECT 291.555 -157.245 291.885 -156.915 ;
        RECT 291.555 -158.605 291.885 -158.275 ;
        RECT 291.555 -159.965 291.885 -159.635 ;
        RECT 291.555 -161.325 291.885 -160.995 ;
        RECT 291.555 -162.685 291.885 -162.355 ;
        RECT 291.555 -164.045 291.885 -163.715 ;
        RECT 291.555 -165.405 291.885 -165.075 ;
        RECT 291.555 -166.765 291.885 -166.435 ;
        RECT 291.555 -168.125 291.885 -167.795 ;
        RECT 291.555 -169.485 291.885 -169.155 ;
        RECT 291.555 -170.845 291.885 -170.515 ;
        RECT 291.555 -172.205 291.885 -171.875 ;
        RECT 291.555 -173.565 291.885 -173.235 ;
        RECT 291.555 -174.925 291.885 -174.595 ;
        RECT 291.555 -176.285 291.885 -175.955 ;
        RECT 291.555 -177.645 291.885 -177.315 ;
        RECT 291.555 -183.29 291.885 -182.16 ;
        RECT 291.56 -183.405 291.88 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 292.915 244.04 293.245 245.17 ;
        RECT 292.915 239.875 293.245 240.205 ;
        RECT 292.915 238.515 293.245 238.845 ;
        RECT 292.915 237.155 293.245 237.485 ;
        RECT 292.92 237.155 293.24 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 292.915 -0.845 293.245 -0.515 ;
        RECT 292.915 -2.205 293.245 -1.875 ;
        RECT 292.915 -3.565 293.245 -3.235 ;
        RECT 292.92 -3.565 293.24 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 294.275 244.04 294.605 245.17 ;
        RECT 294.275 239.875 294.605 240.205 ;
        RECT 294.275 238.515 294.605 238.845 ;
        RECT 294.275 237.155 294.605 237.485 ;
        RECT 294.28 237.155 294.6 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 294.275 -0.845 294.605 -0.515 ;
        RECT 294.275 -2.205 294.605 -1.875 ;
        RECT 294.275 -3.565 294.605 -3.235 ;
        RECT 294.28 -3.565 294.6 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 294.275 -91.965 294.605 -91.635 ;
        RECT 294.275 -93.325 294.605 -92.995 ;
        RECT 294.275 -94.685 294.605 -94.355 ;
        RECT 294.275 -96.045 294.605 -95.715 ;
        RECT 294.275 -97.405 294.605 -97.075 ;
        RECT 294.275 -98.765 294.605 -98.435 ;
        RECT 294.275 -100.125 294.605 -99.795 ;
        RECT 294.275 -101.485 294.605 -101.155 ;
        RECT 294.275 -102.845 294.605 -102.515 ;
        RECT 294.275 -104.205 294.605 -103.875 ;
        RECT 294.275 -105.565 294.605 -105.235 ;
        RECT 294.275 -106.925 294.605 -106.595 ;
        RECT 294.275 -108.285 294.605 -107.955 ;
        RECT 294.275 -109.645 294.605 -109.315 ;
        RECT 294.275 -111.005 294.605 -110.675 ;
        RECT 294.275 -112.365 294.605 -112.035 ;
        RECT 294.275 -113.725 294.605 -113.395 ;
        RECT 294.275 -115.085 294.605 -114.755 ;
        RECT 294.275 -116.445 294.605 -116.115 ;
        RECT 294.275 -117.805 294.605 -117.475 ;
        RECT 294.275 -119.165 294.605 -118.835 ;
        RECT 294.275 -120.525 294.605 -120.195 ;
        RECT 294.275 -121.885 294.605 -121.555 ;
        RECT 294.275 -123.245 294.605 -122.915 ;
        RECT 294.275 -124.605 294.605 -124.275 ;
        RECT 294.275 -125.965 294.605 -125.635 ;
        RECT 294.275 -127.325 294.605 -126.995 ;
        RECT 294.275 -128.685 294.605 -128.355 ;
        RECT 294.275 -130.045 294.605 -129.715 ;
        RECT 294.275 -131.405 294.605 -131.075 ;
        RECT 294.275 -132.765 294.605 -132.435 ;
        RECT 294.275 -134.125 294.605 -133.795 ;
        RECT 294.275 -135.485 294.605 -135.155 ;
        RECT 294.275 -136.845 294.605 -136.515 ;
        RECT 294.275 -138.205 294.605 -137.875 ;
        RECT 294.275 -139.565 294.605 -139.235 ;
        RECT 294.275 -140.925 294.605 -140.595 ;
        RECT 294.275 -142.285 294.605 -141.955 ;
        RECT 294.275 -143.645 294.605 -143.315 ;
        RECT 294.275 -145.005 294.605 -144.675 ;
        RECT 294.275 -146.365 294.605 -146.035 ;
        RECT 294.275 -147.725 294.605 -147.395 ;
        RECT 294.275 -149.085 294.605 -148.755 ;
        RECT 294.275 -150.445 294.605 -150.115 ;
        RECT 294.275 -151.805 294.605 -151.475 ;
        RECT 294.275 -153.165 294.605 -152.835 ;
        RECT 294.275 -154.525 294.605 -154.195 ;
        RECT 294.275 -155.885 294.605 -155.555 ;
        RECT 294.275 -157.245 294.605 -156.915 ;
        RECT 294.275 -158.605 294.605 -158.275 ;
        RECT 294.275 -159.965 294.605 -159.635 ;
        RECT 294.275 -161.325 294.605 -160.995 ;
        RECT 294.275 -162.685 294.605 -162.355 ;
        RECT 294.275 -164.045 294.605 -163.715 ;
        RECT 294.275 -165.405 294.605 -165.075 ;
        RECT 294.275 -166.765 294.605 -166.435 ;
        RECT 294.275 -168.125 294.605 -167.795 ;
        RECT 294.275 -169.485 294.605 -169.155 ;
        RECT 294.275 -170.845 294.605 -170.515 ;
        RECT 294.275 -172.205 294.605 -171.875 ;
        RECT 294.275 -173.565 294.605 -173.235 ;
        RECT 294.275 -174.925 294.605 -174.595 ;
        RECT 294.275 -176.285 294.605 -175.955 ;
        RECT 294.275 -177.645 294.605 -177.315 ;
        RECT 294.275 -183.29 294.605 -182.16 ;
        RECT 294.28 -183.405 294.6 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 295.46 -94.075 295.79 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 295.635 244.04 295.965 245.17 ;
        RECT 295.635 239.875 295.965 240.205 ;
        RECT 295.635 238.515 295.965 238.845 ;
        RECT 295.635 237.155 295.965 237.485 ;
        RECT 295.64 237.155 295.96 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 295.635 -96.045 295.965 -95.715 ;
        RECT 295.635 -97.405 295.965 -97.075 ;
        RECT 295.635 -98.765 295.965 -98.435 ;
        RECT 295.635 -100.125 295.965 -99.795 ;
        RECT 295.635 -101.485 295.965 -101.155 ;
        RECT 295.635 -102.845 295.965 -102.515 ;
        RECT 295.635 -104.205 295.965 -103.875 ;
        RECT 295.635 -105.565 295.965 -105.235 ;
        RECT 295.635 -106.925 295.965 -106.595 ;
        RECT 295.635 -108.285 295.965 -107.955 ;
        RECT 295.635 -109.645 295.965 -109.315 ;
        RECT 295.635 -111.005 295.965 -110.675 ;
        RECT 295.635 -112.365 295.965 -112.035 ;
        RECT 295.635 -113.725 295.965 -113.395 ;
        RECT 295.635 -115.085 295.965 -114.755 ;
        RECT 295.635 -116.445 295.965 -116.115 ;
        RECT 295.635 -117.805 295.965 -117.475 ;
        RECT 295.635 -119.165 295.965 -118.835 ;
        RECT 295.635 -120.525 295.965 -120.195 ;
        RECT 295.635 -121.885 295.965 -121.555 ;
        RECT 295.635 -123.245 295.965 -122.915 ;
        RECT 295.635 -124.605 295.965 -124.275 ;
        RECT 295.635 -125.965 295.965 -125.635 ;
        RECT 295.635 -127.325 295.965 -126.995 ;
        RECT 295.635 -128.685 295.965 -128.355 ;
        RECT 295.635 -130.045 295.965 -129.715 ;
        RECT 295.635 -131.405 295.965 -131.075 ;
        RECT 295.635 -132.765 295.965 -132.435 ;
        RECT 295.635 -134.125 295.965 -133.795 ;
        RECT 295.635 -135.485 295.965 -135.155 ;
        RECT 295.635 -136.845 295.965 -136.515 ;
        RECT 295.635 -138.205 295.965 -137.875 ;
        RECT 295.635 -139.565 295.965 -139.235 ;
        RECT 295.635 -140.925 295.965 -140.595 ;
        RECT 295.635 -142.285 295.965 -141.955 ;
        RECT 295.635 -143.645 295.965 -143.315 ;
        RECT 295.635 -145.005 295.965 -144.675 ;
        RECT 295.635 -146.365 295.965 -146.035 ;
        RECT 295.635 -147.725 295.965 -147.395 ;
        RECT 295.635 -149.085 295.965 -148.755 ;
        RECT 295.635 -150.445 295.965 -150.115 ;
        RECT 295.635 -151.805 295.965 -151.475 ;
        RECT 295.635 -153.165 295.965 -152.835 ;
        RECT 295.635 -154.525 295.965 -154.195 ;
        RECT 295.635 -155.885 295.965 -155.555 ;
        RECT 295.635 -157.245 295.965 -156.915 ;
        RECT 295.635 -158.605 295.965 -158.275 ;
        RECT 295.635 -159.965 295.965 -159.635 ;
        RECT 295.635 -161.325 295.965 -160.995 ;
        RECT 295.635 -162.685 295.965 -162.355 ;
        RECT 295.635 -164.045 295.965 -163.715 ;
        RECT 295.635 -165.405 295.965 -165.075 ;
        RECT 295.635 -166.765 295.965 -166.435 ;
        RECT 295.635 -168.125 295.965 -167.795 ;
        RECT 295.635 -169.485 295.965 -169.155 ;
        RECT 295.635 -170.845 295.965 -170.515 ;
        RECT 295.635 -172.205 295.965 -171.875 ;
        RECT 295.635 -173.565 295.965 -173.235 ;
        RECT 295.635 -174.925 295.965 -174.595 ;
        RECT 295.635 -176.285 295.965 -175.955 ;
        RECT 295.635 -177.645 295.965 -177.315 ;
        RECT 295.635 -183.29 295.965 -182.16 ;
        RECT 295.64 -183.405 295.96 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 296.995 244.04 297.325 245.17 ;
        RECT 296.995 239.875 297.325 240.205 ;
        RECT 296.995 238.515 297.325 238.845 ;
        RECT 296.995 237.155 297.325 237.485 ;
        RECT 297 237.155 297.32 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 296.995 -0.845 297.325 -0.515 ;
        RECT 296.995 -2.205 297.325 -1.875 ;
        RECT 296.995 -3.565 297.325 -3.235 ;
        RECT 297 -3.565 297.32 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 298.355 244.04 298.685 245.17 ;
        RECT 298.355 239.875 298.685 240.205 ;
        RECT 298.355 238.515 298.685 238.845 ;
        RECT 298.355 237.155 298.685 237.485 ;
        RECT 298.36 237.155 298.68 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 298.355 -0.845 298.685 -0.515 ;
        RECT 298.355 -2.205 298.685 -1.875 ;
        RECT 298.355 -3.565 298.685 -3.235 ;
        RECT 298.36 -3.565 298.68 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 299.715 244.04 300.045 245.17 ;
        RECT 299.715 239.875 300.045 240.205 ;
        RECT 299.715 238.515 300.045 238.845 ;
        RECT 299.715 237.155 300.045 237.485 ;
        RECT 299.72 237.155 300.04 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 299.715 -0.845 300.045 -0.515 ;
        RECT 299.715 -2.205 300.045 -1.875 ;
        RECT 299.715 -3.565 300.045 -3.235 ;
        RECT 299.72 -3.565 300.04 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 301.075 244.04 301.405 245.17 ;
        RECT 301.075 239.875 301.405 240.205 ;
        RECT 301.075 238.515 301.405 238.845 ;
        RECT 301.075 237.155 301.405 237.485 ;
        RECT 301.08 237.155 301.4 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 301.075 -96.045 301.405 -95.715 ;
        RECT 301.075 -97.405 301.405 -97.075 ;
        RECT 301.075 -98.765 301.405 -98.435 ;
        RECT 301.075 -100.125 301.405 -99.795 ;
        RECT 301.075 -101.485 301.405 -101.155 ;
        RECT 301.075 -102.845 301.405 -102.515 ;
        RECT 301.075 -104.205 301.405 -103.875 ;
        RECT 301.075 -105.565 301.405 -105.235 ;
        RECT 301.075 -106.925 301.405 -106.595 ;
        RECT 301.075 -108.285 301.405 -107.955 ;
        RECT 301.075 -109.645 301.405 -109.315 ;
        RECT 301.075 -111.005 301.405 -110.675 ;
        RECT 301.075 -112.365 301.405 -112.035 ;
        RECT 301.075 -113.725 301.405 -113.395 ;
        RECT 301.075 -115.085 301.405 -114.755 ;
        RECT 301.075 -116.445 301.405 -116.115 ;
        RECT 301.075 -117.805 301.405 -117.475 ;
        RECT 301.075 -119.165 301.405 -118.835 ;
        RECT 301.075 -120.525 301.405 -120.195 ;
        RECT 301.075 -121.885 301.405 -121.555 ;
        RECT 301.075 -123.245 301.405 -122.915 ;
        RECT 301.075 -124.605 301.405 -124.275 ;
        RECT 301.075 -125.965 301.405 -125.635 ;
        RECT 301.075 -127.325 301.405 -126.995 ;
        RECT 301.075 -128.685 301.405 -128.355 ;
        RECT 301.075 -130.045 301.405 -129.715 ;
        RECT 301.075 -131.405 301.405 -131.075 ;
        RECT 301.075 -132.765 301.405 -132.435 ;
        RECT 301.075 -134.125 301.405 -133.795 ;
        RECT 301.075 -135.485 301.405 -135.155 ;
        RECT 301.075 -136.845 301.405 -136.515 ;
        RECT 301.075 -138.205 301.405 -137.875 ;
        RECT 301.075 -139.565 301.405 -139.235 ;
        RECT 301.075 -140.925 301.405 -140.595 ;
        RECT 301.075 -142.285 301.405 -141.955 ;
        RECT 301.075 -143.645 301.405 -143.315 ;
        RECT 301.075 -145.005 301.405 -144.675 ;
        RECT 301.075 -146.365 301.405 -146.035 ;
        RECT 301.075 -147.725 301.405 -147.395 ;
        RECT 301.075 -149.085 301.405 -148.755 ;
        RECT 301.075 -150.445 301.405 -150.115 ;
        RECT 301.075 -151.805 301.405 -151.475 ;
        RECT 301.075 -153.165 301.405 -152.835 ;
        RECT 301.075 -154.525 301.405 -154.195 ;
        RECT 301.075 -155.885 301.405 -155.555 ;
        RECT 301.075 -157.245 301.405 -156.915 ;
        RECT 301.075 -158.605 301.405 -158.275 ;
        RECT 301.075 -159.965 301.405 -159.635 ;
        RECT 301.075 -161.325 301.405 -160.995 ;
        RECT 301.075 -162.685 301.405 -162.355 ;
        RECT 301.075 -164.045 301.405 -163.715 ;
        RECT 301.075 -165.405 301.405 -165.075 ;
        RECT 301.075 -166.765 301.405 -166.435 ;
        RECT 301.075 -168.125 301.405 -167.795 ;
        RECT 301.075 -169.485 301.405 -169.155 ;
        RECT 301.075 -170.845 301.405 -170.515 ;
        RECT 301.075 -172.205 301.405 -171.875 ;
        RECT 301.075 -173.565 301.405 -173.235 ;
        RECT 301.075 -174.925 301.405 -174.595 ;
        RECT 301.075 -176.285 301.405 -175.955 ;
        RECT 301.075 -177.645 301.405 -177.315 ;
        RECT 301.075 -183.29 301.405 -182.16 ;
        RECT 301.08 -183.405 301.4 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 301.56 -94.075 301.89 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 302.435 244.04 302.765 245.17 ;
        RECT 302.435 239.875 302.765 240.205 ;
        RECT 302.435 238.515 302.765 238.845 ;
        RECT 302.435 237.155 302.765 237.485 ;
        RECT 302.44 237.155 302.76 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 303.795 244.04 304.125 245.17 ;
        RECT 303.795 239.875 304.125 240.205 ;
        RECT 303.795 238.515 304.125 238.845 ;
        RECT 303.795 237.155 304.125 237.485 ;
        RECT 303.8 237.155 304.12 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 303.795 -0.845 304.125 -0.515 ;
        RECT 303.795 -2.205 304.125 -1.875 ;
        RECT 303.795 -3.565 304.125 -3.235 ;
        RECT 303.8 -3.565 304.12 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 303.795 -91.965 304.125 -91.635 ;
        RECT 303.795 -93.325 304.125 -92.995 ;
        RECT 303.795 -94.685 304.125 -94.355 ;
        RECT 303.795 -96.045 304.125 -95.715 ;
        RECT 303.795 -97.405 304.125 -97.075 ;
        RECT 303.795 -98.765 304.125 -98.435 ;
        RECT 303.795 -100.125 304.125 -99.795 ;
        RECT 303.795 -101.485 304.125 -101.155 ;
        RECT 303.795 -102.845 304.125 -102.515 ;
        RECT 303.795 -104.205 304.125 -103.875 ;
        RECT 303.795 -105.565 304.125 -105.235 ;
        RECT 303.795 -106.925 304.125 -106.595 ;
        RECT 303.795 -108.285 304.125 -107.955 ;
        RECT 303.795 -109.645 304.125 -109.315 ;
        RECT 303.795 -111.005 304.125 -110.675 ;
        RECT 303.795 -112.365 304.125 -112.035 ;
        RECT 303.795 -113.725 304.125 -113.395 ;
        RECT 303.795 -115.085 304.125 -114.755 ;
        RECT 303.795 -116.445 304.125 -116.115 ;
        RECT 303.795 -117.805 304.125 -117.475 ;
        RECT 303.795 -119.165 304.125 -118.835 ;
        RECT 303.795 -120.525 304.125 -120.195 ;
        RECT 303.795 -121.885 304.125 -121.555 ;
        RECT 303.795 -123.245 304.125 -122.915 ;
        RECT 303.795 -124.605 304.125 -124.275 ;
        RECT 303.795 -125.965 304.125 -125.635 ;
        RECT 303.795 -127.325 304.125 -126.995 ;
        RECT 303.795 -128.685 304.125 -128.355 ;
        RECT 303.795 -130.045 304.125 -129.715 ;
        RECT 303.795 -131.405 304.125 -131.075 ;
        RECT 303.795 -132.765 304.125 -132.435 ;
        RECT 303.795 -134.125 304.125 -133.795 ;
        RECT 303.795 -135.485 304.125 -135.155 ;
        RECT 303.795 -136.845 304.125 -136.515 ;
        RECT 303.795 -138.205 304.125 -137.875 ;
        RECT 303.795 -139.565 304.125 -139.235 ;
        RECT 303.795 -140.925 304.125 -140.595 ;
        RECT 303.795 -142.285 304.125 -141.955 ;
        RECT 303.795 -143.645 304.125 -143.315 ;
        RECT 303.795 -145.005 304.125 -144.675 ;
        RECT 303.795 -146.365 304.125 -146.035 ;
        RECT 303.795 -147.725 304.125 -147.395 ;
        RECT 303.795 -149.085 304.125 -148.755 ;
        RECT 303.795 -150.445 304.125 -150.115 ;
        RECT 303.795 -151.805 304.125 -151.475 ;
        RECT 303.795 -153.165 304.125 -152.835 ;
        RECT 303.795 -154.525 304.125 -154.195 ;
        RECT 303.795 -155.885 304.125 -155.555 ;
        RECT 303.795 -157.245 304.125 -156.915 ;
        RECT 303.795 -158.605 304.125 -158.275 ;
        RECT 303.795 -159.965 304.125 -159.635 ;
        RECT 303.795 -161.325 304.125 -160.995 ;
        RECT 303.795 -162.685 304.125 -162.355 ;
        RECT 303.795 -164.045 304.125 -163.715 ;
        RECT 303.795 -165.405 304.125 -165.075 ;
        RECT 303.795 -166.765 304.125 -166.435 ;
        RECT 303.795 -168.125 304.125 -167.795 ;
        RECT 303.795 -169.485 304.125 -169.155 ;
        RECT 303.795 -170.845 304.125 -170.515 ;
        RECT 303.795 -172.205 304.125 -171.875 ;
        RECT 303.795 -173.565 304.125 -173.235 ;
        RECT 303.795 -174.925 304.125 -174.595 ;
        RECT 303.795 -176.285 304.125 -175.955 ;
        RECT 303.795 -177.645 304.125 -177.315 ;
        RECT 303.795 -183.29 304.125 -182.16 ;
        RECT 303.8 -183.405 304.12 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 305.155 244.04 305.485 245.17 ;
        RECT 305.155 239.875 305.485 240.205 ;
        RECT 305.155 238.515 305.485 238.845 ;
        RECT 305.155 237.155 305.485 237.485 ;
        RECT 305.16 237.155 305.48 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 305.155 -0.845 305.485 -0.515 ;
        RECT 305.155 -2.205 305.485 -1.875 ;
        RECT 305.155 -3.565 305.485 -3.235 ;
        RECT 305.16 -3.565 305.48 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 306.515 244.04 306.845 245.17 ;
        RECT 306.515 239.875 306.845 240.205 ;
        RECT 306.515 238.515 306.845 238.845 ;
        RECT 306.515 237.155 306.845 237.485 ;
        RECT 306.52 237.155 306.84 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 234.46 -94.075 234.79 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 235.795 244.04 236.125 245.17 ;
        RECT 235.795 239.875 236.125 240.205 ;
        RECT 235.795 238.515 236.125 238.845 ;
        RECT 235.795 237.155 236.125 237.485 ;
        RECT 235.8 237.155 236.12 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 235.795 -0.845 236.125 -0.515 ;
        RECT 235.795 -2.205 236.125 -1.875 ;
        RECT 235.795 -3.565 236.125 -3.235 ;
        RECT 235.8 -3.565 236.12 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 237.155 244.04 237.485 245.17 ;
        RECT 237.155 239.875 237.485 240.205 ;
        RECT 237.155 238.515 237.485 238.845 ;
        RECT 237.155 237.155 237.485 237.485 ;
        RECT 237.16 237.155 237.48 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 237.155 -0.845 237.485 -0.515 ;
        RECT 237.155 -2.205 237.485 -1.875 ;
        RECT 237.155 -3.565 237.485 -3.235 ;
        RECT 237.16 -3.565 237.48 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 238.515 244.04 238.845 245.17 ;
        RECT 238.515 239.875 238.845 240.205 ;
        RECT 238.515 238.515 238.845 238.845 ;
        RECT 238.515 237.155 238.845 237.485 ;
        RECT 238.52 237.155 238.84 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 238.515 -0.845 238.845 -0.515 ;
        RECT 238.515 -2.205 238.845 -1.875 ;
        RECT 238.515 -3.565 238.845 -3.235 ;
        RECT 238.52 -3.565 238.84 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 238.515 -91.965 238.845 -91.635 ;
        RECT 238.515 -93.325 238.845 -92.995 ;
        RECT 238.515 -94.685 238.845 -94.355 ;
        RECT 238.515 -96.045 238.845 -95.715 ;
        RECT 238.515 -97.405 238.845 -97.075 ;
        RECT 238.515 -98.765 238.845 -98.435 ;
        RECT 238.515 -100.125 238.845 -99.795 ;
        RECT 238.515 -101.485 238.845 -101.155 ;
        RECT 238.515 -102.845 238.845 -102.515 ;
        RECT 238.515 -104.205 238.845 -103.875 ;
        RECT 238.515 -105.565 238.845 -105.235 ;
        RECT 238.515 -106.925 238.845 -106.595 ;
        RECT 238.515 -108.285 238.845 -107.955 ;
        RECT 238.515 -109.645 238.845 -109.315 ;
        RECT 238.515 -111.005 238.845 -110.675 ;
        RECT 238.515 -112.365 238.845 -112.035 ;
        RECT 238.515 -113.725 238.845 -113.395 ;
        RECT 238.515 -115.085 238.845 -114.755 ;
        RECT 238.515 -116.445 238.845 -116.115 ;
        RECT 238.515 -117.805 238.845 -117.475 ;
        RECT 238.515 -119.165 238.845 -118.835 ;
        RECT 238.515 -120.525 238.845 -120.195 ;
        RECT 238.515 -121.885 238.845 -121.555 ;
        RECT 238.515 -123.245 238.845 -122.915 ;
        RECT 238.515 -124.605 238.845 -124.275 ;
        RECT 238.515 -125.965 238.845 -125.635 ;
        RECT 238.515 -127.325 238.845 -126.995 ;
        RECT 238.515 -128.685 238.845 -128.355 ;
        RECT 238.515 -130.045 238.845 -129.715 ;
        RECT 238.515 -131.405 238.845 -131.075 ;
        RECT 238.515 -132.765 238.845 -132.435 ;
        RECT 238.515 -134.125 238.845 -133.795 ;
        RECT 238.515 -135.485 238.845 -135.155 ;
        RECT 238.515 -136.845 238.845 -136.515 ;
        RECT 238.515 -138.205 238.845 -137.875 ;
        RECT 238.515 -139.565 238.845 -139.235 ;
        RECT 238.515 -140.925 238.845 -140.595 ;
        RECT 238.515 -142.285 238.845 -141.955 ;
        RECT 238.515 -143.645 238.845 -143.315 ;
        RECT 238.515 -145.005 238.845 -144.675 ;
        RECT 238.515 -146.365 238.845 -146.035 ;
        RECT 238.515 -147.725 238.845 -147.395 ;
        RECT 238.515 -149.085 238.845 -148.755 ;
        RECT 238.515 -150.445 238.845 -150.115 ;
        RECT 238.515 -151.805 238.845 -151.475 ;
        RECT 238.515 -153.165 238.845 -152.835 ;
        RECT 238.515 -154.525 238.845 -154.195 ;
        RECT 238.515 -155.885 238.845 -155.555 ;
        RECT 238.515 -157.245 238.845 -156.915 ;
        RECT 238.515 -158.605 238.845 -158.275 ;
        RECT 238.515 -159.965 238.845 -159.635 ;
        RECT 238.515 -161.325 238.845 -160.995 ;
        RECT 238.515 -162.685 238.845 -162.355 ;
        RECT 238.515 -164.045 238.845 -163.715 ;
        RECT 238.515 -165.405 238.845 -165.075 ;
        RECT 238.515 -166.765 238.845 -166.435 ;
        RECT 238.515 -168.125 238.845 -167.795 ;
        RECT 238.515 -169.485 238.845 -169.155 ;
        RECT 238.515 -170.845 238.845 -170.515 ;
        RECT 238.515 -172.205 238.845 -171.875 ;
        RECT 238.515 -173.565 238.845 -173.235 ;
        RECT 238.515 -174.925 238.845 -174.595 ;
        RECT 238.515 -176.285 238.845 -175.955 ;
        RECT 238.515 -177.645 238.845 -177.315 ;
        RECT 238.515 -183.29 238.845 -182.16 ;
        RECT 238.52 -183.405 238.84 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 239.875 244.04 240.205 245.17 ;
        RECT 239.875 239.875 240.205 240.205 ;
        RECT 239.875 238.515 240.205 238.845 ;
        RECT 239.875 237.155 240.205 237.485 ;
        RECT 239.88 237.155 240.2 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 239.875 -0.845 240.205 -0.515 ;
        RECT 239.875 -2.205 240.205 -1.875 ;
        RECT 239.875 -3.565 240.205 -3.235 ;
        RECT 239.88 -3.565 240.2 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 239.875 -91.965 240.205 -91.635 ;
        RECT 239.875 -93.325 240.205 -92.995 ;
        RECT 239.875 -94.685 240.205 -94.355 ;
        RECT 239.875 -96.045 240.205 -95.715 ;
        RECT 239.875 -97.405 240.205 -97.075 ;
        RECT 239.875 -98.765 240.205 -98.435 ;
        RECT 239.875 -100.125 240.205 -99.795 ;
        RECT 239.875 -101.485 240.205 -101.155 ;
        RECT 239.875 -102.845 240.205 -102.515 ;
        RECT 239.875 -104.205 240.205 -103.875 ;
        RECT 239.875 -105.565 240.205 -105.235 ;
        RECT 239.875 -106.925 240.205 -106.595 ;
        RECT 239.875 -108.285 240.205 -107.955 ;
        RECT 239.875 -109.645 240.205 -109.315 ;
        RECT 239.875 -111.005 240.205 -110.675 ;
        RECT 239.875 -112.365 240.205 -112.035 ;
        RECT 239.875 -113.725 240.205 -113.395 ;
        RECT 239.875 -115.085 240.205 -114.755 ;
        RECT 239.875 -116.445 240.205 -116.115 ;
        RECT 239.875 -117.805 240.205 -117.475 ;
        RECT 239.875 -119.165 240.205 -118.835 ;
        RECT 239.875 -120.525 240.205 -120.195 ;
        RECT 239.875 -121.885 240.205 -121.555 ;
        RECT 239.875 -123.245 240.205 -122.915 ;
        RECT 239.875 -124.605 240.205 -124.275 ;
        RECT 239.875 -125.965 240.205 -125.635 ;
        RECT 239.875 -127.325 240.205 -126.995 ;
        RECT 239.875 -128.685 240.205 -128.355 ;
        RECT 239.875 -130.045 240.205 -129.715 ;
        RECT 239.875 -131.405 240.205 -131.075 ;
        RECT 239.875 -132.765 240.205 -132.435 ;
        RECT 239.875 -134.125 240.205 -133.795 ;
        RECT 239.875 -135.485 240.205 -135.155 ;
        RECT 239.875 -136.845 240.205 -136.515 ;
        RECT 239.875 -138.205 240.205 -137.875 ;
        RECT 239.875 -139.565 240.205 -139.235 ;
        RECT 239.875 -140.925 240.205 -140.595 ;
        RECT 239.875 -142.285 240.205 -141.955 ;
        RECT 239.875 -143.645 240.205 -143.315 ;
        RECT 239.875 -145.005 240.205 -144.675 ;
        RECT 239.875 -146.365 240.205 -146.035 ;
        RECT 239.875 -147.725 240.205 -147.395 ;
        RECT 239.875 -149.085 240.205 -148.755 ;
        RECT 239.875 -150.445 240.205 -150.115 ;
        RECT 239.875 -151.805 240.205 -151.475 ;
        RECT 239.875 -153.165 240.205 -152.835 ;
        RECT 239.875 -154.525 240.205 -154.195 ;
        RECT 239.875 -155.885 240.205 -155.555 ;
        RECT 239.875 -157.245 240.205 -156.915 ;
        RECT 239.875 -158.605 240.205 -158.275 ;
        RECT 239.875 -159.965 240.205 -159.635 ;
        RECT 239.875 -161.325 240.205 -160.995 ;
        RECT 239.875 -162.685 240.205 -162.355 ;
        RECT 239.875 -164.045 240.205 -163.715 ;
        RECT 239.875 -165.405 240.205 -165.075 ;
        RECT 239.875 -166.765 240.205 -166.435 ;
        RECT 239.875 -168.125 240.205 -167.795 ;
        RECT 239.875 -169.485 240.205 -169.155 ;
        RECT 239.875 -170.845 240.205 -170.515 ;
        RECT 239.875 -172.205 240.205 -171.875 ;
        RECT 239.875 -173.565 240.205 -173.235 ;
        RECT 239.875 -174.925 240.205 -174.595 ;
        RECT 239.875 -176.285 240.205 -175.955 ;
        RECT 239.875 -177.645 240.205 -177.315 ;
        RECT 239.875 -183.29 240.205 -182.16 ;
        RECT 239.88 -183.405 240.2 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 240.56 -94.075 240.89 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 241.235 244.04 241.565 245.17 ;
        RECT 241.235 239.875 241.565 240.205 ;
        RECT 241.235 238.515 241.565 238.845 ;
        RECT 241.235 237.155 241.565 237.485 ;
        RECT 241.24 237.155 241.56 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 242.595 244.04 242.925 245.17 ;
        RECT 242.595 239.875 242.925 240.205 ;
        RECT 242.595 238.515 242.925 238.845 ;
        RECT 242.595 237.155 242.925 237.485 ;
        RECT 242.6 237.155 242.92 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 242.595 -0.845 242.925 -0.515 ;
        RECT 242.595 -2.205 242.925 -1.875 ;
        RECT 242.595 -3.565 242.925 -3.235 ;
        RECT 242.6 -3.565 242.92 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 243.955 244.04 244.285 245.17 ;
        RECT 243.955 239.875 244.285 240.205 ;
        RECT 243.955 238.515 244.285 238.845 ;
        RECT 243.955 237.155 244.285 237.485 ;
        RECT 243.96 237.155 244.28 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 243.955 -0.845 244.285 -0.515 ;
        RECT 243.955 -2.205 244.285 -1.875 ;
        RECT 243.955 -3.565 244.285 -3.235 ;
        RECT 243.96 -3.565 244.28 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 245.315 244.04 245.645 245.17 ;
        RECT 245.315 239.875 245.645 240.205 ;
        RECT 245.315 238.515 245.645 238.845 ;
        RECT 245.315 237.155 245.645 237.485 ;
        RECT 245.32 237.155 245.64 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 245.315 -0.845 245.645 -0.515 ;
        RECT 245.315 -2.205 245.645 -1.875 ;
        RECT 245.315 -3.565 245.645 -3.235 ;
        RECT 245.32 -3.565 245.64 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 245.315 -91.965 245.645 -91.635 ;
        RECT 245.315 -93.325 245.645 -92.995 ;
        RECT 245.315 -94.685 245.645 -94.355 ;
        RECT 245.315 -96.045 245.645 -95.715 ;
        RECT 245.315 -97.405 245.645 -97.075 ;
        RECT 245.315 -98.765 245.645 -98.435 ;
        RECT 245.315 -100.125 245.645 -99.795 ;
        RECT 245.315 -101.485 245.645 -101.155 ;
        RECT 245.315 -102.845 245.645 -102.515 ;
        RECT 245.315 -104.205 245.645 -103.875 ;
        RECT 245.315 -105.565 245.645 -105.235 ;
        RECT 245.315 -106.925 245.645 -106.595 ;
        RECT 245.315 -108.285 245.645 -107.955 ;
        RECT 245.315 -109.645 245.645 -109.315 ;
        RECT 245.315 -111.005 245.645 -110.675 ;
        RECT 245.315 -112.365 245.645 -112.035 ;
        RECT 245.315 -113.725 245.645 -113.395 ;
        RECT 245.315 -115.085 245.645 -114.755 ;
        RECT 245.315 -116.445 245.645 -116.115 ;
        RECT 245.315 -117.805 245.645 -117.475 ;
        RECT 245.315 -119.165 245.645 -118.835 ;
        RECT 245.315 -120.525 245.645 -120.195 ;
        RECT 245.315 -121.885 245.645 -121.555 ;
        RECT 245.315 -123.245 245.645 -122.915 ;
        RECT 245.315 -124.605 245.645 -124.275 ;
        RECT 245.315 -125.965 245.645 -125.635 ;
        RECT 245.315 -127.325 245.645 -126.995 ;
        RECT 245.315 -128.685 245.645 -128.355 ;
        RECT 245.315 -130.045 245.645 -129.715 ;
        RECT 245.315 -131.405 245.645 -131.075 ;
        RECT 245.315 -132.765 245.645 -132.435 ;
        RECT 245.315 -134.125 245.645 -133.795 ;
        RECT 245.315 -135.485 245.645 -135.155 ;
        RECT 245.315 -136.845 245.645 -136.515 ;
        RECT 245.315 -138.205 245.645 -137.875 ;
        RECT 245.315 -139.565 245.645 -139.235 ;
        RECT 245.315 -140.925 245.645 -140.595 ;
        RECT 245.315 -142.285 245.645 -141.955 ;
        RECT 245.315 -143.645 245.645 -143.315 ;
        RECT 245.315 -145.005 245.645 -144.675 ;
        RECT 245.315 -146.365 245.645 -146.035 ;
        RECT 245.315 -147.725 245.645 -147.395 ;
        RECT 245.315 -149.085 245.645 -148.755 ;
        RECT 245.315 -150.445 245.645 -150.115 ;
        RECT 245.315 -151.805 245.645 -151.475 ;
        RECT 245.315 -153.165 245.645 -152.835 ;
        RECT 245.315 -154.525 245.645 -154.195 ;
        RECT 245.315 -155.885 245.645 -155.555 ;
        RECT 245.315 -157.245 245.645 -156.915 ;
        RECT 245.315 -158.605 245.645 -158.275 ;
        RECT 245.315 -159.965 245.645 -159.635 ;
        RECT 245.315 -161.325 245.645 -160.995 ;
        RECT 245.315 -162.685 245.645 -162.355 ;
        RECT 245.315 -164.045 245.645 -163.715 ;
        RECT 245.315 -165.405 245.645 -165.075 ;
        RECT 245.315 -166.765 245.645 -166.435 ;
        RECT 245.315 -168.125 245.645 -167.795 ;
        RECT 245.315 -169.485 245.645 -169.155 ;
        RECT 245.315 -170.845 245.645 -170.515 ;
        RECT 245.315 -172.205 245.645 -171.875 ;
        RECT 245.315 -173.565 245.645 -173.235 ;
        RECT 245.315 -174.925 245.645 -174.595 ;
        RECT 245.315 -176.285 245.645 -175.955 ;
        RECT 245.315 -177.645 245.645 -177.315 ;
        RECT 245.315 -183.29 245.645 -182.16 ;
        RECT 245.32 -183.405 245.64 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 246.66 -94.075 246.99 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 246.675 244.04 247.005 245.17 ;
        RECT 246.675 239.875 247.005 240.205 ;
        RECT 246.675 238.515 247.005 238.845 ;
        RECT 246.675 237.155 247.005 237.485 ;
        RECT 246.68 237.155 247 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 246.675 -96.045 247.005 -95.715 ;
        RECT 246.675 -97.405 247.005 -97.075 ;
        RECT 246.675 -98.765 247.005 -98.435 ;
        RECT 246.675 -100.125 247.005 -99.795 ;
        RECT 246.675 -101.485 247.005 -101.155 ;
        RECT 246.675 -102.845 247.005 -102.515 ;
        RECT 246.675 -104.205 247.005 -103.875 ;
        RECT 246.675 -105.565 247.005 -105.235 ;
        RECT 246.675 -106.925 247.005 -106.595 ;
        RECT 246.675 -108.285 247.005 -107.955 ;
        RECT 246.675 -109.645 247.005 -109.315 ;
        RECT 246.675 -111.005 247.005 -110.675 ;
        RECT 246.675 -112.365 247.005 -112.035 ;
        RECT 246.675 -113.725 247.005 -113.395 ;
        RECT 246.675 -115.085 247.005 -114.755 ;
        RECT 246.675 -116.445 247.005 -116.115 ;
        RECT 246.675 -117.805 247.005 -117.475 ;
        RECT 246.675 -119.165 247.005 -118.835 ;
        RECT 246.675 -120.525 247.005 -120.195 ;
        RECT 246.675 -121.885 247.005 -121.555 ;
        RECT 246.675 -123.245 247.005 -122.915 ;
        RECT 246.675 -124.605 247.005 -124.275 ;
        RECT 246.675 -125.965 247.005 -125.635 ;
        RECT 246.675 -127.325 247.005 -126.995 ;
        RECT 246.675 -128.685 247.005 -128.355 ;
        RECT 246.675 -130.045 247.005 -129.715 ;
        RECT 246.675 -131.405 247.005 -131.075 ;
        RECT 246.675 -132.765 247.005 -132.435 ;
        RECT 246.675 -134.125 247.005 -133.795 ;
        RECT 246.675 -135.485 247.005 -135.155 ;
        RECT 246.675 -136.845 247.005 -136.515 ;
        RECT 246.675 -138.205 247.005 -137.875 ;
        RECT 246.675 -139.565 247.005 -139.235 ;
        RECT 246.675 -140.925 247.005 -140.595 ;
        RECT 246.675 -142.285 247.005 -141.955 ;
        RECT 246.675 -143.645 247.005 -143.315 ;
        RECT 246.675 -145.005 247.005 -144.675 ;
        RECT 246.675 -146.365 247.005 -146.035 ;
        RECT 246.675 -147.725 247.005 -147.395 ;
        RECT 246.675 -149.085 247.005 -148.755 ;
        RECT 246.675 -150.445 247.005 -150.115 ;
        RECT 246.675 -151.805 247.005 -151.475 ;
        RECT 246.675 -153.165 247.005 -152.835 ;
        RECT 246.675 -154.525 247.005 -154.195 ;
        RECT 246.675 -155.885 247.005 -155.555 ;
        RECT 246.675 -157.245 247.005 -156.915 ;
        RECT 246.675 -158.605 247.005 -158.275 ;
        RECT 246.675 -159.965 247.005 -159.635 ;
        RECT 246.675 -161.325 247.005 -160.995 ;
        RECT 246.675 -162.685 247.005 -162.355 ;
        RECT 246.675 -164.045 247.005 -163.715 ;
        RECT 246.675 -165.405 247.005 -165.075 ;
        RECT 246.675 -166.765 247.005 -166.435 ;
        RECT 246.675 -168.125 247.005 -167.795 ;
        RECT 246.675 -169.485 247.005 -169.155 ;
        RECT 246.675 -170.845 247.005 -170.515 ;
        RECT 246.675 -172.205 247.005 -171.875 ;
        RECT 246.675 -173.565 247.005 -173.235 ;
        RECT 246.675 -174.925 247.005 -174.595 ;
        RECT 246.675 -176.285 247.005 -175.955 ;
        RECT 246.675 -177.645 247.005 -177.315 ;
        RECT 246.675 -183.29 247.005 -182.16 ;
        RECT 246.68 -183.405 247 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 248.035 244.04 248.365 245.17 ;
        RECT 248.035 239.875 248.365 240.205 ;
        RECT 248.035 238.515 248.365 238.845 ;
        RECT 248.035 237.155 248.365 237.485 ;
        RECT 248.04 237.155 248.36 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 248.035 -0.845 248.365 -0.515 ;
        RECT 248.035 -2.205 248.365 -1.875 ;
        RECT 248.035 -3.565 248.365 -3.235 ;
        RECT 248.04 -3.565 248.36 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 249.395 244.04 249.725 245.17 ;
        RECT 249.395 239.875 249.725 240.205 ;
        RECT 249.395 238.515 249.725 238.845 ;
        RECT 249.395 237.155 249.725 237.485 ;
        RECT 249.4 237.155 249.72 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 249.395 -0.845 249.725 -0.515 ;
        RECT 249.395 -2.205 249.725 -1.875 ;
        RECT 249.395 -3.565 249.725 -3.235 ;
        RECT 249.4 -3.565 249.72 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 250.755 244.04 251.085 245.17 ;
        RECT 250.755 239.875 251.085 240.205 ;
        RECT 250.755 238.515 251.085 238.845 ;
        RECT 250.755 237.155 251.085 237.485 ;
        RECT 250.76 237.155 251.08 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 250.755 -0.845 251.085 -0.515 ;
        RECT 250.755 -2.205 251.085 -1.875 ;
        RECT 250.755 -3.565 251.085 -3.235 ;
        RECT 250.76 -3.565 251.08 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 252.115 244.04 252.445 245.17 ;
        RECT 252.115 239.875 252.445 240.205 ;
        RECT 252.115 238.515 252.445 238.845 ;
        RECT 252.115 237.155 252.445 237.485 ;
        RECT 252.12 237.155 252.44 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 252.115 -96.045 252.445 -95.715 ;
        RECT 252.115 -97.405 252.445 -97.075 ;
        RECT 252.115 -98.765 252.445 -98.435 ;
        RECT 252.115 -100.125 252.445 -99.795 ;
        RECT 252.115 -101.485 252.445 -101.155 ;
        RECT 252.115 -102.845 252.445 -102.515 ;
        RECT 252.115 -104.205 252.445 -103.875 ;
        RECT 252.115 -105.565 252.445 -105.235 ;
        RECT 252.115 -106.925 252.445 -106.595 ;
        RECT 252.115 -108.285 252.445 -107.955 ;
        RECT 252.115 -109.645 252.445 -109.315 ;
        RECT 252.115 -111.005 252.445 -110.675 ;
        RECT 252.115 -112.365 252.445 -112.035 ;
        RECT 252.115 -113.725 252.445 -113.395 ;
        RECT 252.115 -115.085 252.445 -114.755 ;
        RECT 252.115 -116.445 252.445 -116.115 ;
        RECT 252.115 -117.805 252.445 -117.475 ;
        RECT 252.115 -119.165 252.445 -118.835 ;
        RECT 252.115 -120.525 252.445 -120.195 ;
        RECT 252.115 -121.885 252.445 -121.555 ;
        RECT 252.115 -123.245 252.445 -122.915 ;
        RECT 252.115 -124.605 252.445 -124.275 ;
        RECT 252.115 -125.965 252.445 -125.635 ;
        RECT 252.115 -127.325 252.445 -126.995 ;
        RECT 252.115 -128.685 252.445 -128.355 ;
        RECT 252.115 -130.045 252.445 -129.715 ;
        RECT 252.115 -131.405 252.445 -131.075 ;
        RECT 252.115 -132.765 252.445 -132.435 ;
        RECT 252.115 -134.125 252.445 -133.795 ;
        RECT 252.115 -135.485 252.445 -135.155 ;
        RECT 252.115 -136.845 252.445 -136.515 ;
        RECT 252.115 -138.205 252.445 -137.875 ;
        RECT 252.115 -139.565 252.445 -139.235 ;
        RECT 252.115 -140.925 252.445 -140.595 ;
        RECT 252.115 -142.285 252.445 -141.955 ;
        RECT 252.115 -143.645 252.445 -143.315 ;
        RECT 252.115 -145.005 252.445 -144.675 ;
        RECT 252.115 -146.365 252.445 -146.035 ;
        RECT 252.115 -147.725 252.445 -147.395 ;
        RECT 252.115 -149.085 252.445 -148.755 ;
        RECT 252.115 -150.445 252.445 -150.115 ;
        RECT 252.115 -151.805 252.445 -151.475 ;
        RECT 252.115 -153.165 252.445 -152.835 ;
        RECT 252.115 -154.525 252.445 -154.195 ;
        RECT 252.115 -155.885 252.445 -155.555 ;
        RECT 252.115 -157.245 252.445 -156.915 ;
        RECT 252.115 -158.605 252.445 -158.275 ;
        RECT 252.115 -159.965 252.445 -159.635 ;
        RECT 252.115 -161.325 252.445 -160.995 ;
        RECT 252.115 -162.685 252.445 -162.355 ;
        RECT 252.115 -164.045 252.445 -163.715 ;
        RECT 252.115 -165.405 252.445 -165.075 ;
        RECT 252.115 -166.765 252.445 -166.435 ;
        RECT 252.115 -168.125 252.445 -167.795 ;
        RECT 252.115 -169.485 252.445 -169.155 ;
        RECT 252.115 -170.845 252.445 -170.515 ;
        RECT 252.115 -172.205 252.445 -171.875 ;
        RECT 252.115 -173.565 252.445 -173.235 ;
        RECT 252.115 -174.925 252.445 -174.595 ;
        RECT 252.115 -176.285 252.445 -175.955 ;
        RECT 252.115 -177.645 252.445 -177.315 ;
        RECT 252.115 -183.29 252.445 -182.16 ;
        RECT 252.12 -183.405 252.44 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 252.76 -94.075 253.09 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 253.475 244.04 253.805 245.17 ;
        RECT 253.475 239.875 253.805 240.205 ;
        RECT 253.475 238.515 253.805 238.845 ;
        RECT 253.475 237.155 253.805 237.485 ;
        RECT 253.48 237.155 253.8 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 254.835 244.04 255.165 245.17 ;
        RECT 254.835 239.875 255.165 240.205 ;
        RECT 254.835 238.515 255.165 238.845 ;
        RECT 254.835 237.155 255.165 237.485 ;
        RECT 254.84 237.155 255.16 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 254.835 -0.845 255.165 -0.515 ;
        RECT 254.835 -2.205 255.165 -1.875 ;
        RECT 254.835 -3.565 255.165 -3.235 ;
        RECT 254.84 -3.565 255.16 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 256.195 244.04 256.525 245.17 ;
        RECT 256.195 239.875 256.525 240.205 ;
        RECT 256.195 238.515 256.525 238.845 ;
        RECT 256.195 237.155 256.525 237.485 ;
        RECT 256.2 237.155 256.52 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 256.195 -0.845 256.525 -0.515 ;
        RECT 256.195 -2.205 256.525 -1.875 ;
        RECT 256.195 -3.565 256.525 -3.235 ;
        RECT 256.2 -3.565 256.52 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 257.555 244.04 257.885 245.17 ;
        RECT 257.555 239.875 257.885 240.205 ;
        RECT 257.555 238.515 257.885 238.845 ;
        RECT 257.555 237.155 257.885 237.485 ;
        RECT 257.56 237.155 257.88 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 257.555 -0.845 257.885 -0.515 ;
        RECT 257.555 -2.205 257.885 -1.875 ;
        RECT 257.555 -3.565 257.885 -3.235 ;
        RECT 257.56 -3.565 257.88 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 257.555 -91.965 257.885 -91.635 ;
        RECT 257.555 -93.325 257.885 -92.995 ;
        RECT 257.555 -94.685 257.885 -94.355 ;
        RECT 257.555 -96.045 257.885 -95.715 ;
        RECT 257.555 -97.405 257.885 -97.075 ;
        RECT 257.555 -98.765 257.885 -98.435 ;
        RECT 257.555 -100.125 257.885 -99.795 ;
        RECT 257.555 -101.485 257.885 -101.155 ;
        RECT 257.555 -102.845 257.885 -102.515 ;
        RECT 257.555 -104.205 257.885 -103.875 ;
        RECT 257.555 -105.565 257.885 -105.235 ;
        RECT 257.555 -106.925 257.885 -106.595 ;
        RECT 257.555 -108.285 257.885 -107.955 ;
        RECT 257.555 -109.645 257.885 -109.315 ;
        RECT 257.555 -111.005 257.885 -110.675 ;
        RECT 257.555 -112.365 257.885 -112.035 ;
        RECT 257.555 -113.725 257.885 -113.395 ;
        RECT 257.555 -115.085 257.885 -114.755 ;
        RECT 257.555 -116.445 257.885 -116.115 ;
        RECT 257.555 -117.805 257.885 -117.475 ;
        RECT 257.555 -119.165 257.885 -118.835 ;
        RECT 257.555 -120.525 257.885 -120.195 ;
        RECT 257.555 -121.885 257.885 -121.555 ;
        RECT 257.555 -123.245 257.885 -122.915 ;
        RECT 257.555 -124.605 257.885 -124.275 ;
        RECT 257.555 -125.965 257.885 -125.635 ;
        RECT 257.555 -127.325 257.885 -126.995 ;
        RECT 257.555 -128.685 257.885 -128.355 ;
        RECT 257.555 -130.045 257.885 -129.715 ;
        RECT 257.555 -131.405 257.885 -131.075 ;
        RECT 257.555 -132.765 257.885 -132.435 ;
        RECT 257.555 -134.125 257.885 -133.795 ;
        RECT 257.555 -135.485 257.885 -135.155 ;
        RECT 257.555 -136.845 257.885 -136.515 ;
        RECT 257.555 -138.205 257.885 -137.875 ;
        RECT 257.555 -139.565 257.885 -139.235 ;
        RECT 257.555 -140.925 257.885 -140.595 ;
        RECT 257.555 -142.285 257.885 -141.955 ;
        RECT 257.555 -143.645 257.885 -143.315 ;
        RECT 257.555 -145.005 257.885 -144.675 ;
        RECT 257.555 -146.365 257.885 -146.035 ;
        RECT 257.555 -147.725 257.885 -147.395 ;
        RECT 257.555 -149.085 257.885 -148.755 ;
        RECT 257.555 -150.445 257.885 -150.115 ;
        RECT 257.555 -151.805 257.885 -151.475 ;
        RECT 257.555 -153.165 257.885 -152.835 ;
        RECT 257.555 -154.525 257.885 -154.195 ;
        RECT 257.555 -155.885 257.885 -155.555 ;
        RECT 257.555 -157.245 257.885 -156.915 ;
        RECT 257.555 -158.605 257.885 -158.275 ;
        RECT 257.555 -159.965 257.885 -159.635 ;
        RECT 257.555 -161.325 257.885 -160.995 ;
        RECT 257.555 -162.685 257.885 -162.355 ;
        RECT 257.555 -164.045 257.885 -163.715 ;
        RECT 257.555 -165.405 257.885 -165.075 ;
        RECT 257.555 -166.765 257.885 -166.435 ;
        RECT 257.555 -168.125 257.885 -167.795 ;
        RECT 257.555 -169.485 257.885 -169.155 ;
        RECT 257.555 -170.845 257.885 -170.515 ;
        RECT 257.555 -172.205 257.885 -171.875 ;
        RECT 257.555 -173.565 257.885 -173.235 ;
        RECT 257.555 -174.925 257.885 -174.595 ;
        RECT 257.555 -176.285 257.885 -175.955 ;
        RECT 257.555 -177.645 257.885 -177.315 ;
        RECT 257.555 -183.29 257.885 -182.16 ;
        RECT 257.56 -183.405 257.88 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 258.86 -94.075 259.19 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 258.915 244.04 259.245 245.17 ;
        RECT 258.915 239.875 259.245 240.205 ;
        RECT 258.915 238.515 259.245 238.845 ;
        RECT 258.915 237.155 259.245 237.485 ;
        RECT 258.92 237.155 259.24 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 258.915 -96.045 259.245 -95.715 ;
        RECT 258.915 -97.405 259.245 -97.075 ;
        RECT 258.915 -98.765 259.245 -98.435 ;
        RECT 258.915 -100.125 259.245 -99.795 ;
        RECT 258.915 -101.485 259.245 -101.155 ;
        RECT 258.915 -102.845 259.245 -102.515 ;
        RECT 258.915 -104.205 259.245 -103.875 ;
        RECT 258.915 -105.565 259.245 -105.235 ;
        RECT 258.915 -106.925 259.245 -106.595 ;
        RECT 258.915 -108.285 259.245 -107.955 ;
        RECT 258.915 -109.645 259.245 -109.315 ;
        RECT 258.915 -111.005 259.245 -110.675 ;
        RECT 258.915 -112.365 259.245 -112.035 ;
        RECT 258.915 -113.725 259.245 -113.395 ;
        RECT 258.915 -115.085 259.245 -114.755 ;
        RECT 258.915 -116.445 259.245 -116.115 ;
        RECT 258.915 -117.805 259.245 -117.475 ;
        RECT 258.915 -119.165 259.245 -118.835 ;
        RECT 258.915 -120.525 259.245 -120.195 ;
        RECT 258.915 -121.885 259.245 -121.555 ;
        RECT 258.915 -123.245 259.245 -122.915 ;
        RECT 258.915 -124.605 259.245 -124.275 ;
        RECT 258.915 -125.965 259.245 -125.635 ;
        RECT 258.915 -127.325 259.245 -126.995 ;
        RECT 258.915 -128.685 259.245 -128.355 ;
        RECT 258.915 -130.045 259.245 -129.715 ;
        RECT 258.915 -131.405 259.245 -131.075 ;
        RECT 258.915 -132.765 259.245 -132.435 ;
        RECT 258.915 -134.125 259.245 -133.795 ;
        RECT 258.915 -135.485 259.245 -135.155 ;
        RECT 258.915 -136.845 259.245 -136.515 ;
        RECT 258.915 -138.205 259.245 -137.875 ;
        RECT 258.915 -139.565 259.245 -139.235 ;
        RECT 258.915 -140.925 259.245 -140.595 ;
        RECT 258.915 -142.285 259.245 -141.955 ;
        RECT 258.915 -143.645 259.245 -143.315 ;
        RECT 258.915 -145.005 259.245 -144.675 ;
        RECT 258.915 -146.365 259.245 -146.035 ;
        RECT 258.915 -147.725 259.245 -147.395 ;
        RECT 258.915 -149.085 259.245 -148.755 ;
        RECT 258.915 -150.445 259.245 -150.115 ;
        RECT 258.915 -151.805 259.245 -151.475 ;
        RECT 258.915 -153.165 259.245 -152.835 ;
        RECT 258.915 -154.525 259.245 -154.195 ;
        RECT 258.915 -155.885 259.245 -155.555 ;
        RECT 258.915 -157.245 259.245 -156.915 ;
        RECT 258.915 -158.605 259.245 -158.275 ;
        RECT 258.915 -159.965 259.245 -159.635 ;
        RECT 258.915 -161.325 259.245 -160.995 ;
        RECT 258.915 -162.685 259.245 -162.355 ;
        RECT 258.915 -164.045 259.245 -163.715 ;
        RECT 258.915 -165.405 259.245 -165.075 ;
        RECT 258.915 -166.765 259.245 -166.435 ;
        RECT 258.915 -168.125 259.245 -167.795 ;
        RECT 258.915 -169.485 259.245 -169.155 ;
        RECT 258.915 -170.845 259.245 -170.515 ;
        RECT 258.915 -172.205 259.245 -171.875 ;
        RECT 258.915 -173.565 259.245 -173.235 ;
        RECT 258.915 -174.925 259.245 -174.595 ;
        RECT 258.915 -176.285 259.245 -175.955 ;
        RECT 258.915 -177.645 259.245 -177.315 ;
        RECT 258.915 -183.29 259.245 -182.16 ;
        RECT 258.92 -183.405 259.24 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 260.275 244.04 260.605 245.17 ;
        RECT 260.275 239.875 260.605 240.205 ;
        RECT 260.275 238.515 260.605 238.845 ;
        RECT 260.275 237.155 260.605 237.485 ;
        RECT 260.28 237.155 260.6 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 260.275 -0.845 260.605 -0.515 ;
        RECT 260.275 -2.205 260.605 -1.875 ;
        RECT 260.275 -3.565 260.605 -3.235 ;
        RECT 260.28 -3.565 260.6 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 261.635 244.04 261.965 245.17 ;
        RECT 261.635 239.875 261.965 240.205 ;
        RECT 261.635 238.515 261.965 238.845 ;
        RECT 261.635 237.155 261.965 237.485 ;
        RECT 261.64 237.155 261.96 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 261.635 -0.845 261.965 -0.515 ;
        RECT 261.635 -2.205 261.965 -1.875 ;
        RECT 261.635 -3.565 261.965 -3.235 ;
        RECT 261.64 -3.565 261.96 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 262.995 244.04 263.325 245.17 ;
        RECT 262.995 239.875 263.325 240.205 ;
        RECT 262.995 238.515 263.325 238.845 ;
        RECT 262.995 237.155 263.325 237.485 ;
        RECT 263 237.155 263.32 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 262.995 -0.845 263.325 -0.515 ;
        RECT 262.995 -2.205 263.325 -1.875 ;
        RECT 262.995 -3.565 263.325 -3.235 ;
        RECT 263 -3.565 263.32 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 262.995 -91.965 263.325 -91.635 ;
        RECT 262.995 -93.325 263.325 -92.995 ;
        RECT 262.995 -94.685 263.325 -94.355 ;
        RECT 262.995 -96.045 263.325 -95.715 ;
        RECT 262.995 -97.405 263.325 -97.075 ;
        RECT 262.995 -98.765 263.325 -98.435 ;
        RECT 262.995 -100.125 263.325 -99.795 ;
        RECT 262.995 -101.485 263.325 -101.155 ;
        RECT 262.995 -102.845 263.325 -102.515 ;
        RECT 262.995 -104.205 263.325 -103.875 ;
        RECT 262.995 -105.565 263.325 -105.235 ;
        RECT 262.995 -106.925 263.325 -106.595 ;
        RECT 262.995 -108.285 263.325 -107.955 ;
        RECT 262.995 -109.645 263.325 -109.315 ;
        RECT 262.995 -111.005 263.325 -110.675 ;
        RECT 262.995 -112.365 263.325 -112.035 ;
        RECT 262.995 -113.725 263.325 -113.395 ;
        RECT 262.995 -115.085 263.325 -114.755 ;
        RECT 262.995 -116.445 263.325 -116.115 ;
        RECT 262.995 -117.805 263.325 -117.475 ;
        RECT 262.995 -119.165 263.325 -118.835 ;
        RECT 262.995 -120.525 263.325 -120.195 ;
        RECT 262.995 -121.885 263.325 -121.555 ;
        RECT 262.995 -123.245 263.325 -122.915 ;
        RECT 262.995 -124.605 263.325 -124.275 ;
        RECT 262.995 -125.965 263.325 -125.635 ;
        RECT 262.995 -127.325 263.325 -126.995 ;
        RECT 262.995 -128.685 263.325 -128.355 ;
        RECT 262.995 -130.045 263.325 -129.715 ;
        RECT 262.995 -131.405 263.325 -131.075 ;
        RECT 262.995 -132.765 263.325 -132.435 ;
        RECT 262.995 -134.125 263.325 -133.795 ;
        RECT 262.995 -135.485 263.325 -135.155 ;
        RECT 262.995 -136.845 263.325 -136.515 ;
        RECT 262.995 -138.205 263.325 -137.875 ;
        RECT 262.995 -139.565 263.325 -139.235 ;
        RECT 262.995 -140.925 263.325 -140.595 ;
        RECT 262.995 -142.285 263.325 -141.955 ;
        RECT 262.995 -143.645 263.325 -143.315 ;
        RECT 262.995 -145.005 263.325 -144.675 ;
        RECT 262.995 -146.365 263.325 -146.035 ;
        RECT 262.995 -147.725 263.325 -147.395 ;
        RECT 262.995 -149.085 263.325 -148.755 ;
        RECT 262.995 -150.445 263.325 -150.115 ;
        RECT 262.995 -151.805 263.325 -151.475 ;
        RECT 262.995 -153.165 263.325 -152.835 ;
        RECT 262.995 -154.525 263.325 -154.195 ;
        RECT 262.995 -155.885 263.325 -155.555 ;
        RECT 262.995 -157.245 263.325 -156.915 ;
        RECT 262.995 -158.605 263.325 -158.275 ;
        RECT 262.995 -159.965 263.325 -159.635 ;
        RECT 262.995 -161.325 263.325 -160.995 ;
        RECT 262.995 -162.685 263.325 -162.355 ;
        RECT 262.995 -164.045 263.325 -163.715 ;
        RECT 262.995 -165.405 263.325 -165.075 ;
        RECT 262.995 -166.765 263.325 -166.435 ;
        RECT 262.995 -168.125 263.325 -167.795 ;
        RECT 262.995 -169.485 263.325 -169.155 ;
        RECT 262.995 -170.845 263.325 -170.515 ;
        RECT 262.995 -172.205 263.325 -171.875 ;
        RECT 262.995 -173.565 263.325 -173.235 ;
        RECT 262.995 -174.925 263.325 -174.595 ;
        RECT 262.995 -176.285 263.325 -175.955 ;
        RECT 262.995 -177.645 263.325 -177.315 ;
        RECT 262.995 -183.29 263.325 -182.16 ;
        RECT 263 -183.405 263.32 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 264.355 244.04 264.685 245.17 ;
        RECT 264.355 239.875 264.685 240.205 ;
        RECT 264.355 238.515 264.685 238.845 ;
        RECT 264.355 237.155 264.685 237.485 ;
        RECT 264.36 237.155 264.68 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 264.355 -96.045 264.685 -95.715 ;
        RECT 264.355 -97.405 264.685 -97.075 ;
        RECT 264.355 -98.765 264.685 -98.435 ;
        RECT 264.355 -100.125 264.685 -99.795 ;
        RECT 264.355 -101.485 264.685 -101.155 ;
        RECT 264.355 -102.845 264.685 -102.515 ;
        RECT 264.355 -104.205 264.685 -103.875 ;
        RECT 264.355 -105.565 264.685 -105.235 ;
        RECT 264.355 -106.925 264.685 -106.595 ;
        RECT 264.355 -108.285 264.685 -107.955 ;
        RECT 264.355 -109.645 264.685 -109.315 ;
        RECT 264.355 -111.005 264.685 -110.675 ;
        RECT 264.355 -112.365 264.685 -112.035 ;
        RECT 264.355 -113.725 264.685 -113.395 ;
        RECT 264.355 -115.085 264.685 -114.755 ;
        RECT 264.355 -116.445 264.685 -116.115 ;
        RECT 264.355 -117.805 264.685 -117.475 ;
        RECT 264.355 -119.165 264.685 -118.835 ;
        RECT 264.355 -120.525 264.685 -120.195 ;
        RECT 264.355 -121.885 264.685 -121.555 ;
        RECT 264.355 -123.245 264.685 -122.915 ;
        RECT 264.355 -124.605 264.685 -124.275 ;
        RECT 264.355 -125.965 264.685 -125.635 ;
        RECT 264.355 -127.325 264.685 -126.995 ;
        RECT 264.355 -128.685 264.685 -128.355 ;
        RECT 264.355 -130.045 264.685 -129.715 ;
        RECT 264.355 -131.405 264.685 -131.075 ;
        RECT 264.355 -132.765 264.685 -132.435 ;
        RECT 264.355 -134.125 264.685 -133.795 ;
        RECT 264.355 -135.485 264.685 -135.155 ;
        RECT 264.355 -136.845 264.685 -136.515 ;
        RECT 264.355 -138.205 264.685 -137.875 ;
        RECT 264.355 -139.565 264.685 -139.235 ;
        RECT 264.355 -140.925 264.685 -140.595 ;
        RECT 264.355 -142.285 264.685 -141.955 ;
        RECT 264.355 -143.645 264.685 -143.315 ;
        RECT 264.355 -145.005 264.685 -144.675 ;
        RECT 264.355 -146.365 264.685 -146.035 ;
        RECT 264.355 -147.725 264.685 -147.395 ;
        RECT 264.355 -149.085 264.685 -148.755 ;
        RECT 264.355 -150.445 264.685 -150.115 ;
        RECT 264.355 -151.805 264.685 -151.475 ;
        RECT 264.355 -153.165 264.685 -152.835 ;
        RECT 264.355 -154.525 264.685 -154.195 ;
        RECT 264.355 -155.885 264.685 -155.555 ;
        RECT 264.355 -157.245 264.685 -156.915 ;
        RECT 264.355 -158.605 264.685 -158.275 ;
        RECT 264.355 -159.965 264.685 -159.635 ;
        RECT 264.355 -161.325 264.685 -160.995 ;
        RECT 264.355 -162.685 264.685 -162.355 ;
        RECT 264.355 -164.045 264.685 -163.715 ;
        RECT 264.355 -165.405 264.685 -165.075 ;
        RECT 264.355 -166.765 264.685 -166.435 ;
        RECT 264.355 -168.125 264.685 -167.795 ;
        RECT 264.355 -169.485 264.685 -169.155 ;
        RECT 264.355 -170.845 264.685 -170.515 ;
        RECT 264.355 -172.205 264.685 -171.875 ;
        RECT 264.355 -173.565 264.685 -173.235 ;
        RECT 264.355 -174.925 264.685 -174.595 ;
        RECT 264.355 -176.285 264.685 -175.955 ;
        RECT 264.355 -177.645 264.685 -177.315 ;
        RECT 264.355 -183.29 264.685 -182.16 ;
        RECT 264.36 -183.405 264.68 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 264.96 -94.075 265.29 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 265.715 244.04 266.045 245.17 ;
        RECT 265.715 239.875 266.045 240.205 ;
        RECT 265.715 238.515 266.045 238.845 ;
        RECT 265.715 237.155 266.045 237.485 ;
        RECT 265.72 237.155 266.04 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 267.075 244.04 267.405 245.17 ;
        RECT 267.075 239.875 267.405 240.205 ;
        RECT 267.075 238.515 267.405 238.845 ;
        RECT 267.075 237.155 267.405 237.485 ;
        RECT 267.08 237.155 267.4 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 267.075 -0.845 267.405 -0.515 ;
        RECT 267.075 -2.205 267.405 -1.875 ;
        RECT 267.075 -3.565 267.405 -3.235 ;
        RECT 267.08 -3.565 267.4 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 267.075 -91.965 267.405 -91.635 ;
        RECT 267.075 -93.325 267.405 -92.995 ;
        RECT 267.075 -94.685 267.405 -94.355 ;
        RECT 267.075 -96.045 267.405 -95.715 ;
        RECT 267.075 -97.405 267.405 -97.075 ;
        RECT 267.075 -98.765 267.405 -98.435 ;
        RECT 267.075 -100.125 267.405 -99.795 ;
        RECT 267.075 -101.485 267.405 -101.155 ;
        RECT 267.075 -102.845 267.405 -102.515 ;
        RECT 267.075 -104.205 267.405 -103.875 ;
        RECT 267.075 -105.565 267.405 -105.235 ;
        RECT 267.075 -106.925 267.405 -106.595 ;
        RECT 267.075 -108.285 267.405 -107.955 ;
        RECT 267.075 -109.645 267.405 -109.315 ;
        RECT 267.075 -111.005 267.405 -110.675 ;
        RECT 267.075 -112.365 267.405 -112.035 ;
        RECT 267.075 -113.725 267.405 -113.395 ;
        RECT 267.075 -115.085 267.405 -114.755 ;
        RECT 267.075 -116.445 267.405 -116.115 ;
        RECT 267.075 -117.805 267.405 -117.475 ;
        RECT 267.075 -119.165 267.405 -118.835 ;
        RECT 267.075 -120.525 267.405 -120.195 ;
        RECT 267.075 -121.885 267.405 -121.555 ;
        RECT 267.075 -123.245 267.405 -122.915 ;
        RECT 267.075 -124.605 267.405 -124.275 ;
        RECT 267.075 -125.965 267.405 -125.635 ;
        RECT 267.075 -127.325 267.405 -126.995 ;
        RECT 267.075 -128.685 267.405 -128.355 ;
        RECT 267.075 -130.045 267.405 -129.715 ;
        RECT 267.075 -131.405 267.405 -131.075 ;
        RECT 267.075 -132.765 267.405 -132.435 ;
        RECT 267.075 -134.125 267.405 -133.795 ;
        RECT 267.075 -135.485 267.405 -135.155 ;
        RECT 267.075 -136.845 267.405 -136.515 ;
        RECT 267.075 -138.205 267.405 -137.875 ;
        RECT 267.075 -139.565 267.405 -139.235 ;
        RECT 267.075 -140.925 267.405 -140.595 ;
        RECT 267.075 -142.285 267.405 -141.955 ;
        RECT 267.075 -143.645 267.405 -143.315 ;
        RECT 267.075 -145.005 267.405 -144.675 ;
        RECT 267.075 -146.365 267.405 -146.035 ;
        RECT 267.075 -147.725 267.405 -147.395 ;
        RECT 267.075 -149.085 267.405 -148.755 ;
        RECT 267.075 -150.445 267.405 -150.115 ;
        RECT 267.075 -151.805 267.405 -151.475 ;
        RECT 267.075 -153.165 267.405 -152.835 ;
        RECT 267.075 -154.525 267.405 -154.195 ;
        RECT 267.075 -155.885 267.405 -155.555 ;
        RECT 267.075 -157.245 267.405 -156.915 ;
        RECT 267.075 -158.605 267.405 -158.275 ;
        RECT 267.075 -159.965 267.405 -159.635 ;
        RECT 267.075 -161.325 267.405 -160.995 ;
        RECT 267.075 -162.685 267.405 -162.355 ;
        RECT 267.075 -164.045 267.405 -163.715 ;
        RECT 267.075 -165.405 267.405 -165.075 ;
        RECT 267.075 -166.765 267.405 -166.435 ;
        RECT 267.075 -168.125 267.405 -167.795 ;
        RECT 267.075 -169.485 267.405 -169.155 ;
        RECT 267.075 -170.845 267.405 -170.515 ;
        RECT 267.075 -172.205 267.405 -171.875 ;
        RECT 267.075 -173.565 267.405 -173.235 ;
        RECT 267.075 -174.925 267.405 -174.595 ;
        RECT 267.075 -176.285 267.405 -175.955 ;
        RECT 267.075 -177.645 267.405 -177.315 ;
        RECT 267.075 -183.29 267.405 -182.16 ;
        RECT 267.08 -183.405 267.4 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 268.435 244.04 268.765 245.17 ;
        RECT 268.435 239.875 268.765 240.205 ;
        RECT 268.435 238.515 268.765 238.845 ;
        RECT 268.435 237.155 268.765 237.485 ;
        RECT 268.44 237.155 268.76 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 268.435 -0.845 268.765 -0.515 ;
        RECT 268.435 -2.205 268.765 -1.875 ;
        RECT 268.435 -3.565 268.765 -3.235 ;
        RECT 268.44 -3.565 268.76 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 269.795 244.04 270.125 245.17 ;
        RECT 269.795 239.875 270.125 240.205 ;
        RECT 269.795 238.515 270.125 238.845 ;
        RECT 269.795 237.155 270.125 237.485 ;
        RECT 269.8 237.155 270.12 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 269.795 -0.845 270.125 -0.515 ;
        RECT 269.795 -2.205 270.125 -1.875 ;
        RECT 269.795 -3.565 270.125 -3.235 ;
        RECT 269.8 -3.565 270.12 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 269.795 -91.965 270.125 -91.635 ;
        RECT 269.795 -93.325 270.125 -92.995 ;
        RECT 269.795 -94.685 270.125 -94.355 ;
        RECT 269.795 -96.045 270.125 -95.715 ;
        RECT 269.795 -97.405 270.125 -97.075 ;
        RECT 269.795 -98.765 270.125 -98.435 ;
        RECT 269.795 -100.125 270.125 -99.795 ;
        RECT 269.795 -101.485 270.125 -101.155 ;
        RECT 269.795 -102.845 270.125 -102.515 ;
        RECT 269.795 -104.205 270.125 -103.875 ;
        RECT 269.795 -105.565 270.125 -105.235 ;
        RECT 269.795 -106.925 270.125 -106.595 ;
        RECT 269.795 -108.285 270.125 -107.955 ;
        RECT 269.795 -109.645 270.125 -109.315 ;
        RECT 269.795 -111.005 270.125 -110.675 ;
        RECT 269.795 -112.365 270.125 -112.035 ;
        RECT 269.795 -113.725 270.125 -113.395 ;
        RECT 269.795 -115.085 270.125 -114.755 ;
        RECT 269.795 -116.445 270.125 -116.115 ;
        RECT 269.795 -117.805 270.125 -117.475 ;
        RECT 269.795 -119.165 270.125 -118.835 ;
        RECT 269.795 -120.525 270.125 -120.195 ;
        RECT 269.795 -121.885 270.125 -121.555 ;
        RECT 269.795 -123.245 270.125 -122.915 ;
        RECT 269.795 -124.605 270.125 -124.275 ;
        RECT 269.795 -125.965 270.125 -125.635 ;
        RECT 269.795 -127.325 270.125 -126.995 ;
        RECT 269.795 -128.685 270.125 -128.355 ;
        RECT 269.795 -130.045 270.125 -129.715 ;
        RECT 269.795 -131.405 270.125 -131.075 ;
        RECT 269.795 -132.765 270.125 -132.435 ;
        RECT 269.795 -134.125 270.125 -133.795 ;
        RECT 269.795 -135.485 270.125 -135.155 ;
        RECT 269.795 -136.845 270.125 -136.515 ;
        RECT 269.795 -138.205 270.125 -137.875 ;
        RECT 269.795 -139.565 270.125 -139.235 ;
        RECT 269.795 -140.925 270.125 -140.595 ;
        RECT 269.795 -142.285 270.125 -141.955 ;
        RECT 269.795 -143.645 270.125 -143.315 ;
        RECT 269.795 -145.005 270.125 -144.675 ;
        RECT 269.795 -146.365 270.125 -146.035 ;
        RECT 269.795 -147.725 270.125 -147.395 ;
        RECT 269.795 -149.085 270.125 -148.755 ;
        RECT 269.795 -150.445 270.125 -150.115 ;
        RECT 269.795 -151.805 270.125 -151.475 ;
        RECT 269.795 -153.165 270.125 -152.835 ;
        RECT 269.795 -154.525 270.125 -154.195 ;
        RECT 269.795 -155.885 270.125 -155.555 ;
        RECT 269.795 -157.245 270.125 -156.915 ;
        RECT 269.795 -158.605 270.125 -158.275 ;
        RECT 269.795 -159.965 270.125 -159.635 ;
        RECT 269.795 -161.325 270.125 -160.995 ;
        RECT 269.795 -162.685 270.125 -162.355 ;
        RECT 269.795 -164.045 270.125 -163.715 ;
        RECT 269.795 -165.405 270.125 -165.075 ;
        RECT 269.795 -166.765 270.125 -166.435 ;
        RECT 269.795 -168.125 270.125 -167.795 ;
        RECT 269.795 -169.485 270.125 -169.155 ;
        RECT 269.795 -170.845 270.125 -170.515 ;
        RECT 269.795 -172.205 270.125 -171.875 ;
        RECT 269.795 -173.565 270.125 -173.235 ;
        RECT 269.795 -174.925 270.125 -174.595 ;
        RECT 269.795 -176.285 270.125 -175.955 ;
        RECT 269.795 -177.645 270.125 -177.315 ;
        RECT 269.795 -183.29 270.125 -182.16 ;
        RECT 269.8 -183.405 270.12 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 271.06 -94.075 271.39 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 271.155 244.04 271.485 245.17 ;
        RECT 271.155 239.875 271.485 240.205 ;
        RECT 271.155 238.515 271.485 238.845 ;
        RECT 271.155 237.155 271.485 237.485 ;
        RECT 271.16 237.155 271.48 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 271.155 -123.245 271.485 -122.915 ;
        RECT 271.155 -124.605 271.485 -124.275 ;
        RECT 271.155 -125.965 271.485 -125.635 ;
        RECT 271.155 -127.325 271.485 -126.995 ;
        RECT 271.155 -128.685 271.485 -128.355 ;
        RECT 271.155 -130.045 271.485 -129.715 ;
        RECT 271.155 -131.405 271.485 -131.075 ;
        RECT 271.155 -132.765 271.485 -132.435 ;
        RECT 271.155 -134.125 271.485 -133.795 ;
        RECT 271.155 -135.485 271.485 -135.155 ;
        RECT 271.155 -136.845 271.485 -136.515 ;
        RECT 271.155 -138.205 271.485 -137.875 ;
        RECT 271.155 -139.565 271.485 -139.235 ;
        RECT 271.155 -140.925 271.485 -140.595 ;
        RECT 271.155 -142.285 271.485 -141.955 ;
        RECT 271.155 -143.645 271.485 -143.315 ;
        RECT 271.155 -145.005 271.485 -144.675 ;
        RECT 271.155 -146.365 271.485 -146.035 ;
        RECT 271.155 -147.725 271.485 -147.395 ;
        RECT 271.155 -149.085 271.485 -148.755 ;
        RECT 271.155 -150.445 271.485 -150.115 ;
        RECT 271.155 -151.805 271.485 -151.475 ;
        RECT 271.155 -153.165 271.485 -152.835 ;
        RECT 271.155 -154.525 271.485 -154.195 ;
        RECT 271.155 -155.885 271.485 -155.555 ;
        RECT 271.155 -157.245 271.485 -156.915 ;
        RECT 271.155 -158.605 271.485 -158.275 ;
        RECT 271.155 -159.965 271.485 -159.635 ;
        RECT 271.155 -161.325 271.485 -160.995 ;
        RECT 271.155 -162.685 271.485 -162.355 ;
        RECT 271.155 -164.045 271.485 -163.715 ;
        RECT 271.155 -165.405 271.485 -165.075 ;
        RECT 271.155 -166.765 271.485 -166.435 ;
        RECT 271.155 -168.125 271.485 -167.795 ;
        RECT 271.155 -169.485 271.485 -169.155 ;
        RECT 271.155 -170.845 271.485 -170.515 ;
        RECT 271.155 -172.205 271.485 -171.875 ;
        RECT 271.155 -173.565 271.485 -173.235 ;
        RECT 271.155 -174.925 271.485 -174.595 ;
        RECT 271.155 -176.285 271.485 -175.955 ;
        RECT 271.155 -177.645 271.485 -177.315 ;
        RECT 271.155 -183.29 271.485 -182.16 ;
        RECT 271.16 -183.405 271.48 -95.04 ;
        RECT 271.155 -96.045 271.485 -95.715 ;
        RECT 271.155 -97.405 271.485 -97.075 ;
        RECT 271.155 -98.765 271.485 -98.435 ;
        RECT 271.155 -100.125 271.485 -99.795 ;
        RECT 271.155 -101.485 271.485 -101.155 ;
        RECT 271.155 -102.845 271.485 -102.515 ;
        RECT 271.155 -104.205 271.485 -103.875 ;
        RECT 271.155 -105.565 271.485 -105.235 ;
        RECT 271.155 -106.925 271.485 -106.595 ;
        RECT 271.155 -108.285 271.485 -107.955 ;
        RECT 271.155 -109.645 271.485 -109.315 ;
        RECT 271.155 -111.005 271.485 -110.675 ;
        RECT 271.155 -112.365 271.485 -112.035 ;
        RECT 271.155 -113.725 271.485 -113.395 ;
        RECT 271.155 -115.085 271.485 -114.755 ;
        RECT 271.155 -116.445 271.485 -116.115 ;
        RECT 271.155 -117.805 271.485 -117.475 ;
        RECT 271.155 -119.165 271.485 -118.835 ;
        RECT 271.155 -120.525 271.485 -120.195 ;
        RECT 271.155 -121.885 271.485 -121.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 203.96 -94.075 204.29 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 204.515 244.04 204.845 245.17 ;
        RECT 204.515 239.875 204.845 240.205 ;
        RECT 204.515 238.515 204.845 238.845 ;
        RECT 204.515 237.155 204.845 237.485 ;
        RECT 204.52 237.155 204.84 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 204.515 -96.045 204.845 -95.715 ;
        RECT 204.515 -97.405 204.845 -97.075 ;
        RECT 204.515 -98.765 204.845 -98.435 ;
        RECT 204.515 -100.125 204.845 -99.795 ;
        RECT 204.515 -101.485 204.845 -101.155 ;
        RECT 204.515 -102.845 204.845 -102.515 ;
        RECT 204.515 -104.205 204.845 -103.875 ;
        RECT 204.515 -105.565 204.845 -105.235 ;
        RECT 204.515 -106.925 204.845 -106.595 ;
        RECT 204.515 -108.285 204.845 -107.955 ;
        RECT 204.515 -109.645 204.845 -109.315 ;
        RECT 204.515 -111.005 204.845 -110.675 ;
        RECT 204.515 -112.365 204.845 -112.035 ;
        RECT 204.515 -113.725 204.845 -113.395 ;
        RECT 204.515 -115.085 204.845 -114.755 ;
        RECT 204.515 -116.445 204.845 -116.115 ;
        RECT 204.515 -117.805 204.845 -117.475 ;
        RECT 204.515 -119.165 204.845 -118.835 ;
        RECT 204.515 -120.525 204.845 -120.195 ;
        RECT 204.515 -121.885 204.845 -121.555 ;
        RECT 204.515 -123.245 204.845 -122.915 ;
        RECT 204.515 -124.605 204.845 -124.275 ;
        RECT 204.515 -125.965 204.845 -125.635 ;
        RECT 204.515 -127.325 204.845 -126.995 ;
        RECT 204.515 -128.685 204.845 -128.355 ;
        RECT 204.515 -130.045 204.845 -129.715 ;
        RECT 204.515 -131.405 204.845 -131.075 ;
        RECT 204.515 -132.765 204.845 -132.435 ;
        RECT 204.515 -134.125 204.845 -133.795 ;
        RECT 204.515 -135.485 204.845 -135.155 ;
        RECT 204.515 -136.845 204.845 -136.515 ;
        RECT 204.515 -138.205 204.845 -137.875 ;
        RECT 204.515 -139.565 204.845 -139.235 ;
        RECT 204.515 -140.925 204.845 -140.595 ;
        RECT 204.515 -142.285 204.845 -141.955 ;
        RECT 204.515 -143.645 204.845 -143.315 ;
        RECT 204.515 -145.005 204.845 -144.675 ;
        RECT 204.515 -146.365 204.845 -146.035 ;
        RECT 204.515 -147.725 204.845 -147.395 ;
        RECT 204.515 -149.085 204.845 -148.755 ;
        RECT 204.515 -150.445 204.845 -150.115 ;
        RECT 204.515 -151.805 204.845 -151.475 ;
        RECT 204.515 -153.165 204.845 -152.835 ;
        RECT 204.515 -154.525 204.845 -154.195 ;
        RECT 204.515 -155.885 204.845 -155.555 ;
        RECT 204.515 -157.245 204.845 -156.915 ;
        RECT 204.515 -158.605 204.845 -158.275 ;
        RECT 204.515 -159.965 204.845 -159.635 ;
        RECT 204.515 -161.325 204.845 -160.995 ;
        RECT 204.515 -162.685 204.845 -162.355 ;
        RECT 204.515 -164.045 204.845 -163.715 ;
        RECT 204.515 -165.405 204.845 -165.075 ;
        RECT 204.515 -166.765 204.845 -166.435 ;
        RECT 204.515 -168.125 204.845 -167.795 ;
        RECT 204.515 -169.485 204.845 -169.155 ;
        RECT 204.515 -170.845 204.845 -170.515 ;
        RECT 204.515 -172.205 204.845 -171.875 ;
        RECT 204.515 -173.565 204.845 -173.235 ;
        RECT 204.515 -174.925 204.845 -174.595 ;
        RECT 204.515 -176.285 204.845 -175.955 ;
        RECT 204.515 -177.645 204.845 -177.315 ;
        RECT 204.515 -183.29 204.845 -182.16 ;
        RECT 204.52 -183.405 204.84 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 205.875 244.04 206.205 245.17 ;
        RECT 205.875 239.875 206.205 240.205 ;
        RECT 205.875 238.515 206.205 238.845 ;
        RECT 205.875 237.155 206.205 237.485 ;
        RECT 205.88 237.155 206.2 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 205.875 -0.845 206.205 -0.515 ;
        RECT 205.875 -2.205 206.205 -1.875 ;
        RECT 205.875 -3.565 206.205 -3.235 ;
        RECT 205.88 -3.565 206.2 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 207.235 244.04 207.565 245.17 ;
        RECT 207.235 239.875 207.565 240.205 ;
        RECT 207.235 238.515 207.565 238.845 ;
        RECT 207.235 237.155 207.565 237.485 ;
        RECT 207.24 237.155 207.56 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 207.235 -0.845 207.565 -0.515 ;
        RECT 207.235 -2.205 207.565 -1.875 ;
        RECT 207.235 -3.565 207.565 -3.235 ;
        RECT 207.24 -3.565 207.56 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 208.595 244.04 208.925 245.17 ;
        RECT 208.595 239.875 208.925 240.205 ;
        RECT 208.595 238.515 208.925 238.845 ;
        RECT 208.595 237.155 208.925 237.485 ;
        RECT 208.6 237.155 208.92 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 208.595 -0.845 208.925 -0.515 ;
        RECT 208.595 -2.205 208.925 -1.875 ;
        RECT 208.595 -3.565 208.925 -3.235 ;
        RECT 208.6 -3.565 208.92 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 208.595 -91.965 208.925 -91.635 ;
        RECT 208.595 -93.325 208.925 -92.995 ;
        RECT 208.595 -94.685 208.925 -94.355 ;
        RECT 208.595 -96.045 208.925 -95.715 ;
        RECT 208.595 -97.405 208.925 -97.075 ;
        RECT 208.595 -98.765 208.925 -98.435 ;
        RECT 208.595 -100.125 208.925 -99.795 ;
        RECT 208.595 -101.485 208.925 -101.155 ;
        RECT 208.595 -102.845 208.925 -102.515 ;
        RECT 208.595 -104.205 208.925 -103.875 ;
        RECT 208.595 -105.565 208.925 -105.235 ;
        RECT 208.595 -106.925 208.925 -106.595 ;
        RECT 208.595 -108.285 208.925 -107.955 ;
        RECT 208.595 -109.645 208.925 -109.315 ;
        RECT 208.595 -111.005 208.925 -110.675 ;
        RECT 208.595 -112.365 208.925 -112.035 ;
        RECT 208.595 -113.725 208.925 -113.395 ;
        RECT 208.595 -115.085 208.925 -114.755 ;
        RECT 208.595 -116.445 208.925 -116.115 ;
        RECT 208.595 -117.805 208.925 -117.475 ;
        RECT 208.595 -119.165 208.925 -118.835 ;
        RECT 208.595 -120.525 208.925 -120.195 ;
        RECT 208.595 -121.885 208.925 -121.555 ;
        RECT 208.595 -123.245 208.925 -122.915 ;
        RECT 208.595 -124.605 208.925 -124.275 ;
        RECT 208.595 -125.965 208.925 -125.635 ;
        RECT 208.595 -127.325 208.925 -126.995 ;
        RECT 208.595 -128.685 208.925 -128.355 ;
        RECT 208.595 -130.045 208.925 -129.715 ;
        RECT 208.595 -131.405 208.925 -131.075 ;
        RECT 208.595 -132.765 208.925 -132.435 ;
        RECT 208.595 -134.125 208.925 -133.795 ;
        RECT 208.595 -135.485 208.925 -135.155 ;
        RECT 208.595 -136.845 208.925 -136.515 ;
        RECT 208.595 -138.205 208.925 -137.875 ;
        RECT 208.595 -139.565 208.925 -139.235 ;
        RECT 208.595 -140.925 208.925 -140.595 ;
        RECT 208.595 -142.285 208.925 -141.955 ;
        RECT 208.595 -143.645 208.925 -143.315 ;
        RECT 208.595 -145.005 208.925 -144.675 ;
        RECT 208.595 -146.365 208.925 -146.035 ;
        RECT 208.595 -147.725 208.925 -147.395 ;
        RECT 208.595 -149.085 208.925 -148.755 ;
        RECT 208.595 -150.445 208.925 -150.115 ;
        RECT 208.595 -151.805 208.925 -151.475 ;
        RECT 208.595 -153.165 208.925 -152.835 ;
        RECT 208.595 -154.525 208.925 -154.195 ;
        RECT 208.595 -155.885 208.925 -155.555 ;
        RECT 208.595 -157.245 208.925 -156.915 ;
        RECT 208.595 -158.605 208.925 -158.275 ;
        RECT 208.595 -159.965 208.925 -159.635 ;
        RECT 208.595 -161.325 208.925 -160.995 ;
        RECT 208.595 -162.685 208.925 -162.355 ;
        RECT 208.595 -164.045 208.925 -163.715 ;
        RECT 208.595 -165.405 208.925 -165.075 ;
        RECT 208.595 -166.765 208.925 -166.435 ;
        RECT 208.595 -168.125 208.925 -167.795 ;
        RECT 208.595 -169.485 208.925 -169.155 ;
        RECT 208.595 -170.845 208.925 -170.515 ;
        RECT 208.595 -172.205 208.925 -171.875 ;
        RECT 208.595 -173.565 208.925 -173.235 ;
        RECT 208.595 -174.925 208.925 -174.595 ;
        RECT 208.595 -176.285 208.925 -175.955 ;
        RECT 208.595 -177.645 208.925 -177.315 ;
        RECT 208.595 -183.29 208.925 -182.16 ;
        RECT 208.6 -183.405 208.92 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 209.955 244.04 210.285 245.17 ;
        RECT 209.955 239.875 210.285 240.205 ;
        RECT 209.955 238.515 210.285 238.845 ;
        RECT 209.955 237.155 210.285 237.485 ;
        RECT 209.96 237.155 210.28 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 209.955 -96.045 210.285 -95.715 ;
        RECT 209.955 -97.405 210.285 -97.075 ;
        RECT 209.955 -98.765 210.285 -98.435 ;
        RECT 209.955 -100.125 210.285 -99.795 ;
        RECT 209.955 -101.485 210.285 -101.155 ;
        RECT 209.955 -102.845 210.285 -102.515 ;
        RECT 209.955 -104.205 210.285 -103.875 ;
        RECT 209.955 -105.565 210.285 -105.235 ;
        RECT 209.955 -106.925 210.285 -106.595 ;
        RECT 209.955 -108.285 210.285 -107.955 ;
        RECT 209.955 -109.645 210.285 -109.315 ;
        RECT 209.955 -111.005 210.285 -110.675 ;
        RECT 209.955 -112.365 210.285 -112.035 ;
        RECT 209.955 -113.725 210.285 -113.395 ;
        RECT 209.955 -115.085 210.285 -114.755 ;
        RECT 209.955 -116.445 210.285 -116.115 ;
        RECT 209.955 -117.805 210.285 -117.475 ;
        RECT 209.955 -119.165 210.285 -118.835 ;
        RECT 209.955 -120.525 210.285 -120.195 ;
        RECT 209.955 -121.885 210.285 -121.555 ;
        RECT 209.955 -123.245 210.285 -122.915 ;
        RECT 209.955 -124.605 210.285 -124.275 ;
        RECT 209.955 -125.965 210.285 -125.635 ;
        RECT 209.955 -127.325 210.285 -126.995 ;
        RECT 209.955 -128.685 210.285 -128.355 ;
        RECT 209.955 -130.045 210.285 -129.715 ;
        RECT 209.955 -131.405 210.285 -131.075 ;
        RECT 209.955 -132.765 210.285 -132.435 ;
        RECT 209.955 -134.125 210.285 -133.795 ;
        RECT 209.955 -135.485 210.285 -135.155 ;
        RECT 209.955 -136.845 210.285 -136.515 ;
        RECT 209.955 -138.205 210.285 -137.875 ;
        RECT 209.955 -139.565 210.285 -139.235 ;
        RECT 209.955 -140.925 210.285 -140.595 ;
        RECT 209.955 -142.285 210.285 -141.955 ;
        RECT 209.955 -143.645 210.285 -143.315 ;
        RECT 209.955 -145.005 210.285 -144.675 ;
        RECT 209.955 -146.365 210.285 -146.035 ;
        RECT 209.955 -147.725 210.285 -147.395 ;
        RECT 209.955 -149.085 210.285 -148.755 ;
        RECT 209.955 -150.445 210.285 -150.115 ;
        RECT 209.955 -151.805 210.285 -151.475 ;
        RECT 209.955 -153.165 210.285 -152.835 ;
        RECT 209.955 -154.525 210.285 -154.195 ;
        RECT 209.955 -155.885 210.285 -155.555 ;
        RECT 209.955 -157.245 210.285 -156.915 ;
        RECT 209.955 -158.605 210.285 -158.275 ;
        RECT 209.955 -159.965 210.285 -159.635 ;
        RECT 209.955 -161.325 210.285 -160.995 ;
        RECT 209.955 -162.685 210.285 -162.355 ;
        RECT 209.955 -164.045 210.285 -163.715 ;
        RECT 209.955 -165.405 210.285 -165.075 ;
        RECT 209.955 -166.765 210.285 -166.435 ;
        RECT 209.955 -168.125 210.285 -167.795 ;
        RECT 209.955 -169.485 210.285 -169.155 ;
        RECT 209.955 -170.845 210.285 -170.515 ;
        RECT 209.955 -172.205 210.285 -171.875 ;
        RECT 209.955 -173.565 210.285 -173.235 ;
        RECT 209.955 -174.925 210.285 -174.595 ;
        RECT 209.955 -176.285 210.285 -175.955 ;
        RECT 209.955 -177.645 210.285 -177.315 ;
        RECT 209.955 -183.29 210.285 -182.16 ;
        RECT 209.96 -183.405 210.28 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 210.06 -94.075 210.39 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 211.315 244.04 211.645 245.17 ;
        RECT 211.315 239.875 211.645 240.205 ;
        RECT 211.315 238.515 211.645 238.845 ;
        RECT 211.315 237.155 211.645 237.485 ;
        RECT 211.32 237.155 211.64 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 212.675 244.04 213.005 245.17 ;
        RECT 212.675 239.875 213.005 240.205 ;
        RECT 212.675 238.515 213.005 238.845 ;
        RECT 212.675 237.155 213.005 237.485 ;
        RECT 212.68 237.155 213 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 212.675 -0.845 213.005 -0.515 ;
        RECT 212.675 -2.205 213.005 -1.875 ;
        RECT 212.675 -3.565 213.005 -3.235 ;
        RECT 212.68 -3.565 213 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 214.035 244.04 214.365 245.17 ;
        RECT 214.035 239.875 214.365 240.205 ;
        RECT 214.035 238.515 214.365 238.845 ;
        RECT 214.035 237.155 214.365 237.485 ;
        RECT 214.04 237.155 214.36 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 214.035 -0.845 214.365 -0.515 ;
        RECT 214.035 -2.205 214.365 -1.875 ;
        RECT 214.035 -3.565 214.365 -3.235 ;
        RECT 214.04 -3.565 214.36 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 214.035 -91.965 214.365 -91.635 ;
        RECT 214.035 -93.325 214.365 -92.995 ;
        RECT 214.035 -94.685 214.365 -94.355 ;
        RECT 214.035 -96.045 214.365 -95.715 ;
        RECT 214.035 -97.405 214.365 -97.075 ;
        RECT 214.035 -98.765 214.365 -98.435 ;
        RECT 214.035 -100.125 214.365 -99.795 ;
        RECT 214.035 -101.485 214.365 -101.155 ;
        RECT 214.035 -102.845 214.365 -102.515 ;
        RECT 214.035 -104.205 214.365 -103.875 ;
        RECT 214.035 -105.565 214.365 -105.235 ;
        RECT 214.035 -106.925 214.365 -106.595 ;
        RECT 214.035 -108.285 214.365 -107.955 ;
        RECT 214.035 -109.645 214.365 -109.315 ;
        RECT 214.035 -111.005 214.365 -110.675 ;
        RECT 214.035 -112.365 214.365 -112.035 ;
        RECT 214.035 -113.725 214.365 -113.395 ;
        RECT 214.035 -115.085 214.365 -114.755 ;
        RECT 214.035 -116.445 214.365 -116.115 ;
        RECT 214.035 -117.805 214.365 -117.475 ;
        RECT 214.035 -119.165 214.365 -118.835 ;
        RECT 214.035 -120.525 214.365 -120.195 ;
        RECT 214.035 -121.885 214.365 -121.555 ;
        RECT 214.035 -123.245 214.365 -122.915 ;
        RECT 214.035 -124.605 214.365 -124.275 ;
        RECT 214.035 -125.965 214.365 -125.635 ;
        RECT 214.035 -127.325 214.365 -126.995 ;
        RECT 214.035 -128.685 214.365 -128.355 ;
        RECT 214.035 -130.045 214.365 -129.715 ;
        RECT 214.035 -131.405 214.365 -131.075 ;
        RECT 214.035 -132.765 214.365 -132.435 ;
        RECT 214.035 -134.125 214.365 -133.795 ;
        RECT 214.035 -135.485 214.365 -135.155 ;
        RECT 214.035 -136.845 214.365 -136.515 ;
        RECT 214.035 -138.205 214.365 -137.875 ;
        RECT 214.035 -139.565 214.365 -139.235 ;
        RECT 214.035 -140.925 214.365 -140.595 ;
        RECT 214.035 -142.285 214.365 -141.955 ;
        RECT 214.035 -143.645 214.365 -143.315 ;
        RECT 214.035 -145.005 214.365 -144.675 ;
        RECT 214.035 -146.365 214.365 -146.035 ;
        RECT 214.035 -147.725 214.365 -147.395 ;
        RECT 214.035 -149.085 214.365 -148.755 ;
        RECT 214.035 -150.445 214.365 -150.115 ;
        RECT 214.035 -151.805 214.365 -151.475 ;
        RECT 214.035 -153.165 214.365 -152.835 ;
        RECT 214.035 -154.525 214.365 -154.195 ;
        RECT 214.035 -155.885 214.365 -155.555 ;
        RECT 214.035 -157.245 214.365 -156.915 ;
        RECT 214.035 -158.605 214.365 -158.275 ;
        RECT 214.035 -159.965 214.365 -159.635 ;
        RECT 214.035 -161.325 214.365 -160.995 ;
        RECT 214.035 -162.685 214.365 -162.355 ;
        RECT 214.035 -164.045 214.365 -163.715 ;
        RECT 214.035 -165.405 214.365 -165.075 ;
        RECT 214.035 -166.765 214.365 -166.435 ;
        RECT 214.035 -168.125 214.365 -167.795 ;
        RECT 214.035 -169.485 214.365 -169.155 ;
        RECT 214.035 -170.845 214.365 -170.515 ;
        RECT 214.035 -172.205 214.365 -171.875 ;
        RECT 214.035 -173.565 214.365 -173.235 ;
        RECT 214.035 -174.925 214.365 -174.595 ;
        RECT 214.035 -176.285 214.365 -175.955 ;
        RECT 214.035 -177.645 214.365 -177.315 ;
        RECT 214.035 -183.29 214.365 -182.16 ;
        RECT 214.04 -183.405 214.36 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 215.395 244.04 215.725 245.17 ;
        RECT 215.395 239.875 215.725 240.205 ;
        RECT 215.395 238.515 215.725 238.845 ;
        RECT 215.395 237.155 215.725 237.485 ;
        RECT 215.4 237.155 215.72 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 215.395 -0.845 215.725 -0.515 ;
        RECT 215.395 -2.205 215.725 -1.875 ;
        RECT 215.395 -3.565 215.725 -3.235 ;
        RECT 215.4 -3.565 215.72 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 215.395 -91.965 215.725 -91.635 ;
        RECT 215.395 -93.325 215.725 -92.995 ;
        RECT 215.395 -94.685 215.725 -94.355 ;
        RECT 215.395 -96.045 215.725 -95.715 ;
        RECT 215.395 -97.405 215.725 -97.075 ;
        RECT 215.395 -98.765 215.725 -98.435 ;
        RECT 215.395 -100.125 215.725 -99.795 ;
        RECT 215.395 -101.485 215.725 -101.155 ;
        RECT 215.395 -102.845 215.725 -102.515 ;
        RECT 215.395 -104.205 215.725 -103.875 ;
        RECT 215.395 -105.565 215.725 -105.235 ;
        RECT 215.395 -106.925 215.725 -106.595 ;
        RECT 215.395 -108.285 215.725 -107.955 ;
        RECT 215.395 -109.645 215.725 -109.315 ;
        RECT 215.395 -111.005 215.725 -110.675 ;
        RECT 215.395 -112.365 215.725 -112.035 ;
        RECT 215.395 -113.725 215.725 -113.395 ;
        RECT 215.395 -115.085 215.725 -114.755 ;
        RECT 215.395 -116.445 215.725 -116.115 ;
        RECT 215.395 -117.805 215.725 -117.475 ;
        RECT 215.395 -119.165 215.725 -118.835 ;
        RECT 215.395 -120.525 215.725 -120.195 ;
        RECT 215.395 -121.885 215.725 -121.555 ;
        RECT 215.395 -123.245 215.725 -122.915 ;
        RECT 215.395 -124.605 215.725 -124.275 ;
        RECT 215.395 -125.965 215.725 -125.635 ;
        RECT 215.395 -127.325 215.725 -126.995 ;
        RECT 215.395 -128.685 215.725 -128.355 ;
        RECT 215.395 -130.045 215.725 -129.715 ;
        RECT 215.395 -131.405 215.725 -131.075 ;
        RECT 215.395 -132.765 215.725 -132.435 ;
        RECT 215.395 -134.125 215.725 -133.795 ;
        RECT 215.395 -135.485 215.725 -135.155 ;
        RECT 215.395 -136.845 215.725 -136.515 ;
        RECT 215.395 -138.205 215.725 -137.875 ;
        RECT 215.395 -139.565 215.725 -139.235 ;
        RECT 215.395 -140.925 215.725 -140.595 ;
        RECT 215.395 -142.285 215.725 -141.955 ;
        RECT 215.395 -143.645 215.725 -143.315 ;
        RECT 215.395 -145.005 215.725 -144.675 ;
        RECT 215.395 -146.365 215.725 -146.035 ;
        RECT 215.395 -147.725 215.725 -147.395 ;
        RECT 215.395 -149.085 215.725 -148.755 ;
        RECT 215.395 -150.445 215.725 -150.115 ;
        RECT 215.395 -151.805 215.725 -151.475 ;
        RECT 215.395 -153.165 215.725 -152.835 ;
        RECT 215.395 -154.525 215.725 -154.195 ;
        RECT 215.395 -155.885 215.725 -155.555 ;
        RECT 215.395 -157.245 215.725 -156.915 ;
        RECT 215.395 -158.605 215.725 -158.275 ;
        RECT 215.395 -159.965 215.725 -159.635 ;
        RECT 215.395 -161.325 215.725 -160.995 ;
        RECT 215.395 -162.685 215.725 -162.355 ;
        RECT 215.395 -164.045 215.725 -163.715 ;
        RECT 215.395 -165.405 215.725 -165.075 ;
        RECT 215.395 -166.765 215.725 -166.435 ;
        RECT 215.395 -168.125 215.725 -167.795 ;
        RECT 215.395 -169.485 215.725 -169.155 ;
        RECT 215.395 -170.845 215.725 -170.515 ;
        RECT 215.395 -172.205 215.725 -171.875 ;
        RECT 215.395 -173.565 215.725 -173.235 ;
        RECT 215.395 -174.925 215.725 -174.595 ;
        RECT 215.395 -176.285 215.725 -175.955 ;
        RECT 215.395 -177.645 215.725 -177.315 ;
        RECT 215.395 -183.29 215.725 -182.16 ;
        RECT 215.4 -183.405 215.72 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 216.16 -94.075 216.49 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 216.755 244.04 217.085 245.17 ;
        RECT 216.755 239.875 217.085 240.205 ;
        RECT 216.755 238.515 217.085 238.845 ;
        RECT 216.755 237.155 217.085 237.485 ;
        RECT 216.76 237.155 217.08 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 216.755 -96.045 217.085 -95.715 ;
        RECT 216.755 -97.405 217.085 -97.075 ;
        RECT 216.755 -98.765 217.085 -98.435 ;
        RECT 216.755 -100.125 217.085 -99.795 ;
        RECT 216.755 -101.485 217.085 -101.155 ;
        RECT 216.755 -102.845 217.085 -102.515 ;
        RECT 216.755 -104.205 217.085 -103.875 ;
        RECT 216.755 -105.565 217.085 -105.235 ;
        RECT 216.755 -106.925 217.085 -106.595 ;
        RECT 216.755 -108.285 217.085 -107.955 ;
        RECT 216.755 -109.645 217.085 -109.315 ;
        RECT 216.755 -111.005 217.085 -110.675 ;
        RECT 216.755 -112.365 217.085 -112.035 ;
        RECT 216.755 -113.725 217.085 -113.395 ;
        RECT 216.755 -115.085 217.085 -114.755 ;
        RECT 216.755 -116.445 217.085 -116.115 ;
        RECT 216.755 -117.805 217.085 -117.475 ;
        RECT 216.755 -119.165 217.085 -118.835 ;
        RECT 216.755 -120.525 217.085 -120.195 ;
        RECT 216.755 -121.885 217.085 -121.555 ;
        RECT 216.755 -123.245 217.085 -122.915 ;
        RECT 216.755 -124.605 217.085 -124.275 ;
        RECT 216.755 -125.965 217.085 -125.635 ;
        RECT 216.755 -127.325 217.085 -126.995 ;
        RECT 216.755 -128.685 217.085 -128.355 ;
        RECT 216.755 -130.045 217.085 -129.715 ;
        RECT 216.755 -131.405 217.085 -131.075 ;
        RECT 216.755 -132.765 217.085 -132.435 ;
        RECT 216.755 -134.125 217.085 -133.795 ;
        RECT 216.755 -135.485 217.085 -135.155 ;
        RECT 216.755 -136.845 217.085 -136.515 ;
        RECT 216.755 -138.205 217.085 -137.875 ;
        RECT 216.755 -139.565 217.085 -139.235 ;
        RECT 216.755 -140.925 217.085 -140.595 ;
        RECT 216.755 -142.285 217.085 -141.955 ;
        RECT 216.755 -143.645 217.085 -143.315 ;
        RECT 216.755 -145.005 217.085 -144.675 ;
        RECT 216.755 -146.365 217.085 -146.035 ;
        RECT 216.755 -147.725 217.085 -147.395 ;
        RECT 216.755 -149.085 217.085 -148.755 ;
        RECT 216.755 -150.445 217.085 -150.115 ;
        RECT 216.755 -151.805 217.085 -151.475 ;
        RECT 216.755 -153.165 217.085 -152.835 ;
        RECT 216.755 -154.525 217.085 -154.195 ;
        RECT 216.755 -155.885 217.085 -155.555 ;
        RECT 216.755 -157.245 217.085 -156.915 ;
        RECT 216.755 -158.605 217.085 -158.275 ;
        RECT 216.755 -159.965 217.085 -159.635 ;
        RECT 216.755 -161.325 217.085 -160.995 ;
        RECT 216.755 -162.685 217.085 -162.355 ;
        RECT 216.755 -164.045 217.085 -163.715 ;
        RECT 216.755 -165.405 217.085 -165.075 ;
        RECT 216.755 -166.765 217.085 -166.435 ;
        RECT 216.755 -168.125 217.085 -167.795 ;
        RECT 216.755 -169.485 217.085 -169.155 ;
        RECT 216.755 -170.845 217.085 -170.515 ;
        RECT 216.755 -172.205 217.085 -171.875 ;
        RECT 216.755 -173.565 217.085 -173.235 ;
        RECT 216.755 -174.925 217.085 -174.595 ;
        RECT 216.755 -176.285 217.085 -175.955 ;
        RECT 216.755 -177.645 217.085 -177.315 ;
        RECT 216.755 -183.29 217.085 -182.16 ;
        RECT 216.76 -183.405 217.08 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 218.115 244.04 218.445 245.17 ;
        RECT 218.115 239.875 218.445 240.205 ;
        RECT 218.115 238.515 218.445 238.845 ;
        RECT 218.115 237.155 218.445 237.485 ;
        RECT 218.12 237.155 218.44 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 218.115 -0.845 218.445 -0.515 ;
        RECT 218.115 -2.205 218.445 -1.875 ;
        RECT 218.115 -3.565 218.445 -3.235 ;
        RECT 218.12 -3.565 218.44 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 219.475 244.04 219.805 245.17 ;
        RECT 219.475 239.875 219.805 240.205 ;
        RECT 219.475 238.515 219.805 238.845 ;
        RECT 219.475 237.155 219.805 237.485 ;
        RECT 219.48 237.155 219.8 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 219.475 -0.845 219.805 -0.515 ;
        RECT 219.475 -2.205 219.805 -1.875 ;
        RECT 219.475 -3.565 219.805 -3.235 ;
        RECT 219.48 -3.565 219.8 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 220.835 244.04 221.165 245.17 ;
        RECT 220.835 239.875 221.165 240.205 ;
        RECT 220.835 238.515 221.165 238.845 ;
        RECT 220.835 237.155 221.165 237.485 ;
        RECT 220.84 237.155 221.16 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 220.835 -0.845 221.165 -0.515 ;
        RECT 220.835 -2.205 221.165 -1.875 ;
        RECT 220.835 -3.565 221.165 -3.235 ;
        RECT 220.84 -3.565 221.16 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 220.835 -91.965 221.165 -91.635 ;
        RECT 220.835 -93.325 221.165 -92.995 ;
        RECT 220.835 -94.685 221.165 -94.355 ;
        RECT 220.835 -96.045 221.165 -95.715 ;
        RECT 220.835 -97.405 221.165 -97.075 ;
        RECT 220.835 -98.765 221.165 -98.435 ;
        RECT 220.835 -100.125 221.165 -99.795 ;
        RECT 220.835 -101.485 221.165 -101.155 ;
        RECT 220.835 -102.845 221.165 -102.515 ;
        RECT 220.835 -104.205 221.165 -103.875 ;
        RECT 220.835 -105.565 221.165 -105.235 ;
        RECT 220.835 -106.925 221.165 -106.595 ;
        RECT 220.835 -108.285 221.165 -107.955 ;
        RECT 220.835 -109.645 221.165 -109.315 ;
        RECT 220.835 -111.005 221.165 -110.675 ;
        RECT 220.835 -112.365 221.165 -112.035 ;
        RECT 220.835 -113.725 221.165 -113.395 ;
        RECT 220.835 -115.085 221.165 -114.755 ;
        RECT 220.835 -116.445 221.165 -116.115 ;
        RECT 220.835 -117.805 221.165 -117.475 ;
        RECT 220.835 -119.165 221.165 -118.835 ;
        RECT 220.835 -120.525 221.165 -120.195 ;
        RECT 220.835 -121.885 221.165 -121.555 ;
        RECT 220.835 -123.245 221.165 -122.915 ;
        RECT 220.835 -124.605 221.165 -124.275 ;
        RECT 220.835 -125.965 221.165 -125.635 ;
        RECT 220.835 -127.325 221.165 -126.995 ;
        RECT 220.835 -128.685 221.165 -128.355 ;
        RECT 220.835 -130.045 221.165 -129.715 ;
        RECT 220.835 -131.405 221.165 -131.075 ;
        RECT 220.835 -132.765 221.165 -132.435 ;
        RECT 220.835 -134.125 221.165 -133.795 ;
        RECT 220.835 -135.485 221.165 -135.155 ;
        RECT 220.835 -136.845 221.165 -136.515 ;
        RECT 220.835 -138.205 221.165 -137.875 ;
        RECT 220.835 -139.565 221.165 -139.235 ;
        RECT 220.835 -140.925 221.165 -140.595 ;
        RECT 220.835 -142.285 221.165 -141.955 ;
        RECT 220.835 -143.645 221.165 -143.315 ;
        RECT 220.835 -145.005 221.165 -144.675 ;
        RECT 220.835 -146.365 221.165 -146.035 ;
        RECT 220.835 -147.725 221.165 -147.395 ;
        RECT 220.835 -149.085 221.165 -148.755 ;
        RECT 220.835 -150.445 221.165 -150.115 ;
        RECT 220.835 -151.805 221.165 -151.475 ;
        RECT 220.835 -153.165 221.165 -152.835 ;
        RECT 220.835 -154.525 221.165 -154.195 ;
        RECT 220.835 -155.885 221.165 -155.555 ;
        RECT 220.835 -157.245 221.165 -156.915 ;
        RECT 220.835 -158.605 221.165 -158.275 ;
        RECT 220.835 -159.965 221.165 -159.635 ;
        RECT 220.835 -161.325 221.165 -160.995 ;
        RECT 220.835 -162.685 221.165 -162.355 ;
        RECT 220.835 -164.045 221.165 -163.715 ;
        RECT 220.835 -165.405 221.165 -165.075 ;
        RECT 220.835 -166.765 221.165 -166.435 ;
        RECT 220.835 -168.125 221.165 -167.795 ;
        RECT 220.835 -169.485 221.165 -169.155 ;
        RECT 220.835 -170.845 221.165 -170.515 ;
        RECT 220.835 -172.205 221.165 -171.875 ;
        RECT 220.835 -173.565 221.165 -173.235 ;
        RECT 220.835 -174.925 221.165 -174.595 ;
        RECT 220.835 -176.285 221.165 -175.955 ;
        RECT 220.835 -177.645 221.165 -177.315 ;
        RECT 220.835 -183.29 221.165 -182.16 ;
        RECT 220.84 -183.405 221.16 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 222.195 244.04 222.525 245.17 ;
        RECT 222.195 239.875 222.525 240.205 ;
        RECT 222.195 238.515 222.525 238.845 ;
        RECT 222.195 237.155 222.525 237.485 ;
        RECT 222.2 237.155 222.52 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 222.195 -96.045 222.525 -95.715 ;
        RECT 222.195 -97.405 222.525 -97.075 ;
        RECT 222.195 -98.765 222.525 -98.435 ;
        RECT 222.195 -100.125 222.525 -99.795 ;
        RECT 222.195 -101.485 222.525 -101.155 ;
        RECT 222.195 -102.845 222.525 -102.515 ;
        RECT 222.195 -104.205 222.525 -103.875 ;
        RECT 222.195 -105.565 222.525 -105.235 ;
        RECT 222.195 -106.925 222.525 -106.595 ;
        RECT 222.195 -108.285 222.525 -107.955 ;
        RECT 222.195 -109.645 222.525 -109.315 ;
        RECT 222.195 -111.005 222.525 -110.675 ;
        RECT 222.195 -112.365 222.525 -112.035 ;
        RECT 222.195 -113.725 222.525 -113.395 ;
        RECT 222.195 -115.085 222.525 -114.755 ;
        RECT 222.195 -116.445 222.525 -116.115 ;
        RECT 222.195 -117.805 222.525 -117.475 ;
        RECT 222.195 -119.165 222.525 -118.835 ;
        RECT 222.195 -120.525 222.525 -120.195 ;
        RECT 222.195 -121.885 222.525 -121.555 ;
        RECT 222.195 -123.245 222.525 -122.915 ;
        RECT 222.195 -124.605 222.525 -124.275 ;
        RECT 222.195 -125.965 222.525 -125.635 ;
        RECT 222.195 -127.325 222.525 -126.995 ;
        RECT 222.195 -128.685 222.525 -128.355 ;
        RECT 222.195 -130.045 222.525 -129.715 ;
        RECT 222.195 -131.405 222.525 -131.075 ;
        RECT 222.195 -132.765 222.525 -132.435 ;
        RECT 222.195 -134.125 222.525 -133.795 ;
        RECT 222.195 -135.485 222.525 -135.155 ;
        RECT 222.195 -136.845 222.525 -136.515 ;
        RECT 222.195 -138.205 222.525 -137.875 ;
        RECT 222.195 -139.565 222.525 -139.235 ;
        RECT 222.195 -140.925 222.525 -140.595 ;
        RECT 222.195 -142.285 222.525 -141.955 ;
        RECT 222.195 -143.645 222.525 -143.315 ;
        RECT 222.195 -145.005 222.525 -144.675 ;
        RECT 222.195 -146.365 222.525 -146.035 ;
        RECT 222.195 -147.725 222.525 -147.395 ;
        RECT 222.195 -149.085 222.525 -148.755 ;
        RECT 222.195 -150.445 222.525 -150.115 ;
        RECT 222.195 -151.805 222.525 -151.475 ;
        RECT 222.195 -153.165 222.525 -152.835 ;
        RECT 222.195 -154.525 222.525 -154.195 ;
        RECT 222.195 -155.885 222.525 -155.555 ;
        RECT 222.195 -157.245 222.525 -156.915 ;
        RECT 222.195 -158.605 222.525 -158.275 ;
        RECT 222.195 -159.965 222.525 -159.635 ;
        RECT 222.195 -161.325 222.525 -160.995 ;
        RECT 222.195 -162.685 222.525 -162.355 ;
        RECT 222.195 -164.045 222.525 -163.715 ;
        RECT 222.195 -165.405 222.525 -165.075 ;
        RECT 222.195 -166.765 222.525 -166.435 ;
        RECT 222.195 -168.125 222.525 -167.795 ;
        RECT 222.195 -169.485 222.525 -169.155 ;
        RECT 222.195 -170.845 222.525 -170.515 ;
        RECT 222.195 -172.205 222.525 -171.875 ;
        RECT 222.195 -173.565 222.525 -173.235 ;
        RECT 222.195 -174.925 222.525 -174.595 ;
        RECT 222.195 -176.285 222.525 -175.955 ;
        RECT 222.195 -177.645 222.525 -177.315 ;
        RECT 222.195 -183.29 222.525 -182.16 ;
        RECT 222.2 -183.405 222.52 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 222.26 -94.075 222.59 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 223.555 244.04 223.885 245.17 ;
        RECT 223.555 239.875 223.885 240.205 ;
        RECT 223.555 238.515 223.885 238.845 ;
        RECT 223.555 237.155 223.885 237.485 ;
        RECT 223.56 237.155 223.88 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 224.915 244.04 225.245 245.17 ;
        RECT 224.915 239.875 225.245 240.205 ;
        RECT 224.915 238.515 225.245 238.845 ;
        RECT 224.915 237.155 225.245 237.485 ;
        RECT 224.92 237.155 225.24 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 224.915 -0.845 225.245 -0.515 ;
        RECT 224.915 -2.205 225.245 -1.875 ;
        RECT 224.915 -3.565 225.245 -3.235 ;
        RECT 224.92 -3.565 225.24 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 226.275 244.04 226.605 245.17 ;
        RECT 226.275 239.875 226.605 240.205 ;
        RECT 226.275 238.515 226.605 238.845 ;
        RECT 226.275 237.155 226.605 237.485 ;
        RECT 226.28 237.155 226.6 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 226.275 -0.845 226.605 -0.515 ;
        RECT 226.275 -2.205 226.605 -1.875 ;
        RECT 226.275 -3.565 226.605 -3.235 ;
        RECT 226.28 -3.565 226.6 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 226.275 -91.965 226.605 -91.635 ;
        RECT 226.275 -93.325 226.605 -92.995 ;
        RECT 226.275 -94.685 226.605 -94.355 ;
        RECT 226.275 -96.045 226.605 -95.715 ;
        RECT 226.275 -97.405 226.605 -97.075 ;
        RECT 226.275 -98.765 226.605 -98.435 ;
        RECT 226.275 -100.125 226.605 -99.795 ;
        RECT 226.275 -101.485 226.605 -101.155 ;
        RECT 226.275 -102.845 226.605 -102.515 ;
        RECT 226.275 -104.205 226.605 -103.875 ;
        RECT 226.275 -105.565 226.605 -105.235 ;
        RECT 226.275 -106.925 226.605 -106.595 ;
        RECT 226.275 -108.285 226.605 -107.955 ;
        RECT 226.275 -109.645 226.605 -109.315 ;
        RECT 226.275 -111.005 226.605 -110.675 ;
        RECT 226.275 -112.365 226.605 -112.035 ;
        RECT 226.275 -113.725 226.605 -113.395 ;
        RECT 226.275 -115.085 226.605 -114.755 ;
        RECT 226.275 -116.445 226.605 -116.115 ;
        RECT 226.275 -117.805 226.605 -117.475 ;
        RECT 226.275 -119.165 226.605 -118.835 ;
        RECT 226.275 -120.525 226.605 -120.195 ;
        RECT 226.275 -121.885 226.605 -121.555 ;
        RECT 226.275 -123.245 226.605 -122.915 ;
        RECT 226.275 -124.605 226.605 -124.275 ;
        RECT 226.275 -125.965 226.605 -125.635 ;
        RECT 226.275 -127.325 226.605 -126.995 ;
        RECT 226.275 -128.685 226.605 -128.355 ;
        RECT 226.275 -130.045 226.605 -129.715 ;
        RECT 226.275 -131.405 226.605 -131.075 ;
        RECT 226.275 -132.765 226.605 -132.435 ;
        RECT 226.275 -134.125 226.605 -133.795 ;
        RECT 226.275 -135.485 226.605 -135.155 ;
        RECT 226.275 -136.845 226.605 -136.515 ;
        RECT 226.275 -138.205 226.605 -137.875 ;
        RECT 226.275 -139.565 226.605 -139.235 ;
        RECT 226.275 -140.925 226.605 -140.595 ;
        RECT 226.275 -142.285 226.605 -141.955 ;
        RECT 226.275 -143.645 226.605 -143.315 ;
        RECT 226.275 -145.005 226.605 -144.675 ;
        RECT 226.275 -146.365 226.605 -146.035 ;
        RECT 226.275 -147.725 226.605 -147.395 ;
        RECT 226.275 -149.085 226.605 -148.755 ;
        RECT 226.275 -150.445 226.605 -150.115 ;
        RECT 226.275 -151.805 226.605 -151.475 ;
        RECT 226.275 -153.165 226.605 -152.835 ;
        RECT 226.275 -154.525 226.605 -154.195 ;
        RECT 226.275 -155.885 226.605 -155.555 ;
        RECT 226.275 -157.245 226.605 -156.915 ;
        RECT 226.275 -158.605 226.605 -158.275 ;
        RECT 226.275 -159.965 226.605 -159.635 ;
        RECT 226.275 -161.325 226.605 -160.995 ;
        RECT 226.275 -162.685 226.605 -162.355 ;
        RECT 226.275 -164.045 226.605 -163.715 ;
        RECT 226.275 -165.405 226.605 -165.075 ;
        RECT 226.275 -166.765 226.605 -166.435 ;
        RECT 226.275 -168.125 226.605 -167.795 ;
        RECT 226.275 -169.485 226.605 -169.155 ;
        RECT 226.275 -170.845 226.605 -170.515 ;
        RECT 226.275 -172.205 226.605 -171.875 ;
        RECT 226.275 -173.565 226.605 -173.235 ;
        RECT 226.275 -174.925 226.605 -174.595 ;
        RECT 226.275 -176.285 226.605 -175.955 ;
        RECT 226.275 -177.645 226.605 -177.315 ;
        RECT 226.275 -183.29 226.605 -182.16 ;
        RECT 226.28 -183.405 226.6 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 227.635 244.04 227.965 245.17 ;
        RECT 227.635 239.875 227.965 240.205 ;
        RECT 227.635 238.515 227.965 238.845 ;
        RECT 227.635 237.155 227.965 237.485 ;
        RECT 227.64 237.155 227.96 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 227.635 -0.845 227.965 -0.515 ;
        RECT 227.635 -2.205 227.965 -1.875 ;
        RECT 227.635 -3.565 227.965 -3.235 ;
        RECT 227.64 -3.565 227.96 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 227.635 -91.965 227.965 -91.635 ;
        RECT 227.635 -93.325 227.965 -92.995 ;
        RECT 227.635 -94.685 227.965 -94.355 ;
        RECT 227.635 -96.045 227.965 -95.715 ;
        RECT 227.635 -97.405 227.965 -97.075 ;
        RECT 227.635 -98.765 227.965 -98.435 ;
        RECT 227.635 -100.125 227.965 -99.795 ;
        RECT 227.635 -101.485 227.965 -101.155 ;
        RECT 227.635 -102.845 227.965 -102.515 ;
        RECT 227.635 -104.205 227.965 -103.875 ;
        RECT 227.635 -105.565 227.965 -105.235 ;
        RECT 227.635 -106.925 227.965 -106.595 ;
        RECT 227.635 -108.285 227.965 -107.955 ;
        RECT 227.635 -109.645 227.965 -109.315 ;
        RECT 227.635 -111.005 227.965 -110.675 ;
        RECT 227.635 -112.365 227.965 -112.035 ;
        RECT 227.635 -113.725 227.965 -113.395 ;
        RECT 227.635 -115.085 227.965 -114.755 ;
        RECT 227.635 -116.445 227.965 -116.115 ;
        RECT 227.635 -117.805 227.965 -117.475 ;
        RECT 227.635 -119.165 227.965 -118.835 ;
        RECT 227.635 -120.525 227.965 -120.195 ;
        RECT 227.635 -121.885 227.965 -121.555 ;
        RECT 227.635 -123.245 227.965 -122.915 ;
        RECT 227.635 -124.605 227.965 -124.275 ;
        RECT 227.635 -125.965 227.965 -125.635 ;
        RECT 227.635 -127.325 227.965 -126.995 ;
        RECT 227.635 -128.685 227.965 -128.355 ;
        RECT 227.635 -130.045 227.965 -129.715 ;
        RECT 227.635 -131.405 227.965 -131.075 ;
        RECT 227.635 -132.765 227.965 -132.435 ;
        RECT 227.635 -134.125 227.965 -133.795 ;
        RECT 227.635 -135.485 227.965 -135.155 ;
        RECT 227.635 -136.845 227.965 -136.515 ;
        RECT 227.635 -138.205 227.965 -137.875 ;
        RECT 227.635 -139.565 227.965 -139.235 ;
        RECT 227.635 -140.925 227.965 -140.595 ;
        RECT 227.635 -142.285 227.965 -141.955 ;
        RECT 227.635 -143.645 227.965 -143.315 ;
        RECT 227.635 -145.005 227.965 -144.675 ;
        RECT 227.635 -146.365 227.965 -146.035 ;
        RECT 227.635 -147.725 227.965 -147.395 ;
        RECT 227.635 -149.085 227.965 -148.755 ;
        RECT 227.635 -150.445 227.965 -150.115 ;
        RECT 227.635 -151.805 227.965 -151.475 ;
        RECT 227.635 -153.165 227.965 -152.835 ;
        RECT 227.635 -154.525 227.965 -154.195 ;
        RECT 227.635 -155.885 227.965 -155.555 ;
        RECT 227.635 -157.245 227.965 -156.915 ;
        RECT 227.635 -158.605 227.965 -158.275 ;
        RECT 227.635 -159.965 227.965 -159.635 ;
        RECT 227.635 -161.325 227.965 -160.995 ;
        RECT 227.635 -162.685 227.965 -162.355 ;
        RECT 227.635 -164.045 227.965 -163.715 ;
        RECT 227.635 -165.405 227.965 -165.075 ;
        RECT 227.635 -166.765 227.965 -166.435 ;
        RECT 227.635 -168.125 227.965 -167.795 ;
        RECT 227.635 -169.485 227.965 -169.155 ;
        RECT 227.635 -170.845 227.965 -170.515 ;
        RECT 227.635 -172.205 227.965 -171.875 ;
        RECT 227.635 -173.565 227.965 -173.235 ;
        RECT 227.635 -174.925 227.965 -174.595 ;
        RECT 227.635 -176.285 227.965 -175.955 ;
        RECT 227.635 -177.645 227.965 -177.315 ;
        RECT 227.635 -183.29 227.965 -182.16 ;
        RECT 227.64 -183.405 227.96 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 228.36 -94.075 228.69 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 228.995 244.04 229.325 245.17 ;
        RECT 228.995 239.875 229.325 240.205 ;
        RECT 228.995 238.515 229.325 238.845 ;
        RECT 228.995 237.155 229.325 237.485 ;
        RECT 229 237.155 229.32 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 228.995 -96.045 229.325 -95.715 ;
        RECT 228.995 -97.405 229.325 -97.075 ;
        RECT 228.995 -98.765 229.325 -98.435 ;
        RECT 228.995 -100.125 229.325 -99.795 ;
        RECT 228.995 -101.485 229.325 -101.155 ;
        RECT 228.995 -102.845 229.325 -102.515 ;
        RECT 228.995 -104.205 229.325 -103.875 ;
        RECT 228.995 -105.565 229.325 -105.235 ;
        RECT 228.995 -106.925 229.325 -106.595 ;
        RECT 228.995 -108.285 229.325 -107.955 ;
        RECT 228.995 -109.645 229.325 -109.315 ;
        RECT 228.995 -111.005 229.325 -110.675 ;
        RECT 228.995 -112.365 229.325 -112.035 ;
        RECT 228.995 -113.725 229.325 -113.395 ;
        RECT 228.995 -115.085 229.325 -114.755 ;
        RECT 228.995 -116.445 229.325 -116.115 ;
        RECT 228.995 -117.805 229.325 -117.475 ;
        RECT 228.995 -119.165 229.325 -118.835 ;
        RECT 228.995 -120.525 229.325 -120.195 ;
        RECT 228.995 -121.885 229.325 -121.555 ;
        RECT 228.995 -123.245 229.325 -122.915 ;
        RECT 228.995 -124.605 229.325 -124.275 ;
        RECT 228.995 -125.965 229.325 -125.635 ;
        RECT 228.995 -127.325 229.325 -126.995 ;
        RECT 228.995 -128.685 229.325 -128.355 ;
        RECT 228.995 -130.045 229.325 -129.715 ;
        RECT 228.995 -131.405 229.325 -131.075 ;
        RECT 228.995 -132.765 229.325 -132.435 ;
        RECT 228.995 -134.125 229.325 -133.795 ;
        RECT 228.995 -135.485 229.325 -135.155 ;
        RECT 228.995 -136.845 229.325 -136.515 ;
        RECT 228.995 -138.205 229.325 -137.875 ;
        RECT 228.995 -139.565 229.325 -139.235 ;
        RECT 228.995 -140.925 229.325 -140.595 ;
        RECT 228.995 -142.285 229.325 -141.955 ;
        RECT 228.995 -143.645 229.325 -143.315 ;
        RECT 228.995 -145.005 229.325 -144.675 ;
        RECT 228.995 -146.365 229.325 -146.035 ;
        RECT 228.995 -147.725 229.325 -147.395 ;
        RECT 228.995 -149.085 229.325 -148.755 ;
        RECT 228.995 -150.445 229.325 -150.115 ;
        RECT 228.995 -151.805 229.325 -151.475 ;
        RECT 228.995 -153.165 229.325 -152.835 ;
        RECT 228.995 -154.525 229.325 -154.195 ;
        RECT 228.995 -155.885 229.325 -155.555 ;
        RECT 228.995 -157.245 229.325 -156.915 ;
        RECT 228.995 -158.605 229.325 -158.275 ;
        RECT 228.995 -159.965 229.325 -159.635 ;
        RECT 228.995 -161.325 229.325 -160.995 ;
        RECT 228.995 -162.685 229.325 -162.355 ;
        RECT 228.995 -164.045 229.325 -163.715 ;
        RECT 228.995 -165.405 229.325 -165.075 ;
        RECT 228.995 -166.765 229.325 -166.435 ;
        RECT 228.995 -168.125 229.325 -167.795 ;
        RECT 228.995 -169.485 229.325 -169.155 ;
        RECT 228.995 -170.845 229.325 -170.515 ;
        RECT 228.995 -172.205 229.325 -171.875 ;
        RECT 228.995 -173.565 229.325 -173.235 ;
        RECT 228.995 -174.925 229.325 -174.595 ;
        RECT 228.995 -176.285 229.325 -175.955 ;
        RECT 228.995 -177.645 229.325 -177.315 ;
        RECT 228.995 -183.29 229.325 -182.16 ;
        RECT 229 -183.405 229.32 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 230.355 244.04 230.685 245.17 ;
        RECT 230.355 239.875 230.685 240.205 ;
        RECT 230.355 238.515 230.685 238.845 ;
        RECT 230.355 237.155 230.685 237.485 ;
        RECT 230.36 237.155 230.68 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 230.355 -0.845 230.685 -0.515 ;
        RECT 230.355 -2.205 230.685 -1.875 ;
        RECT 230.355 -3.565 230.685 -3.235 ;
        RECT 230.36 -3.565 230.68 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 231.715 244.04 232.045 245.17 ;
        RECT 231.715 239.875 232.045 240.205 ;
        RECT 231.715 238.515 232.045 238.845 ;
        RECT 231.715 237.155 232.045 237.485 ;
        RECT 231.72 237.155 232.04 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 231.715 -0.845 232.045 -0.515 ;
        RECT 231.715 -2.205 232.045 -1.875 ;
        RECT 231.715 -3.565 232.045 -3.235 ;
        RECT 231.72 -3.565 232.04 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 233.075 244.04 233.405 245.17 ;
        RECT 233.075 239.875 233.405 240.205 ;
        RECT 233.075 238.515 233.405 238.845 ;
        RECT 233.075 237.155 233.405 237.485 ;
        RECT 233.08 237.155 233.4 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 233.075 -0.845 233.405 -0.515 ;
        RECT 233.075 -2.205 233.405 -1.875 ;
        RECT 233.075 -3.565 233.405 -3.235 ;
        RECT 233.08 -3.565 233.4 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 233.075 -91.965 233.405 -91.635 ;
        RECT 233.075 -93.325 233.405 -92.995 ;
        RECT 233.075 -94.685 233.405 -94.355 ;
        RECT 233.075 -96.045 233.405 -95.715 ;
        RECT 233.075 -97.405 233.405 -97.075 ;
        RECT 233.075 -98.765 233.405 -98.435 ;
        RECT 233.075 -100.125 233.405 -99.795 ;
        RECT 233.075 -101.485 233.405 -101.155 ;
        RECT 233.075 -102.845 233.405 -102.515 ;
        RECT 233.075 -104.205 233.405 -103.875 ;
        RECT 233.075 -105.565 233.405 -105.235 ;
        RECT 233.075 -106.925 233.405 -106.595 ;
        RECT 233.075 -108.285 233.405 -107.955 ;
        RECT 233.075 -109.645 233.405 -109.315 ;
        RECT 233.075 -111.005 233.405 -110.675 ;
        RECT 233.075 -112.365 233.405 -112.035 ;
        RECT 233.075 -113.725 233.405 -113.395 ;
        RECT 233.075 -115.085 233.405 -114.755 ;
        RECT 233.075 -116.445 233.405 -116.115 ;
        RECT 233.075 -117.805 233.405 -117.475 ;
        RECT 233.075 -119.165 233.405 -118.835 ;
        RECT 233.075 -120.525 233.405 -120.195 ;
        RECT 233.075 -121.885 233.405 -121.555 ;
        RECT 233.075 -123.245 233.405 -122.915 ;
        RECT 233.075 -124.605 233.405 -124.275 ;
        RECT 233.075 -125.965 233.405 -125.635 ;
        RECT 233.075 -127.325 233.405 -126.995 ;
        RECT 233.075 -128.685 233.405 -128.355 ;
        RECT 233.075 -130.045 233.405 -129.715 ;
        RECT 233.075 -131.405 233.405 -131.075 ;
        RECT 233.075 -132.765 233.405 -132.435 ;
        RECT 233.075 -134.125 233.405 -133.795 ;
        RECT 233.075 -135.485 233.405 -135.155 ;
        RECT 233.075 -136.845 233.405 -136.515 ;
        RECT 233.075 -138.205 233.405 -137.875 ;
        RECT 233.075 -139.565 233.405 -139.235 ;
        RECT 233.075 -140.925 233.405 -140.595 ;
        RECT 233.075 -142.285 233.405 -141.955 ;
        RECT 233.075 -143.645 233.405 -143.315 ;
        RECT 233.075 -145.005 233.405 -144.675 ;
        RECT 233.075 -146.365 233.405 -146.035 ;
        RECT 233.075 -147.725 233.405 -147.395 ;
        RECT 233.075 -149.085 233.405 -148.755 ;
        RECT 233.075 -150.445 233.405 -150.115 ;
        RECT 233.075 -151.805 233.405 -151.475 ;
        RECT 233.075 -153.165 233.405 -152.835 ;
        RECT 233.075 -154.525 233.405 -154.195 ;
        RECT 233.075 -155.885 233.405 -155.555 ;
        RECT 233.075 -157.245 233.405 -156.915 ;
        RECT 233.075 -158.605 233.405 -158.275 ;
        RECT 233.075 -159.965 233.405 -159.635 ;
        RECT 233.075 -161.325 233.405 -160.995 ;
        RECT 233.075 -162.685 233.405 -162.355 ;
        RECT 233.075 -164.045 233.405 -163.715 ;
        RECT 233.075 -165.405 233.405 -165.075 ;
        RECT 233.075 -166.765 233.405 -166.435 ;
        RECT 233.075 -168.125 233.405 -167.795 ;
        RECT 233.075 -169.485 233.405 -169.155 ;
        RECT 233.075 -170.845 233.405 -170.515 ;
        RECT 233.075 -172.205 233.405 -171.875 ;
        RECT 233.075 -173.565 233.405 -173.235 ;
        RECT 233.075 -174.925 233.405 -174.595 ;
        RECT 233.075 -176.285 233.405 -175.955 ;
        RECT 233.075 -177.645 233.405 -177.315 ;
        RECT 233.075 -183.29 233.405 -182.16 ;
        RECT 233.08 -183.405 233.4 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 234.435 244.04 234.765 245.17 ;
        RECT 234.435 239.875 234.765 240.205 ;
        RECT 234.435 238.515 234.765 238.845 ;
        RECT 234.435 237.155 234.765 237.485 ;
        RECT 234.44 237.155 234.76 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 234.435 -130.045 234.765 -129.715 ;
        RECT 234.435 -131.405 234.765 -131.075 ;
        RECT 234.435 -132.765 234.765 -132.435 ;
        RECT 234.435 -134.125 234.765 -133.795 ;
        RECT 234.435 -135.485 234.765 -135.155 ;
        RECT 234.435 -136.845 234.765 -136.515 ;
        RECT 234.435 -138.205 234.765 -137.875 ;
        RECT 234.435 -139.565 234.765 -139.235 ;
        RECT 234.435 -140.925 234.765 -140.595 ;
        RECT 234.435 -142.285 234.765 -141.955 ;
        RECT 234.435 -143.645 234.765 -143.315 ;
        RECT 234.435 -145.005 234.765 -144.675 ;
        RECT 234.435 -146.365 234.765 -146.035 ;
        RECT 234.435 -147.725 234.765 -147.395 ;
        RECT 234.435 -149.085 234.765 -148.755 ;
        RECT 234.435 -150.445 234.765 -150.115 ;
        RECT 234.435 -151.805 234.765 -151.475 ;
        RECT 234.435 -153.165 234.765 -152.835 ;
        RECT 234.435 -154.525 234.765 -154.195 ;
        RECT 234.435 -155.885 234.765 -155.555 ;
        RECT 234.435 -157.245 234.765 -156.915 ;
        RECT 234.435 -158.605 234.765 -158.275 ;
        RECT 234.435 -159.965 234.765 -159.635 ;
        RECT 234.435 -161.325 234.765 -160.995 ;
        RECT 234.435 -162.685 234.765 -162.355 ;
        RECT 234.435 -164.045 234.765 -163.715 ;
        RECT 234.435 -165.405 234.765 -165.075 ;
        RECT 234.435 -166.765 234.765 -166.435 ;
        RECT 234.435 -168.125 234.765 -167.795 ;
        RECT 234.435 -169.485 234.765 -169.155 ;
        RECT 234.435 -170.845 234.765 -170.515 ;
        RECT 234.435 -172.205 234.765 -171.875 ;
        RECT 234.435 -173.565 234.765 -173.235 ;
        RECT 234.435 -174.925 234.765 -174.595 ;
        RECT 234.435 -176.285 234.765 -175.955 ;
        RECT 234.435 -177.645 234.765 -177.315 ;
        RECT 234.435 -183.29 234.765 -182.16 ;
        RECT 234.44 -183.405 234.76 -95.04 ;
        RECT 234.435 -96.045 234.765 -95.715 ;
        RECT 234.435 -97.405 234.765 -97.075 ;
        RECT 234.435 -98.765 234.765 -98.435 ;
        RECT 234.435 -100.125 234.765 -99.795 ;
        RECT 234.435 -101.485 234.765 -101.155 ;
        RECT 234.435 -102.845 234.765 -102.515 ;
        RECT 234.435 -104.205 234.765 -103.875 ;
        RECT 234.435 -105.565 234.765 -105.235 ;
        RECT 234.435 -106.925 234.765 -106.595 ;
        RECT 234.435 -108.285 234.765 -107.955 ;
        RECT 234.435 -109.645 234.765 -109.315 ;
        RECT 234.435 -111.005 234.765 -110.675 ;
        RECT 234.435 -112.365 234.765 -112.035 ;
        RECT 234.435 -113.725 234.765 -113.395 ;
        RECT 234.435 -115.085 234.765 -114.755 ;
        RECT 234.435 -116.445 234.765 -116.115 ;
        RECT 234.435 -117.805 234.765 -117.475 ;
        RECT 234.435 -119.165 234.765 -118.835 ;
        RECT 234.435 -120.525 234.765 -120.195 ;
        RECT 234.435 -121.885 234.765 -121.555 ;
        RECT 234.435 -123.245 234.765 -122.915 ;
        RECT 234.435 -124.605 234.765 -124.275 ;
        RECT 234.435 -125.965 234.765 -125.635 ;
        RECT 234.435 -127.325 234.765 -126.995 ;
        RECT 234.435 -128.685 234.765 -128.355 ;
    END
    PORT
      LAYER met3 ;
        RECT 173.235 244.04 173.565 245.17 ;
        RECT 173.235 239.875 173.565 240.205 ;
        RECT 173.235 238.515 173.565 238.845 ;
        RECT 173.235 237.155 173.565 237.485 ;
        RECT 173.24 237.155 173.56 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 173.235 -96.045 173.565 -95.715 ;
        RECT 173.235 -97.405 173.565 -97.075 ;
        RECT 173.235 -98.765 173.565 -98.435 ;
        RECT 173.235 -100.125 173.565 -99.795 ;
        RECT 173.235 -101.485 173.565 -101.155 ;
        RECT 173.235 -102.845 173.565 -102.515 ;
        RECT 173.235 -104.205 173.565 -103.875 ;
        RECT 173.235 -105.565 173.565 -105.235 ;
        RECT 173.235 -106.925 173.565 -106.595 ;
        RECT 173.235 -108.285 173.565 -107.955 ;
        RECT 173.235 -109.645 173.565 -109.315 ;
        RECT 173.235 -111.005 173.565 -110.675 ;
        RECT 173.235 -112.365 173.565 -112.035 ;
        RECT 173.235 -113.725 173.565 -113.395 ;
        RECT 173.235 -115.085 173.565 -114.755 ;
        RECT 173.235 -116.445 173.565 -116.115 ;
        RECT 173.235 -117.805 173.565 -117.475 ;
        RECT 173.235 -119.165 173.565 -118.835 ;
        RECT 173.235 -120.525 173.565 -120.195 ;
        RECT 173.235 -121.885 173.565 -121.555 ;
        RECT 173.235 -123.245 173.565 -122.915 ;
        RECT 173.235 -124.605 173.565 -124.275 ;
        RECT 173.235 -125.965 173.565 -125.635 ;
        RECT 173.235 -127.325 173.565 -126.995 ;
        RECT 173.235 -128.685 173.565 -128.355 ;
        RECT 173.235 -130.045 173.565 -129.715 ;
        RECT 173.235 -131.405 173.565 -131.075 ;
        RECT 173.235 -132.765 173.565 -132.435 ;
        RECT 173.235 -134.125 173.565 -133.795 ;
        RECT 173.235 -135.485 173.565 -135.155 ;
        RECT 173.235 -136.845 173.565 -136.515 ;
        RECT 173.235 -138.205 173.565 -137.875 ;
        RECT 173.235 -139.565 173.565 -139.235 ;
        RECT 173.235 -140.925 173.565 -140.595 ;
        RECT 173.235 -142.285 173.565 -141.955 ;
        RECT 173.235 -143.645 173.565 -143.315 ;
        RECT 173.235 -145.005 173.565 -144.675 ;
        RECT 173.235 -146.365 173.565 -146.035 ;
        RECT 173.235 -147.725 173.565 -147.395 ;
        RECT 173.235 -149.085 173.565 -148.755 ;
        RECT 173.235 -150.445 173.565 -150.115 ;
        RECT 173.235 -151.805 173.565 -151.475 ;
        RECT 173.235 -153.165 173.565 -152.835 ;
        RECT 173.235 -154.525 173.565 -154.195 ;
        RECT 173.235 -155.885 173.565 -155.555 ;
        RECT 173.235 -157.245 173.565 -156.915 ;
        RECT 173.235 -158.605 173.565 -158.275 ;
        RECT 173.235 -159.965 173.565 -159.635 ;
        RECT 173.235 -161.325 173.565 -160.995 ;
        RECT 173.235 -162.685 173.565 -162.355 ;
        RECT 173.235 -164.045 173.565 -163.715 ;
        RECT 173.235 -165.405 173.565 -165.075 ;
        RECT 173.235 -166.765 173.565 -166.435 ;
        RECT 173.235 -168.125 173.565 -167.795 ;
        RECT 173.235 -169.485 173.565 -169.155 ;
        RECT 173.235 -170.845 173.565 -170.515 ;
        RECT 173.235 -172.205 173.565 -171.875 ;
        RECT 173.235 -173.565 173.565 -173.235 ;
        RECT 173.235 -174.925 173.565 -174.595 ;
        RECT 173.235 -176.285 173.565 -175.955 ;
        RECT 173.235 -177.645 173.565 -177.315 ;
        RECT 173.235 -183.29 173.565 -182.16 ;
        RECT 173.24 -183.405 173.56 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 173.46 -94.075 173.79 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 174.595 244.04 174.925 245.17 ;
        RECT 174.595 239.875 174.925 240.205 ;
        RECT 174.595 238.515 174.925 238.845 ;
        RECT 174.595 237.155 174.925 237.485 ;
        RECT 174.6 237.155 174.92 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 175.955 244.04 176.285 245.17 ;
        RECT 175.955 239.875 176.285 240.205 ;
        RECT 175.955 238.515 176.285 238.845 ;
        RECT 175.955 237.155 176.285 237.485 ;
        RECT 175.96 237.155 176.28 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 175.955 -0.845 176.285 -0.515 ;
        RECT 175.955 -2.205 176.285 -1.875 ;
        RECT 175.955 -3.565 176.285 -3.235 ;
        RECT 175.96 -3.565 176.28 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 177.315 244.04 177.645 245.17 ;
        RECT 177.315 239.875 177.645 240.205 ;
        RECT 177.315 238.515 177.645 238.845 ;
        RECT 177.315 237.155 177.645 237.485 ;
        RECT 177.32 237.155 177.64 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 177.315 -0.845 177.645 -0.515 ;
        RECT 177.315 -2.205 177.645 -1.875 ;
        RECT 177.315 -3.565 177.645 -3.235 ;
        RECT 177.32 -3.565 177.64 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 177.315 -91.965 177.645 -91.635 ;
        RECT 177.315 -93.325 177.645 -92.995 ;
        RECT 177.315 -94.685 177.645 -94.355 ;
        RECT 177.315 -96.045 177.645 -95.715 ;
        RECT 177.315 -97.405 177.645 -97.075 ;
        RECT 177.315 -98.765 177.645 -98.435 ;
        RECT 177.315 -100.125 177.645 -99.795 ;
        RECT 177.315 -101.485 177.645 -101.155 ;
        RECT 177.315 -102.845 177.645 -102.515 ;
        RECT 177.315 -104.205 177.645 -103.875 ;
        RECT 177.315 -105.565 177.645 -105.235 ;
        RECT 177.315 -106.925 177.645 -106.595 ;
        RECT 177.315 -108.285 177.645 -107.955 ;
        RECT 177.315 -109.645 177.645 -109.315 ;
        RECT 177.315 -111.005 177.645 -110.675 ;
        RECT 177.315 -112.365 177.645 -112.035 ;
        RECT 177.315 -113.725 177.645 -113.395 ;
        RECT 177.315 -115.085 177.645 -114.755 ;
        RECT 177.315 -116.445 177.645 -116.115 ;
        RECT 177.315 -117.805 177.645 -117.475 ;
        RECT 177.315 -119.165 177.645 -118.835 ;
        RECT 177.315 -120.525 177.645 -120.195 ;
        RECT 177.315 -121.885 177.645 -121.555 ;
        RECT 177.315 -123.245 177.645 -122.915 ;
        RECT 177.315 -124.605 177.645 -124.275 ;
        RECT 177.315 -125.965 177.645 -125.635 ;
        RECT 177.315 -127.325 177.645 -126.995 ;
        RECT 177.315 -128.685 177.645 -128.355 ;
        RECT 177.315 -130.045 177.645 -129.715 ;
        RECT 177.315 -131.405 177.645 -131.075 ;
        RECT 177.315 -132.765 177.645 -132.435 ;
        RECT 177.315 -134.125 177.645 -133.795 ;
        RECT 177.315 -135.485 177.645 -135.155 ;
        RECT 177.315 -136.845 177.645 -136.515 ;
        RECT 177.315 -138.205 177.645 -137.875 ;
        RECT 177.315 -139.565 177.645 -139.235 ;
        RECT 177.315 -140.925 177.645 -140.595 ;
        RECT 177.315 -142.285 177.645 -141.955 ;
        RECT 177.315 -143.645 177.645 -143.315 ;
        RECT 177.315 -145.005 177.645 -144.675 ;
        RECT 177.315 -146.365 177.645 -146.035 ;
        RECT 177.315 -147.725 177.645 -147.395 ;
        RECT 177.315 -149.085 177.645 -148.755 ;
        RECT 177.315 -150.445 177.645 -150.115 ;
        RECT 177.315 -151.805 177.645 -151.475 ;
        RECT 177.315 -153.165 177.645 -152.835 ;
        RECT 177.315 -154.525 177.645 -154.195 ;
        RECT 177.315 -155.885 177.645 -155.555 ;
        RECT 177.315 -157.245 177.645 -156.915 ;
        RECT 177.315 -158.605 177.645 -158.275 ;
        RECT 177.315 -159.965 177.645 -159.635 ;
        RECT 177.315 -161.325 177.645 -160.995 ;
        RECT 177.315 -162.685 177.645 -162.355 ;
        RECT 177.315 -164.045 177.645 -163.715 ;
        RECT 177.315 -165.405 177.645 -165.075 ;
        RECT 177.315 -166.765 177.645 -166.435 ;
        RECT 177.315 -168.125 177.645 -167.795 ;
        RECT 177.315 -169.485 177.645 -169.155 ;
        RECT 177.315 -170.845 177.645 -170.515 ;
        RECT 177.315 -172.205 177.645 -171.875 ;
        RECT 177.315 -173.565 177.645 -173.235 ;
        RECT 177.315 -174.925 177.645 -174.595 ;
        RECT 177.315 -176.285 177.645 -175.955 ;
        RECT 177.315 -177.645 177.645 -177.315 ;
        RECT 177.315 -183.29 177.645 -182.16 ;
        RECT 177.32 -183.405 177.64 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 178.675 244.04 179.005 245.17 ;
        RECT 178.675 239.875 179.005 240.205 ;
        RECT 178.675 238.515 179.005 238.845 ;
        RECT 178.675 237.155 179.005 237.485 ;
        RECT 178.68 237.155 179 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 178.675 -0.845 179.005 -0.515 ;
        RECT 178.675 -2.205 179.005 -1.875 ;
        RECT 178.675 -3.565 179.005 -3.235 ;
        RECT 178.68 -3.565 179 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 178.675 -91.965 179.005 -91.635 ;
        RECT 178.675 -93.325 179.005 -92.995 ;
        RECT 178.675 -94.685 179.005 -94.355 ;
        RECT 178.675 -96.045 179.005 -95.715 ;
        RECT 178.675 -97.405 179.005 -97.075 ;
        RECT 178.675 -98.765 179.005 -98.435 ;
        RECT 178.675 -100.125 179.005 -99.795 ;
        RECT 178.675 -101.485 179.005 -101.155 ;
        RECT 178.675 -102.845 179.005 -102.515 ;
        RECT 178.675 -104.205 179.005 -103.875 ;
        RECT 178.675 -105.565 179.005 -105.235 ;
        RECT 178.675 -106.925 179.005 -106.595 ;
        RECT 178.675 -108.285 179.005 -107.955 ;
        RECT 178.675 -109.645 179.005 -109.315 ;
        RECT 178.675 -111.005 179.005 -110.675 ;
        RECT 178.675 -112.365 179.005 -112.035 ;
        RECT 178.675 -113.725 179.005 -113.395 ;
        RECT 178.675 -115.085 179.005 -114.755 ;
        RECT 178.675 -116.445 179.005 -116.115 ;
        RECT 178.675 -117.805 179.005 -117.475 ;
        RECT 178.675 -119.165 179.005 -118.835 ;
        RECT 178.675 -120.525 179.005 -120.195 ;
        RECT 178.675 -121.885 179.005 -121.555 ;
        RECT 178.675 -123.245 179.005 -122.915 ;
        RECT 178.675 -124.605 179.005 -124.275 ;
        RECT 178.675 -125.965 179.005 -125.635 ;
        RECT 178.675 -127.325 179.005 -126.995 ;
        RECT 178.675 -128.685 179.005 -128.355 ;
        RECT 178.675 -130.045 179.005 -129.715 ;
        RECT 178.675 -131.405 179.005 -131.075 ;
        RECT 178.675 -132.765 179.005 -132.435 ;
        RECT 178.675 -134.125 179.005 -133.795 ;
        RECT 178.675 -135.485 179.005 -135.155 ;
        RECT 178.675 -136.845 179.005 -136.515 ;
        RECT 178.675 -138.205 179.005 -137.875 ;
        RECT 178.675 -139.565 179.005 -139.235 ;
        RECT 178.675 -140.925 179.005 -140.595 ;
        RECT 178.675 -142.285 179.005 -141.955 ;
        RECT 178.675 -143.645 179.005 -143.315 ;
        RECT 178.675 -145.005 179.005 -144.675 ;
        RECT 178.675 -146.365 179.005 -146.035 ;
        RECT 178.675 -147.725 179.005 -147.395 ;
        RECT 178.675 -149.085 179.005 -148.755 ;
        RECT 178.675 -150.445 179.005 -150.115 ;
        RECT 178.675 -151.805 179.005 -151.475 ;
        RECT 178.675 -153.165 179.005 -152.835 ;
        RECT 178.675 -154.525 179.005 -154.195 ;
        RECT 178.675 -155.885 179.005 -155.555 ;
        RECT 178.675 -157.245 179.005 -156.915 ;
        RECT 178.675 -158.605 179.005 -158.275 ;
        RECT 178.675 -159.965 179.005 -159.635 ;
        RECT 178.675 -161.325 179.005 -160.995 ;
        RECT 178.675 -162.685 179.005 -162.355 ;
        RECT 178.675 -164.045 179.005 -163.715 ;
        RECT 178.675 -165.405 179.005 -165.075 ;
        RECT 178.675 -166.765 179.005 -166.435 ;
        RECT 178.675 -168.125 179.005 -167.795 ;
        RECT 178.675 -169.485 179.005 -169.155 ;
        RECT 178.675 -170.845 179.005 -170.515 ;
        RECT 178.675 -172.205 179.005 -171.875 ;
        RECT 178.675 -173.565 179.005 -173.235 ;
        RECT 178.675 -174.925 179.005 -174.595 ;
        RECT 178.675 -176.285 179.005 -175.955 ;
        RECT 178.675 -177.645 179.005 -177.315 ;
        RECT 178.675 -183.29 179.005 -182.16 ;
        RECT 178.68 -183.405 179 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 179.56 -94.075 179.89 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 180.035 244.04 180.365 245.17 ;
        RECT 180.035 239.875 180.365 240.205 ;
        RECT 180.035 238.515 180.365 238.845 ;
        RECT 180.035 237.155 180.365 237.485 ;
        RECT 180.04 237.155 180.36 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 180.035 -96.045 180.365 -95.715 ;
        RECT 180.035 -97.405 180.365 -97.075 ;
        RECT 180.035 -98.765 180.365 -98.435 ;
        RECT 180.035 -100.125 180.365 -99.795 ;
        RECT 180.035 -101.485 180.365 -101.155 ;
        RECT 180.035 -102.845 180.365 -102.515 ;
        RECT 180.035 -104.205 180.365 -103.875 ;
        RECT 180.035 -105.565 180.365 -105.235 ;
        RECT 180.035 -106.925 180.365 -106.595 ;
        RECT 180.035 -108.285 180.365 -107.955 ;
        RECT 180.035 -109.645 180.365 -109.315 ;
        RECT 180.035 -111.005 180.365 -110.675 ;
        RECT 180.035 -112.365 180.365 -112.035 ;
        RECT 180.035 -113.725 180.365 -113.395 ;
        RECT 180.035 -115.085 180.365 -114.755 ;
        RECT 180.035 -116.445 180.365 -116.115 ;
        RECT 180.035 -117.805 180.365 -117.475 ;
        RECT 180.035 -119.165 180.365 -118.835 ;
        RECT 180.035 -120.525 180.365 -120.195 ;
        RECT 180.035 -121.885 180.365 -121.555 ;
        RECT 180.035 -123.245 180.365 -122.915 ;
        RECT 180.035 -124.605 180.365 -124.275 ;
        RECT 180.035 -125.965 180.365 -125.635 ;
        RECT 180.035 -127.325 180.365 -126.995 ;
        RECT 180.035 -128.685 180.365 -128.355 ;
        RECT 180.035 -130.045 180.365 -129.715 ;
        RECT 180.035 -131.405 180.365 -131.075 ;
        RECT 180.035 -132.765 180.365 -132.435 ;
        RECT 180.035 -134.125 180.365 -133.795 ;
        RECT 180.035 -135.485 180.365 -135.155 ;
        RECT 180.035 -136.845 180.365 -136.515 ;
        RECT 180.035 -138.205 180.365 -137.875 ;
        RECT 180.035 -139.565 180.365 -139.235 ;
        RECT 180.035 -140.925 180.365 -140.595 ;
        RECT 180.035 -142.285 180.365 -141.955 ;
        RECT 180.035 -143.645 180.365 -143.315 ;
        RECT 180.035 -145.005 180.365 -144.675 ;
        RECT 180.035 -146.365 180.365 -146.035 ;
        RECT 180.035 -147.725 180.365 -147.395 ;
        RECT 180.035 -149.085 180.365 -148.755 ;
        RECT 180.035 -150.445 180.365 -150.115 ;
        RECT 180.035 -151.805 180.365 -151.475 ;
        RECT 180.035 -153.165 180.365 -152.835 ;
        RECT 180.035 -154.525 180.365 -154.195 ;
        RECT 180.035 -155.885 180.365 -155.555 ;
        RECT 180.035 -157.245 180.365 -156.915 ;
        RECT 180.035 -158.605 180.365 -158.275 ;
        RECT 180.035 -159.965 180.365 -159.635 ;
        RECT 180.035 -161.325 180.365 -160.995 ;
        RECT 180.035 -162.685 180.365 -162.355 ;
        RECT 180.035 -164.045 180.365 -163.715 ;
        RECT 180.035 -165.405 180.365 -165.075 ;
        RECT 180.035 -166.765 180.365 -166.435 ;
        RECT 180.035 -168.125 180.365 -167.795 ;
        RECT 180.035 -169.485 180.365 -169.155 ;
        RECT 180.035 -170.845 180.365 -170.515 ;
        RECT 180.035 -172.205 180.365 -171.875 ;
        RECT 180.035 -173.565 180.365 -173.235 ;
        RECT 180.035 -174.925 180.365 -174.595 ;
        RECT 180.035 -176.285 180.365 -175.955 ;
        RECT 180.035 -177.645 180.365 -177.315 ;
        RECT 180.035 -183.29 180.365 -182.16 ;
        RECT 180.04 -183.405 180.36 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 181.395 244.04 181.725 245.17 ;
        RECT 181.395 239.875 181.725 240.205 ;
        RECT 181.395 238.515 181.725 238.845 ;
        RECT 181.395 237.155 181.725 237.485 ;
        RECT 181.4 237.155 181.72 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 181.395 -0.845 181.725 -0.515 ;
        RECT 181.395 -2.205 181.725 -1.875 ;
        RECT 181.395 -3.565 181.725 -3.235 ;
        RECT 181.4 -3.565 181.72 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 182.755 244.04 183.085 245.17 ;
        RECT 182.755 239.875 183.085 240.205 ;
        RECT 182.755 238.515 183.085 238.845 ;
        RECT 182.755 237.155 183.085 237.485 ;
        RECT 182.76 237.155 183.08 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 182.755 -0.845 183.085 -0.515 ;
        RECT 182.755 -2.205 183.085 -1.875 ;
        RECT 182.755 -3.565 183.085 -3.235 ;
        RECT 182.76 -3.565 183.08 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 184.115 244.04 184.445 245.17 ;
        RECT 184.115 239.875 184.445 240.205 ;
        RECT 184.115 238.515 184.445 238.845 ;
        RECT 184.115 237.155 184.445 237.485 ;
        RECT 184.12 237.155 184.44 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 184.115 -0.845 184.445 -0.515 ;
        RECT 184.115 -2.205 184.445 -1.875 ;
        RECT 184.115 -3.565 184.445 -3.235 ;
        RECT 184.12 -3.565 184.44 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 184.115 -91.965 184.445 -91.635 ;
        RECT 184.115 -93.325 184.445 -92.995 ;
        RECT 184.115 -94.685 184.445 -94.355 ;
        RECT 184.115 -96.045 184.445 -95.715 ;
        RECT 184.115 -97.405 184.445 -97.075 ;
        RECT 184.115 -98.765 184.445 -98.435 ;
        RECT 184.115 -100.125 184.445 -99.795 ;
        RECT 184.115 -101.485 184.445 -101.155 ;
        RECT 184.115 -102.845 184.445 -102.515 ;
        RECT 184.115 -104.205 184.445 -103.875 ;
        RECT 184.115 -105.565 184.445 -105.235 ;
        RECT 184.115 -106.925 184.445 -106.595 ;
        RECT 184.115 -108.285 184.445 -107.955 ;
        RECT 184.115 -109.645 184.445 -109.315 ;
        RECT 184.115 -111.005 184.445 -110.675 ;
        RECT 184.115 -112.365 184.445 -112.035 ;
        RECT 184.115 -113.725 184.445 -113.395 ;
        RECT 184.115 -115.085 184.445 -114.755 ;
        RECT 184.115 -116.445 184.445 -116.115 ;
        RECT 184.115 -117.805 184.445 -117.475 ;
        RECT 184.115 -119.165 184.445 -118.835 ;
        RECT 184.115 -120.525 184.445 -120.195 ;
        RECT 184.115 -121.885 184.445 -121.555 ;
        RECT 184.115 -123.245 184.445 -122.915 ;
        RECT 184.115 -124.605 184.445 -124.275 ;
        RECT 184.115 -125.965 184.445 -125.635 ;
        RECT 184.115 -127.325 184.445 -126.995 ;
        RECT 184.115 -128.685 184.445 -128.355 ;
        RECT 184.115 -130.045 184.445 -129.715 ;
        RECT 184.115 -131.405 184.445 -131.075 ;
        RECT 184.115 -132.765 184.445 -132.435 ;
        RECT 184.115 -134.125 184.445 -133.795 ;
        RECT 184.115 -135.485 184.445 -135.155 ;
        RECT 184.115 -136.845 184.445 -136.515 ;
        RECT 184.115 -138.205 184.445 -137.875 ;
        RECT 184.115 -139.565 184.445 -139.235 ;
        RECT 184.115 -140.925 184.445 -140.595 ;
        RECT 184.115 -142.285 184.445 -141.955 ;
        RECT 184.115 -143.645 184.445 -143.315 ;
        RECT 184.115 -145.005 184.445 -144.675 ;
        RECT 184.115 -146.365 184.445 -146.035 ;
        RECT 184.115 -147.725 184.445 -147.395 ;
        RECT 184.115 -149.085 184.445 -148.755 ;
        RECT 184.115 -150.445 184.445 -150.115 ;
        RECT 184.115 -151.805 184.445 -151.475 ;
        RECT 184.115 -153.165 184.445 -152.835 ;
        RECT 184.115 -154.525 184.445 -154.195 ;
        RECT 184.115 -155.885 184.445 -155.555 ;
        RECT 184.115 -157.245 184.445 -156.915 ;
        RECT 184.115 -158.605 184.445 -158.275 ;
        RECT 184.115 -159.965 184.445 -159.635 ;
        RECT 184.115 -161.325 184.445 -160.995 ;
        RECT 184.115 -162.685 184.445 -162.355 ;
        RECT 184.115 -164.045 184.445 -163.715 ;
        RECT 184.115 -165.405 184.445 -165.075 ;
        RECT 184.115 -166.765 184.445 -166.435 ;
        RECT 184.115 -168.125 184.445 -167.795 ;
        RECT 184.115 -169.485 184.445 -169.155 ;
        RECT 184.115 -170.845 184.445 -170.515 ;
        RECT 184.115 -172.205 184.445 -171.875 ;
        RECT 184.115 -173.565 184.445 -173.235 ;
        RECT 184.115 -174.925 184.445 -174.595 ;
        RECT 184.115 -176.285 184.445 -175.955 ;
        RECT 184.115 -177.645 184.445 -177.315 ;
        RECT 184.115 -183.29 184.445 -182.16 ;
        RECT 184.12 -183.405 184.44 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 185.475 244.04 185.805 245.17 ;
        RECT 185.475 239.875 185.805 240.205 ;
        RECT 185.475 238.515 185.805 238.845 ;
        RECT 185.475 237.155 185.805 237.485 ;
        RECT 185.48 237.155 185.8 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 185.475 -96.045 185.805 -95.715 ;
        RECT 185.475 -97.405 185.805 -97.075 ;
        RECT 185.475 -98.765 185.805 -98.435 ;
        RECT 185.475 -100.125 185.805 -99.795 ;
        RECT 185.475 -101.485 185.805 -101.155 ;
        RECT 185.475 -102.845 185.805 -102.515 ;
        RECT 185.475 -104.205 185.805 -103.875 ;
        RECT 185.475 -105.565 185.805 -105.235 ;
        RECT 185.475 -106.925 185.805 -106.595 ;
        RECT 185.475 -108.285 185.805 -107.955 ;
        RECT 185.475 -109.645 185.805 -109.315 ;
        RECT 185.475 -111.005 185.805 -110.675 ;
        RECT 185.475 -112.365 185.805 -112.035 ;
        RECT 185.475 -113.725 185.805 -113.395 ;
        RECT 185.475 -115.085 185.805 -114.755 ;
        RECT 185.475 -116.445 185.805 -116.115 ;
        RECT 185.475 -117.805 185.805 -117.475 ;
        RECT 185.475 -119.165 185.805 -118.835 ;
        RECT 185.475 -120.525 185.805 -120.195 ;
        RECT 185.475 -121.885 185.805 -121.555 ;
        RECT 185.475 -123.245 185.805 -122.915 ;
        RECT 185.475 -124.605 185.805 -124.275 ;
        RECT 185.475 -125.965 185.805 -125.635 ;
        RECT 185.475 -127.325 185.805 -126.995 ;
        RECT 185.475 -128.685 185.805 -128.355 ;
        RECT 185.475 -130.045 185.805 -129.715 ;
        RECT 185.475 -131.405 185.805 -131.075 ;
        RECT 185.475 -132.765 185.805 -132.435 ;
        RECT 185.475 -134.125 185.805 -133.795 ;
        RECT 185.475 -135.485 185.805 -135.155 ;
        RECT 185.475 -136.845 185.805 -136.515 ;
        RECT 185.475 -138.205 185.805 -137.875 ;
        RECT 185.475 -139.565 185.805 -139.235 ;
        RECT 185.475 -140.925 185.805 -140.595 ;
        RECT 185.475 -142.285 185.805 -141.955 ;
        RECT 185.475 -143.645 185.805 -143.315 ;
        RECT 185.475 -145.005 185.805 -144.675 ;
        RECT 185.475 -146.365 185.805 -146.035 ;
        RECT 185.475 -147.725 185.805 -147.395 ;
        RECT 185.475 -149.085 185.805 -148.755 ;
        RECT 185.475 -150.445 185.805 -150.115 ;
        RECT 185.475 -151.805 185.805 -151.475 ;
        RECT 185.475 -153.165 185.805 -152.835 ;
        RECT 185.475 -154.525 185.805 -154.195 ;
        RECT 185.475 -155.885 185.805 -155.555 ;
        RECT 185.475 -157.245 185.805 -156.915 ;
        RECT 185.475 -158.605 185.805 -158.275 ;
        RECT 185.475 -159.965 185.805 -159.635 ;
        RECT 185.475 -161.325 185.805 -160.995 ;
        RECT 185.475 -162.685 185.805 -162.355 ;
        RECT 185.475 -164.045 185.805 -163.715 ;
        RECT 185.475 -165.405 185.805 -165.075 ;
        RECT 185.475 -166.765 185.805 -166.435 ;
        RECT 185.475 -168.125 185.805 -167.795 ;
        RECT 185.475 -169.485 185.805 -169.155 ;
        RECT 185.475 -170.845 185.805 -170.515 ;
        RECT 185.475 -172.205 185.805 -171.875 ;
        RECT 185.475 -173.565 185.805 -173.235 ;
        RECT 185.475 -174.925 185.805 -174.595 ;
        RECT 185.475 -176.285 185.805 -175.955 ;
        RECT 185.475 -177.645 185.805 -177.315 ;
        RECT 185.475 -183.29 185.805 -182.16 ;
        RECT 185.48 -183.405 185.8 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 185.66 -94.075 185.99 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 186.835 244.04 187.165 245.17 ;
        RECT 186.835 239.875 187.165 240.205 ;
        RECT 186.835 238.515 187.165 238.845 ;
        RECT 186.835 237.155 187.165 237.485 ;
        RECT 186.84 237.155 187.16 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 188.195 244.04 188.525 245.17 ;
        RECT 188.195 239.875 188.525 240.205 ;
        RECT 188.195 238.515 188.525 238.845 ;
        RECT 188.195 237.155 188.525 237.485 ;
        RECT 188.2 237.155 188.52 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 188.195 -0.845 188.525 -0.515 ;
        RECT 188.195 -2.205 188.525 -1.875 ;
        RECT 188.195 -3.565 188.525 -3.235 ;
        RECT 188.2 -3.565 188.52 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 189.555 244.04 189.885 245.17 ;
        RECT 189.555 239.875 189.885 240.205 ;
        RECT 189.555 238.515 189.885 238.845 ;
        RECT 189.555 237.155 189.885 237.485 ;
        RECT 189.56 237.155 189.88 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 189.555 -0.845 189.885 -0.515 ;
        RECT 189.555 -2.205 189.885 -1.875 ;
        RECT 189.555 -3.565 189.885 -3.235 ;
        RECT 189.56 -3.565 189.88 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 189.555 -91.965 189.885 -91.635 ;
        RECT 189.555 -93.325 189.885 -92.995 ;
        RECT 189.555 -94.685 189.885 -94.355 ;
        RECT 189.555 -96.045 189.885 -95.715 ;
        RECT 189.555 -97.405 189.885 -97.075 ;
        RECT 189.555 -98.765 189.885 -98.435 ;
        RECT 189.555 -100.125 189.885 -99.795 ;
        RECT 189.555 -101.485 189.885 -101.155 ;
        RECT 189.555 -102.845 189.885 -102.515 ;
        RECT 189.555 -104.205 189.885 -103.875 ;
        RECT 189.555 -105.565 189.885 -105.235 ;
        RECT 189.555 -106.925 189.885 -106.595 ;
        RECT 189.555 -108.285 189.885 -107.955 ;
        RECT 189.555 -109.645 189.885 -109.315 ;
        RECT 189.555 -111.005 189.885 -110.675 ;
        RECT 189.555 -112.365 189.885 -112.035 ;
        RECT 189.555 -113.725 189.885 -113.395 ;
        RECT 189.555 -115.085 189.885 -114.755 ;
        RECT 189.555 -116.445 189.885 -116.115 ;
        RECT 189.555 -117.805 189.885 -117.475 ;
        RECT 189.555 -119.165 189.885 -118.835 ;
        RECT 189.555 -120.525 189.885 -120.195 ;
        RECT 189.555 -121.885 189.885 -121.555 ;
        RECT 189.555 -123.245 189.885 -122.915 ;
        RECT 189.555 -124.605 189.885 -124.275 ;
        RECT 189.555 -125.965 189.885 -125.635 ;
        RECT 189.555 -127.325 189.885 -126.995 ;
        RECT 189.555 -128.685 189.885 -128.355 ;
        RECT 189.555 -130.045 189.885 -129.715 ;
        RECT 189.555 -131.405 189.885 -131.075 ;
        RECT 189.555 -132.765 189.885 -132.435 ;
        RECT 189.555 -134.125 189.885 -133.795 ;
        RECT 189.555 -135.485 189.885 -135.155 ;
        RECT 189.555 -136.845 189.885 -136.515 ;
        RECT 189.555 -138.205 189.885 -137.875 ;
        RECT 189.555 -139.565 189.885 -139.235 ;
        RECT 189.555 -140.925 189.885 -140.595 ;
        RECT 189.555 -142.285 189.885 -141.955 ;
        RECT 189.555 -143.645 189.885 -143.315 ;
        RECT 189.555 -145.005 189.885 -144.675 ;
        RECT 189.555 -146.365 189.885 -146.035 ;
        RECT 189.555 -147.725 189.885 -147.395 ;
        RECT 189.555 -149.085 189.885 -148.755 ;
        RECT 189.555 -150.445 189.885 -150.115 ;
        RECT 189.555 -151.805 189.885 -151.475 ;
        RECT 189.555 -153.165 189.885 -152.835 ;
        RECT 189.555 -154.525 189.885 -154.195 ;
        RECT 189.555 -155.885 189.885 -155.555 ;
        RECT 189.555 -157.245 189.885 -156.915 ;
        RECT 189.555 -158.605 189.885 -158.275 ;
        RECT 189.555 -159.965 189.885 -159.635 ;
        RECT 189.555 -161.325 189.885 -160.995 ;
        RECT 189.555 -162.685 189.885 -162.355 ;
        RECT 189.555 -164.045 189.885 -163.715 ;
        RECT 189.555 -165.405 189.885 -165.075 ;
        RECT 189.555 -166.765 189.885 -166.435 ;
        RECT 189.555 -168.125 189.885 -167.795 ;
        RECT 189.555 -169.485 189.885 -169.155 ;
        RECT 189.555 -170.845 189.885 -170.515 ;
        RECT 189.555 -172.205 189.885 -171.875 ;
        RECT 189.555 -173.565 189.885 -173.235 ;
        RECT 189.555 -174.925 189.885 -174.595 ;
        RECT 189.555 -176.285 189.885 -175.955 ;
        RECT 189.555 -177.645 189.885 -177.315 ;
        RECT 189.555 -183.29 189.885 -182.16 ;
        RECT 189.56 -183.405 189.88 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 190.915 244.04 191.245 245.17 ;
        RECT 190.915 239.875 191.245 240.205 ;
        RECT 190.915 238.515 191.245 238.845 ;
        RECT 190.915 237.155 191.245 237.485 ;
        RECT 190.92 237.155 191.24 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 190.915 -0.845 191.245 -0.515 ;
        RECT 190.915 -2.205 191.245 -1.875 ;
        RECT 190.915 -3.565 191.245 -3.235 ;
        RECT 190.92 -3.565 191.24 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 190.915 -91.965 191.245 -91.635 ;
        RECT 190.915 -93.325 191.245 -92.995 ;
        RECT 190.915 -94.685 191.245 -94.355 ;
        RECT 190.915 -96.045 191.245 -95.715 ;
        RECT 190.915 -97.405 191.245 -97.075 ;
        RECT 190.915 -98.765 191.245 -98.435 ;
        RECT 190.915 -100.125 191.245 -99.795 ;
        RECT 190.915 -101.485 191.245 -101.155 ;
        RECT 190.915 -102.845 191.245 -102.515 ;
        RECT 190.915 -104.205 191.245 -103.875 ;
        RECT 190.915 -105.565 191.245 -105.235 ;
        RECT 190.915 -106.925 191.245 -106.595 ;
        RECT 190.915 -108.285 191.245 -107.955 ;
        RECT 190.915 -109.645 191.245 -109.315 ;
        RECT 190.915 -111.005 191.245 -110.675 ;
        RECT 190.915 -112.365 191.245 -112.035 ;
        RECT 190.915 -113.725 191.245 -113.395 ;
        RECT 190.915 -115.085 191.245 -114.755 ;
        RECT 190.915 -116.445 191.245 -116.115 ;
        RECT 190.915 -117.805 191.245 -117.475 ;
        RECT 190.915 -119.165 191.245 -118.835 ;
        RECT 190.915 -120.525 191.245 -120.195 ;
        RECT 190.915 -121.885 191.245 -121.555 ;
        RECT 190.915 -123.245 191.245 -122.915 ;
        RECT 190.915 -124.605 191.245 -124.275 ;
        RECT 190.915 -125.965 191.245 -125.635 ;
        RECT 190.915 -127.325 191.245 -126.995 ;
        RECT 190.915 -128.685 191.245 -128.355 ;
        RECT 190.915 -130.045 191.245 -129.715 ;
        RECT 190.915 -131.405 191.245 -131.075 ;
        RECT 190.915 -132.765 191.245 -132.435 ;
        RECT 190.915 -134.125 191.245 -133.795 ;
        RECT 190.915 -135.485 191.245 -135.155 ;
        RECT 190.915 -136.845 191.245 -136.515 ;
        RECT 190.915 -138.205 191.245 -137.875 ;
        RECT 190.915 -139.565 191.245 -139.235 ;
        RECT 190.915 -140.925 191.245 -140.595 ;
        RECT 190.915 -142.285 191.245 -141.955 ;
        RECT 190.915 -143.645 191.245 -143.315 ;
        RECT 190.915 -145.005 191.245 -144.675 ;
        RECT 190.915 -146.365 191.245 -146.035 ;
        RECT 190.915 -147.725 191.245 -147.395 ;
        RECT 190.915 -149.085 191.245 -148.755 ;
        RECT 190.915 -150.445 191.245 -150.115 ;
        RECT 190.915 -151.805 191.245 -151.475 ;
        RECT 190.915 -153.165 191.245 -152.835 ;
        RECT 190.915 -154.525 191.245 -154.195 ;
        RECT 190.915 -155.885 191.245 -155.555 ;
        RECT 190.915 -157.245 191.245 -156.915 ;
        RECT 190.915 -158.605 191.245 -158.275 ;
        RECT 190.915 -159.965 191.245 -159.635 ;
        RECT 190.915 -161.325 191.245 -160.995 ;
        RECT 190.915 -162.685 191.245 -162.355 ;
        RECT 190.915 -164.045 191.245 -163.715 ;
        RECT 190.915 -165.405 191.245 -165.075 ;
        RECT 190.915 -166.765 191.245 -166.435 ;
        RECT 190.915 -168.125 191.245 -167.795 ;
        RECT 190.915 -169.485 191.245 -169.155 ;
        RECT 190.915 -170.845 191.245 -170.515 ;
        RECT 190.915 -172.205 191.245 -171.875 ;
        RECT 190.915 -173.565 191.245 -173.235 ;
        RECT 190.915 -174.925 191.245 -174.595 ;
        RECT 190.915 -176.285 191.245 -175.955 ;
        RECT 190.915 -177.645 191.245 -177.315 ;
        RECT 190.915 -183.29 191.245 -182.16 ;
        RECT 190.92 -183.405 191.24 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 191.76 -94.075 192.09 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 192.275 244.04 192.605 245.17 ;
        RECT 192.275 239.875 192.605 240.205 ;
        RECT 192.275 238.515 192.605 238.845 ;
        RECT 192.275 237.155 192.605 237.485 ;
        RECT 192.28 237.155 192.6 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 192.275 -96.045 192.605 -95.715 ;
        RECT 192.275 -97.405 192.605 -97.075 ;
        RECT 192.275 -98.765 192.605 -98.435 ;
        RECT 192.275 -100.125 192.605 -99.795 ;
        RECT 192.275 -101.485 192.605 -101.155 ;
        RECT 192.275 -102.845 192.605 -102.515 ;
        RECT 192.275 -104.205 192.605 -103.875 ;
        RECT 192.275 -105.565 192.605 -105.235 ;
        RECT 192.275 -106.925 192.605 -106.595 ;
        RECT 192.275 -108.285 192.605 -107.955 ;
        RECT 192.275 -109.645 192.605 -109.315 ;
        RECT 192.275 -111.005 192.605 -110.675 ;
        RECT 192.275 -112.365 192.605 -112.035 ;
        RECT 192.275 -113.725 192.605 -113.395 ;
        RECT 192.275 -115.085 192.605 -114.755 ;
        RECT 192.275 -116.445 192.605 -116.115 ;
        RECT 192.275 -117.805 192.605 -117.475 ;
        RECT 192.275 -119.165 192.605 -118.835 ;
        RECT 192.275 -120.525 192.605 -120.195 ;
        RECT 192.275 -121.885 192.605 -121.555 ;
        RECT 192.275 -123.245 192.605 -122.915 ;
        RECT 192.275 -124.605 192.605 -124.275 ;
        RECT 192.275 -125.965 192.605 -125.635 ;
        RECT 192.275 -127.325 192.605 -126.995 ;
        RECT 192.275 -128.685 192.605 -128.355 ;
        RECT 192.275 -130.045 192.605 -129.715 ;
        RECT 192.275 -131.405 192.605 -131.075 ;
        RECT 192.275 -132.765 192.605 -132.435 ;
        RECT 192.275 -134.125 192.605 -133.795 ;
        RECT 192.275 -135.485 192.605 -135.155 ;
        RECT 192.275 -136.845 192.605 -136.515 ;
        RECT 192.275 -138.205 192.605 -137.875 ;
        RECT 192.275 -139.565 192.605 -139.235 ;
        RECT 192.275 -140.925 192.605 -140.595 ;
        RECT 192.275 -142.285 192.605 -141.955 ;
        RECT 192.275 -143.645 192.605 -143.315 ;
        RECT 192.275 -145.005 192.605 -144.675 ;
        RECT 192.275 -146.365 192.605 -146.035 ;
        RECT 192.275 -147.725 192.605 -147.395 ;
        RECT 192.275 -149.085 192.605 -148.755 ;
        RECT 192.275 -150.445 192.605 -150.115 ;
        RECT 192.275 -151.805 192.605 -151.475 ;
        RECT 192.275 -153.165 192.605 -152.835 ;
        RECT 192.275 -154.525 192.605 -154.195 ;
        RECT 192.275 -155.885 192.605 -155.555 ;
        RECT 192.275 -157.245 192.605 -156.915 ;
        RECT 192.275 -158.605 192.605 -158.275 ;
        RECT 192.275 -159.965 192.605 -159.635 ;
        RECT 192.275 -161.325 192.605 -160.995 ;
        RECT 192.275 -162.685 192.605 -162.355 ;
        RECT 192.275 -164.045 192.605 -163.715 ;
        RECT 192.275 -165.405 192.605 -165.075 ;
        RECT 192.275 -166.765 192.605 -166.435 ;
        RECT 192.275 -168.125 192.605 -167.795 ;
        RECT 192.275 -169.485 192.605 -169.155 ;
        RECT 192.275 -170.845 192.605 -170.515 ;
        RECT 192.275 -172.205 192.605 -171.875 ;
        RECT 192.275 -173.565 192.605 -173.235 ;
        RECT 192.275 -174.925 192.605 -174.595 ;
        RECT 192.275 -176.285 192.605 -175.955 ;
        RECT 192.275 -177.645 192.605 -177.315 ;
        RECT 192.275 -183.29 192.605 -182.16 ;
        RECT 192.28 -183.405 192.6 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 193.635 244.04 193.965 245.17 ;
        RECT 193.635 239.875 193.965 240.205 ;
        RECT 193.635 238.515 193.965 238.845 ;
        RECT 193.635 237.155 193.965 237.485 ;
        RECT 193.64 237.155 193.96 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 193.635 -0.845 193.965 -0.515 ;
        RECT 193.635 -2.205 193.965 -1.875 ;
        RECT 193.635 -3.565 193.965 -3.235 ;
        RECT 193.64 -3.565 193.96 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 194.995 244.04 195.325 245.17 ;
        RECT 194.995 239.875 195.325 240.205 ;
        RECT 194.995 238.515 195.325 238.845 ;
        RECT 194.995 237.155 195.325 237.485 ;
        RECT 195 237.155 195.32 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 194.995 -0.845 195.325 -0.515 ;
        RECT 194.995 -2.205 195.325 -1.875 ;
        RECT 194.995 -3.565 195.325 -3.235 ;
        RECT 195 -3.565 195.32 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 196.355 244.04 196.685 245.17 ;
        RECT 196.355 239.875 196.685 240.205 ;
        RECT 196.355 238.515 196.685 238.845 ;
        RECT 196.355 237.155 196.685 237.485 ;
        RECT 196.36 237.155 196.68 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 196.355 -0.845 196.685 -0.515 ;
        RECT 196.355 -2.205 196.685 -1.875 ;
        RECT 196.355 -3.565 196.685 -3.235 ;
        RECT 196.36 -3.565 196.68 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 196.355 -91.965 196.685 -91.635 ;
        RECT 196.355 -93.325 196.685 -92.995 ;
        RECT 196.355 -94.685 196.685 -94.355 ;
        RECT 196.355 -96.045 196.685 -95.715 ;
        RECT 196.355 -97.405 196.685 -97.075 ;
        RECT 196.355 -98.765 196.685 -98.435 ;
        RECT 196.355 -100.125 196.685 -99.795 ;
        RECT 196.355 -101.485 196.685 -101.155 ;
        RECT 196.355 -102.845 196.685 -102.515 ;
        RECT 196.355 -104.205 196.685 -103.875 ;
        RECT 196.355 -105.565 196.685 -105.235 ;
        RECT 196.355 -106.925 196.685 -106.595 ;
        RECT 196.355 -108.285 196.685 -107.955 ;
        RECT 196.355 -109.645 196.685 -109.315 ;
        RECT 196.355 -111.005 196.685 -110.675 ;
        RECT 196.355 -112.365 196.685 -112.035 ;
        RECT 196.355 -113.725 196.685 -113.395 ;
        RECT 196.355 -115.085 196.685 -114.755 ;
        RECT 196.355 -116.445 196.685 -116.115 ;
        RECT 196.355 -117.805 196.685 -117.475 ;
        RECT 196.355 -119.165 196.685 -118.835 ;
        RECT 196.355 -120.525 196.685 -120.195 ;
        RECT 196.355 -121.885 196.685 -121.555 ;
        RECT 196.355 -123.245 196.685 -122.915 ;
        RECT 196.355 -124.605 196.685 -124.275 ;
        RECT 196.355 -125.965 196.685 -125.635 ;
        RECT 196.355 -127.325 196.685 -126.995 ;
        RECT 196.355 -128.685 196.685 -128.355 ;
        RECT 196.355 -130.045 196.685 -129.715 ;
        RECT 196.355 -131.405 196.685 -131.075 ;
        RECT 196.355 -132.765 196.685 -132.435 ;
        RECT 196.355 -134.125 196.685 -133.795 ;
        RECT 196.355 -135.485 196.685 -135.155 ;
        RECT 196.355 -136.845 196.685 -136.515 ;
        RECT 196.355 -138.205 196.685 -137.875 ;
        RECT 196.355 -139.565 196.685 -139.235 ;
        RECT 196.355 -140.925 196.685 -140.595 ;
        RECT 196.355 -142.285 196.685 -141.955 ;
        RECT 196.355 -143.645 196.685 -143.315 ;
        RECT 196.355 -145.005 196.685 -144.675 ;
        RECT 196.355 -146.365 196.685 -146.035 ;
        RECT 196.355 -147.725 196.685 -147.395 ;
        RECT 196.355 -149.085 196.685 -148.755 ;
        RECT 196.355 -150.445 196.685 -150.115 ;
        RECT 196.355 -151.805 196.685 -151.475 ;
        RECT 196.355 -153.165 196.685 -152.835 ;
        RECT 196.355 -154.525 196.685 -154.195 ;
        RECT 196.355 -155.885 196.685 -155.555 ;
        RECT 196.355 -157.245 196.685 -156.915 ;
        RECT 196.355 -158.605 196.685 -158.275 ;
        RECT 196.355 -159.965 196.685 -159.635 ;
        RECT 196.355 -161.325 196.685 -160.995 ;
        RECT 196.355 -162.685 196.685 -162.355 ;
        RECT 196.355 -164.045 196.685 -163.715 ;
        RECT 196.355 -165.405 196.685 -165.075 ;
        RECT 196.355 -166.765 196.685 -166.435 ;
        RECT 196.355 -168.125 196.685 -167.795 ;
        RECT 196.355 -169.485 196.685 -169.155 ;
        RECT 196.355 -170.845 196.685 -170.515 ;
        RECT 196.355 -172.205 196.685 -171.875 ;
        RECT 196.355 -173.565 196.685 -173.235 ;
        RECT 196.355 -174.925 196.685 -174.595 ;
        RECT 196.355 -176.285 196.685 -175.955 ;
        RECT 196.355 -177.645 196.685 -177.315 ;
        RECT 196.355 -183.29 196.685 -182.16 ;
        RECT 196.36 -183.405 196.68 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 197.715 244.04 198.045 245.17 ;
        RECT 197.715 239.875 198.045 240.205 ;
        RECT 197.715 238.515 198.045 238.845 ;
        RECT 197.715 237.155 198.045 237.485 ;
        RECT 197.72 237.155 198.04 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 197.715 -96.045 198.045 -95.715 ;
        RECT 197.715 -97.405 198.045 -97.075 ;
        RECT 197.715 -98.765 198.045 -98.435 ;
        RECT 197.715 -100.125 198.045 -99.795 ;
        RECT 197.715 -101.485 198.045 -101.155 ;
        RECT 197.715 -102.845 198.045 -102.515 ;
        RECT 197.715 -104.205 198.045 -103.875 ;
        RECT 197.715 -105.565 198.045 -105.235 ;
        RECT 197.715 -106.925 198.045 -106.595 ;
        RECT 197.715 -108.285 198.045 -107.955 ;
        RECT 197.715 -109.645 198.045 -109.315 ;
        RECT 197.715 -111.005 198.045 -110.675 ;
        RECT 197.715 -112.365 198.045 -112.035 ;
        RECT 197.715 -113.725 198.045 -113.395 ;
        RECT 197.715 -115.085 198.045 -114.755 ;
        RECT 197.715 -116.445 198.045 -116.115 ;
        RECT 197.715 -117.805 198.045 -117.475 ;
        RECT 197.715 -119.165 198.045 -118.835 ;
        RECT 197.715 -120.525 198.045 -120.195 ;
        RECT 197.715 -121.885 198.045 -121.555 ;
        RECT 197.715 -123.245 198.045 -122.915 ;
        RECT 197.715 -124.605 198.045 -124.275 ;
        RECT 197.715 -125.965 198.045 -125.635 ;
        RECT 197.715 -127.325 198.045 -126.995 ;
        RECT 197.715 -128.685 198.045 -128.355 ;
        RECT 197.715 -130.045 198.045 -129.715 ;
        RECT 197.715 -131.405 198.045 -131.075 ;
        RECT 197.715 -132.765 198.045 -132.435 ;
        RECT 197.715 -134.125 198.045 -133.795 ;
        RECT 197.715 -135.485 198.045 -135.155 ;
        RECT 197.715 -136.845 198.045 -136.515 ;
        RECT 197.715 -138.205 198.045 -137.875 ;
        RECT 197.715 -139.565 198.045 -139.235 ;
        RECT 197.715 -140.925 198.045 -140.595 ;
        RECT 197.715 -142.285 198.045 -141.955 ;
        RECT 197.715 -143.645 198.045 -143.315 ;
        RECT 197.715 -145.005 198.045 -144.675 ;
        RECT 197.715 -146.365 198.045 -146.035 ;
        RECT 197.715 -147.725 198.045 -147.395 ;
        RECT 197.715 -149.085 198.045 -148.755 ;
        RECT 197.715 -150.445 198.045 -150.115 ;
        RECT 197.715 -151.805 198.045 -151.475 ;
        RECT 197.715 -153.165 198.045 -152.835 ;
        RECT 197.715 -154.525 198.045 -154.195 ;
        RECT 197.715 -155.885 198.045 -155.555 ;
        RECT 197.715 -157.245 198.045 -156.915 ;
        RECT 197.715 -158.605 198.045 -158.275 ;
        RECT 197.715 -159.965 198.045 -159.635 ;
        RECT 197.715 -161.325 198.045 -160.995 ;
        RECT 197.715 -162.685 198.045 -162.355 ;
        RECT 197.715 -164.045 198.045 -163.715 ;
        RECT 197.715 -165.405 198.045 -165.075 ;
        RECT 197.715 -166.765 198.045 -166.435 ;
        RECT 197.715 -168.125 198.045 -167.795 ;
        RECT 197.715 -169.485 198.045 -169.155 ;
        RECT 197.715 -170.845 198.045 -170.515 ;
        RECT 197.715 -172.205 198.045 -171.875 ;
        RECT 197.715 -173.565 198.045 -173.235 ;
        RECT 197.715 -174.925 198.045 -174.595 ;
        RECT 197.715 -176.285 198.045 -175.955 ;
        RECT 197.715 -177.645 198.045 -177.315 ;
        RECT 197.715 -183.29 198.045 -182.16 ;
        RECT 197.72 -183.405 198.04 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 197.86 -94.075 198.19 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 199.075 244.04 199.405 245.17 ;
        RECT 199.075 239.875 199.405 240.205 ;
        RECT 199.075 238.515 199.405 238.845 ;
        RECT 199.075 237.155 199.405 237.485 ;
        RECT 199.08 237.155 199.4 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 200.435 244.04 200.765 245.17 ;
        RECT 200.435 239.875 200.765 240.205 ;
        RECT 200.435 238.515 200.765 238.845 ;
        RECT 200.435 237.155 200.765 237.485 ;
        RECT 200.44 237.155 200.76 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 200.435 -0.845 200.765 -0.515 ;
        RECT 200.435 -2.205 200.765 -1.875 ;
        RECT 200.435 -3.565 200.765 -3.235 ;
        RECT 200.44 -3.565 200.76 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 201.795 244.04 202.125 245.17 ;
        RECT 201.795 239.875 202.125 240.205 ;
        RECT 201.795 238.515 202.125 238.845 ;
        RECT 201.795 237.155 202.125 237.485 ;
        RECT 201.8 237.155 202.12 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 201.795 -0.845 202.125 -0.515 ;
        RECT 201.795 -2.205 202.125 -1.875 ;
        RECT 201.795 -3.565 202.125 -3.235 ;
        RECT 201.8 -3.565 202.12 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 203.155 244.04 203.485 245.17 ;
        RECT 203.155 239.875 203.485 240.205 ;
        RECT 203.155 238.515 203.485 238.845 ;
        RECT 203.155 237.155 203.485 237.485 ;
        RECT 203.16 237.155 203.48 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 203.155 -0.845 203.485 -0.515 ;
        RECT 203.155 -2.205 203.485 -1.875 ;
        RECT 203.155 -3.565 203.485 -3.235 ;
        RECT 203.16 -3.565 203.48 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 203.155 -98.765 203.485 -98.435 ;
        RECT 203.155 -100.125 203.485 -99.795 ;
        RECT 203.155 -101.485 203.485 -101.155 ;
        RECT 203.155 -102.845 203.485 -102.515 ;
        RECT 203.155 -104.205 203.485 -103.875 ;
        RECT 203.155 -105.565 203.485 -105.235 ;
        RECT 203.155 -106.925 203.485 -106.595 ;
        RECT 203.155 -108.285 203.485 -107.955 ;
        RECT 203.155 -109.645 203.485 -109.315 ;
        RECT 203.155 -111.005 203.485 -110.675 ;
        RECT 203.155 -112.365 203.485 -112.035 ;
        RECT 203.155 -113.725 203.485 -113.395 ;
        RECT 203.155 -115.085 203.485 -114.755 ;
        RECT 203.155 -116.445 203.485 -116.115 ;
        RECT 203.155 -117.805 203.485 -117.475 ;
        RECT 203.155 -119.165 203.485 -118.835 ;
        RECT 203.155 -120.525 203.485 -120.195 ;
        RECT 203.155 -121.885 203.485 -121.555 ;
        RECT 203.155 -123.245 203.485 -122.915 ;
        RECT 203.155 -124.605 203.485 -124.275 ;
        RECT 203.155 -125.965 203.485 -125.635 ;
        RECT 203.155 -127.325 203.485 -126.995 ;
        RECT 203.155 -128.685 203.485 -128.355 ;
        RECT 203.155 -130.045 203.485 -129.715 ;
        RECT 203.155 -131.405 203.485 -131.075 ;
        RECT 203.155 -132.765 203.485 -132.435 ;
        RECT 203.155 -134.125 203.485 -133.795 ;
        RECT 203.155 -135.485 203.485 -135.155 ;
        RECT 203.155 -136.845 203.485 -136.515 ;
        RECT 203.155 -138.205 203.485 -137.875 ;
        RECT 203.155 -139.565 203.485 -139.235 ;
        RECT 203.155 -140.925 203.485 -140.595 ;
        RECT 203.155 -142.285 203.485 -141.955 ;
        RECT 203.155 -143.645 203.485 -143.315 ;
        RECT 203.155 -145.005 203.485 -144.675 ;
        RECT 203.155 -146.365 203.485 -146.035 ;
        RECT 203.155 -147.725 203.485 -147.395 ;
        RECT 203.155 -149.085 203.485 -148.755 ;
        RECT 203.155 -150.445 203.485 -150.115 ;
        RECT 203.155 -151.805 203.485 -151.475 ;
        RECT 203.155 -153.165 203.485 -152.835 ;
        RECT 203.155 -154.525 203.485 -154.195 ;
        RECT 203.155 -155.885 203.485 -155.555 ;
        RECT 203.155 -157.245 203.485 -156.915 ;
        RECT 203.155 -158.605 203.485 -158.275 ;
        RECT 203.155 -159.965 203.485 -159.635 ;
        RECT 203.155 -161.325 203.485 -160.995 ;
        RECT 203.155 -162.685 203.485 -162.355 ;
        RECT 203.155 -164.045 203.485 -163.715 ;
        RECT 203.155 -165.405 203.485 -165.075 ;
        RECT 203.155 -166.765 203.485 -166.435 ;
        RECT 203.155 -168.125 203.485 -167.795 ;
        RECT 203.155 -169.485 203.485 -169.155 ;
        RECT 203.155 -170.845 203.485 -170.515 ;
        RECT 203.155 -172.205 203.485 -171.875 ;
        RECT 203.155 -173.565 203.485 -173.235 ;
        RECT 203.155 -174.925 203.485 -174.595 ;
        RECT 203.155 -176.285 203.485 -175.955 ;
        RECT 203.155 -177.645 203.485 -177.315 ;
        RECT 203.155 -183.29 203.485 -182.16 ;
        RECT 203.16 -183.405 203.48 -90.96 ;
        RECT 203.155 -91.965 203.485 -91.635 ;
        RECT 203.155 -93.325 203.485 -92.995 ;
        RECT 203.155 -94.685 203.485 -94.355 ;
        RECT 203.155 -96.045 203.485 -95.715 ;
        RECT 203.155 -97.405 203.485 -97.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 139.235 244.04 139.565 245.17 ;
        RECT 139.235 239.875 139.565 240.205 ;
        RECT 139.235 238.515 139.565 238.845 ;
        RECT 139.235 237.155 139.565 237.485 ;
        RECT 139.24 237.155 139.56 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 139.235 -0.845 139.565 -0.515 ;
        RECT 139.235 -2.205 139.565 -1.875 ;
        RECT 139.235 -3.565 139.565 -3.235 ;
        RECT 139.24 -3.565 139.56 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 140.595 244.04 140.925 245.17 ;
        RECT 140.595 239.875 140.925 240.205 ;
        RECT 140.595 238.515 140.925 238.845 ;
        RECT 140.595 237.155 140.925 237.485 ;
        RECT 140.6 237.155 140.92 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 140.595 -0.845 140.925 -0.515 ;
        RECT 140.595 -2.205 140.925 -1.875 ;
        RECT 140.595 -3.565 140.925 -3.235 ;
        RECT 140.6 -3.565 140.92 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 140.595 -91.965 140.925 -91.635 ;
        RECT 140.595 -93.325 140.925 -92.995 ;
        RECT 140.595 -94.685 140.925 -94.355 ;
        RECT 140.595 -96.045 140.925 -95.715 ;
        RECT 140.595 -97.405 140.925 -97.075 ;
        RECT 140.595 -98.765 140.925 -98.435 ;
        RECT 140.595 -100.125 140.925 -99.795 ;
        RECT 140.595 -101.485 140.925 -101.155 ;
        RECT 140.595 -102.845 140.925 -102.515 ;
        RECT 140.595 -104.205 140.925 -103.875 ;
        RECT 140.595 -105.565 140.925 -105.235 ;
        RECT 140.595 -106.925 140.925 -106.595 ;
        RECT 140.595 -108.285 140.925 -107.955 ;
        RECT 140.595 -109.645 140.925 -109.315 ;
        RECT 140.595 -111.005 140.925 -110.675 ;
        RECT 140.595 -112.365 140.925 -112.035 ;
        RECT 140.595 -113.725 140.925 -113.395 ;
        RECT 140.595 -115.085 140.925 -114.755 ;
        RECT 140.595 -116.445 140.925 -116.115 ;
        RECT 140.595 -117.805 140.925 -117.475 ;
        RECT 140.595 -119.165 140.925 -118.835 ;
        RECT 140.595 -120.525 140.925 -120.195 ;
        RECT 140.595 -121.885 140.925 -121.555 ;
        RECT 140.595 -123.245 140.925 -122.915 ;
        RECT 140.595 -124.605 140.925 -124.275 ;
        RECT 140.595 -125.965 140.925 -125.635 ;
        RECT 140.595 -127.325 140.925 -126.995 ;
        RECT 140.595 -128.685 140.925 -128.355 ;
        RECT 140.595 -130.045 140.925 -129.715 ;
        RECT 140.595 -131.405 140.925 -131.075 ;
        RECT 140.595 -132.765 140.925 -132.435 ;
        RECT 140.595 -134.125 140.925 -133.795 ;
        RECT 140.595 -135.485 140.925 -135.155 ;
        RECT 140.595 -136.845 140.925 -136.515 ;
        RECT 140.595 -138.205 140.925 -137.875 ;
        RECT 140.595 -139.565 140.925 -139.235 ;
        RECT 140.595 -140.925 140.925 -140.595 ;
        RECT 140.595 -142.285 140.925 -141.955 ;
        RECT 140.595 -143.645 140.925 -143.315 ;
        RECT 140.595 -145.005 140.925 -144.675 ;
        RECT 140.595 -146.365 140.925 -146.035 ;
        RECT 140.595 -147.725 140.925 -147.395 ;
        RECT 140.595 -149.085 140.925 -148.755 ;
        RECT 140.595 -150.445 140.925 -150.115 ;
        RECT 140.595 -151.805 140.925 -151.475 ;
        RECT 140.595 -153.165 140.925 -152.835 ;
        RECT 140.595 -154.525 140.925 -154.195 ;
        RECT 140.595 -155.885 140.925 -155.555 ;
        RECT 140.595 -157.245 140.925 -156.915 ;
        RECT 140.595 -158.605 140.925 -158.275 ;
        RECT 140.595 -159.965 140.925 -159.635 ;
        RECT 140.595 -161.325 140.925 -160.995 ;
        RECT 140.595 -162.685 140.925 -162.355 ;
        RECT 140.595 -164.045 140.925 -163.715 ;
        RECT 140.595 -165.405 140.925 -165.075 ;
        RECT 140.595 -166.765 140.925 -166.435 ;
        RECT 140.595 -168.125 140.925 -167.795 ;
        RECT 140.595 -169.485 140.925 -169.155 ;
        RECT 140.595 -170.845 140.925 -170.515 ;
        RECT 140.595 -172.205 140.925 -171.875 ;
        RECT 140.595 -173.565 140.925 -173.235 ;
        RECT 140.595 -174.925 140.925 -174.595 ;
        RECT 140.595 -176.285 140.925 -175.955 ;
        RECT 140.595 -177.645 140.925 -177.315 ;
        RECT 140.595 -183.29 140.925 -182.16 ;
        RECT 140.6 -183.405 140.92 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 141.955 244.04 142.285 245.17 ;
        RECT 141.955 239.875 142.285 240.205 ;
        RECT 141.955 238.515 142.285 238.845 ;
        RECT 141.955 237.155 142.285 237.485 ;
        RECT 141.96 237.155 142.28 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 141.955 -0.845 142.285 -0.515 ;
        RECT 141.955 -2.205 142.285 -1.875 ;
        RECT 141.955 -3.565 142.285 -3.235 ;
        RECT 141.96 -3.565 142.28 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 141.955 -91.965 142.285 -91.635 ;
        RECT 141.955 -93.325 142.285 -92.995 ;
        RECT 141.955 -94.685 142.285 -94.355 ;
        RECT 141.955 -96.045 142.285 -95.715 ;
        RECT 141.955 -97.405 142.285 -97.075 ;
        RECT 141.955 -98.765 142.285 -98.435 ;
        RECT 141.955 -100.125 142.285 -99.795 ;
        RECT 141.955 -101.485 142.285 -101.155 ;
        RECT 141.955 -102.845 142.285 -102.515 ;
        RECT 141.955 -104.205 142.285 -103.875 ;
        RECT 141.955 -105.565 142.285 -105.235 ;
        RECT 141.955 -106.925 142.285 -106.595 ;
        RECT 141.955 -108.285 142.285 -107.955 ;
        RECT 141.955 -109.645 142.285 -109.315 ;
        RECT 141.955 -111.005 142.285 -110.675 ;
        RECT 141.955 -112.365 142.285 -112.035 ;
        RECT 141.955 -113.725 142.285 -113.395 ;
        RECT 141.955 -115.085 142.285 -114.755 ;
        RECT 141.955 -116.445 142.285 -116.115 ;
        RECT 141.955 -117.805 142.285 -117.475 ;
        RECT 141.955 -119.165 142.285 -118.835 ;
        RECT 141.955 -120.525 142.285 -120.195 ;
        RECT 141.955 -121.885 142.285 -121.555 ;
        RECT 141.955 -123.245 142.285 -122.915 ;
        RECT 141.955 -124.605 142.285 -124.275 ;
        RECT 141.955 -125.965 142.285 -125.635 ;
        RECT 141.955 -127.325 142.285 -126.995 ;
        RECT 141.955 -128.685 142.285 -128.355 ;
        RECT 141.955 -130.045 142.285 -129.715 ;
        RECT 141.955 -131.405 142.285 -131.075 ;
        RECT 141.955 -132.765 142.285 -132.435 ;
        RECT 141.955 -134.125 142.285 -133.795 ;
        RECT 141.955 -135.485 142.285 -135.155 ;
        RECT 141.955 -136.845 142.285 -136.515 ;
        RECT 141.955 -138.205 142.285 -137.875 ;
        RECT 141.955 -139.565 142.285 -139.235 ;
        RECT 141.955 -140.925 142.285 -140.595 ;
        RECT 141.955 -142.285 142.285 -141.955 ;
        RECT 141.955 -143.645 142.285 -143.315 ;
        RECT 141.955 -145.005 142.285 -144.675 ;
        RECT 141.955 -146.365 142.285 -146.035 ;
        RECT 141.955 -147.725 142.285 -147.395 ;
        RECT 141.955 -149.085 142.285 -148.755 ;
        RECT 141.955 -150.445 142.285 -150.115 ;
        RECT 141.955 -151.805 142.285 -151.475 ;
        RECT 141.955 -153.165 142.285 -152.835 ;
        RECT 141.955 -154.525 142.285 -154.195 ;
        RECT 141.955 -155.885 142.285 -155.555 ;
        RECT 141.955 -157.245 142.285 -156.915 ;
        RECT 141.955 -158.605 142.285 -158.275 ;
        RECT 141.955 -159.965 142.285 -159.635 ;
        RECT 141.955 -161.325 142.285 -160.995 ;
        RECT 141.955 -162.685 142.285 -162.355 ;
        RECT 141.955 -164.045 142.285 -163.715 ;
        RECT 141.955 -165.405 142.285 -165.075 ;
        RECT 141.955 -166.765 142.285 -166.435 ;
        RECT 141.955 -168.125 142.285 -167.795 ;
        RECT 141.955 -169.485 142.285 -169.155 ;
        RECT 141.955 -170.845 142.285 -170.515 ;
        RECT 141.955 -172.205 142.285 -171.875 ;
        RECT 141.955 -173.565 142.285 -173.235 ;
        RECT 141.955 -174.925 142.285 -174.595 ;
        RECT 141.955 -176.285 142.285 -175.955 ;
        RECT 141.955 -177.645 142.285 -177.315 ;
        RECT 141.955 -183.29 142.285 -182.16 ;
        RECT 141.96 -183.405 142.28 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 142.96 -94.075 143.29 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 143.315 244.04 143.645 245.17 ;
        RECT 143.315 239.875 143.645 240.205 ;
        RECT 143.315 238.515 143.645 238.845 ;
        RECT 143.315 237.155 143.645 237.485 ;
        RECT 143.32 237.155 143.64 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 143.315 -96.045 143.645 -95.715 ;
        RECT 143.315 -97.405 143.645 -97.075 ;
        RECT 143.315 -98.765 143.645 -98.435 ;
        RECT 143.315 -100.125 143.645 -99.795 ;
        RECT 143.315 -101.485 143.645 -101.155 ;
        RECT 143.315 -102.845 143.645 -102.515 ;
        RECT 143.315 -104.205 143.645 -103.875 ;
        RECT 143.315 -105.565 143.645 -105.235 ;
        RECT 143.315 -106.925 143.645 -106.595 ;
        RECT 143.315 -108.285 143.645 -107.955 ;
        RECT 143.315 -109.645 143.645 -109.315 ;
        RECT 143.315 -111.005 143.645 -110.675 ;
        RECT 143.315 -112.365 143.645 -112.035 ;
        RECT 143.315 -113.725 143.645 -113.395 ;
        RECT 143.315 -115.085 143.645 -114.755 ;
        RECT 143.315 -116.445 143.645 -116.115 ;
        RECT 143.315 -117.805 143.645 -117.475 ;
        RECT 143.315 -119.165 143.645 -118.835 ;
        RECT 143.315 -120.525 143.645 -120.195 ;
        RECT 143.315 -121.885 143.645 -121.555 ;
        RECT 143.315 -123.245 143.645 -122.915 ;
        RECT 143.315 -124.605 143.645 -124.275 ;
        RECT 143.315 -125.965 143.645 -125.635 ;
        RECT 143.315 -127.325 143.645 -126.995 ;
        RECT 143.315 -128.685 143.645 -128.355 ;
        RECT 143.315 -130.045 143.645 -129.715 ;
        RECT 143.315 -131.405 143.645 -131.075 ;
        RECT 143.315 -132.765 143.645 -132.435 ;
        RECT 143.315 -134.125 143.645 -133.795 ;
        RECT 143.315 -135.485 143.645 -135.155 ;
        RECT 143.315 -136.845 143.645 -136.515 ;
        RECT 143.315 -138.205 143.645 -137.875 ;
        RECT 143.315 -139.565 143.645 -139.235 ;
        RECT 143.315 -140.925 143.645 -140.595 ;
        RECT 143.315 -142.285 143.645 -141.955 ;
        RECT 143.315 -143.645 143.645 -143.315 ;
        RECT 143.315 -145.005 143.645 -144.675 ;
        RECT 143.315 -146.365 143.645 -146.035 ;
        RECT 143.315 -147.725 143.645 -147.395 ;
        RECT 143.315 -149.085 143.645 -148.755 ;
        RECT 143.315 -150.445 143.645 -150.115 ;
        RECT 143.315 -151.805 143.645 -151.475 ;
        RECT 143.315 -153.165 143.645 -152.835 ;
        RECT 143.315 -154.525 143.645 -154.195 ;
        RECT 143.315 -155.885 143.645 -155.555 ;
        RECT 143.315 -157.245 143.645 -156.915 ;
        RECT 143.315 -158.605 143.645 -158.275 ;
        RECT 143.315 -159.965 143.645 -159.635 ;
        RECT 143.315 -161.325 143.645 -160.995 ;
        RECT 143.315 -162.685 143.645 -162.355 ;
        RECT 143.315 -164.045 143.645 -163.715 ;
        RECT 143.315 -165.405 143.645 -165.075 ;
        RECT 143.315 -166.765 143.645 -166.435 ;
        RECT 143.315 -168.125 143.645 -167.795 ;
        RECT 143.315 -169.485 143.645 -169.155 ;
        RECT 143.315 -170.845 143.645 -170.515 ;
        RECT 143.315 -172.205 143.645 -171.875 ;
        RECT 143.315 -173.565 143.645 -173.235 ;
        RECT 143.315 -174.925 143.645 -174.595 ;
        RECT 143.315 -176.285 143.645 -175.955 ;
        RECT 143.315 -177.645 143.645 -177.315 ;
        RECT 143.315 -183.29 143.645 -182.16 ;
        RECT 143.32 -183.405 143.64 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 144.675 244.04 145.005 245.17 ;
        RECT 144.675 239.875 145.005 240.205 ;
        RECT 144.675 238.515 145.005 238.845 ;
        RECT 144.675 237.155 145.005 237.485 ;
        RECT 144.68 237.155 145 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 144.675 -0.845 145.005 -0.515 ;
        RECT 144.675 -2.205 145.005 -1.875 ;
        RECT 144.675 -3.565 145.005 -3.235 ;
        RECT 144.68 -3.565 145 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 146.035 244.04 146.365 245.17 ;
        RECT 146.035 239.875 146.365 240.205 ;
        RECT 146.035 238.515 146.365 238.845 ;
        RECT 146.035 237.155 146.365 237.485 ;
        RECT 146.04 237.155 146.36 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 146.035 -0.845 146.365 -0.515 ;
        RECT 146.035 -2.205 146.365 -1.875 ;
        RECT 146.035 -3.565 146.365 -3.235 ;
        RECT 146.04 -3.565 146.36 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 147.395 244.04 147.725 245.17 ;
        RECT 147.395 239.875 147.725 240.205 ;
        RECT 147.395 238.515 147.725 238.845 ;
        RECT 147.395 237.155 147.725 237.485 ;
        RECT 147.4 237.155 147.72 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 147.395 -0.845 147.725 -0.515 ;
        RECT 147.395 -2.205 147.725 -1.875 ;
        RECT 147.395 -3.565 147.725 -3.235 ;
        RECT 147.4 -3.565 147.72 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 147.395 -91.965 147.725 -91.635 ;
        RECT 147.395 -93.325 147.725 -92.995 ;
        RECT 147.395 -94.685 147.725 -94.355 ;
        RECT 147.395 -96.045 147.725 -95.715 ;
        RECT 147.395 -97.405 147.725 -97.075 ;
        RECT 147.395 -98.765 147.725 -98.435 ;
        RECT 147.395 -100.125 147.725 -99.795 ;
        RECT 147.395 -101.485 147.725 -101.155 ;
        RECT 147.395 -102.845 147.725 -102.515 ;
        RECT 147.395 -104.205 147.725 -103.875 ;
        RECT 147.395 -105.565 147.725 -105.235 ;
        RECT 147.395 -106.925 147.725 -106.595 ;
        RECT 147.395 -108.285 147.725 -107.955 ;
        RECT 147.395 -109.645 147.725 -109.315 ;
        RECT 147.395 -111.005 147.725 -110.675 ;
        RECT 147.395 -112.365 147.725 -112.035 ;
        RECT 147.395 -113.725 147.725 -113.395 ;
        RECT 147.395 -115.085 147.725 -114.755 ;
        RECT 147.395 -116.445 147.725 -116.115 ;
        RECT 147.395 -117.805 147.725 -117.475 ;
        RECT 147.395 -119.165 147.725 -118.835 ;
        RECT 147.395 -120.525 147.725 -120.195 ;
        RECT 147.395 -121.885 147.725 -121.555 ;
        RECT 147.395 -123.245 147.725 -122.915 ;
        RECT 147.395 -124.605 147.725 -124.275 ;
        RECT 147.395 -125.965 147.725 -125.635 ;
        RECT 147.395 -127.325 147.725 -126.995 ;
        RECT 147.395 -128.685 147.725 -128.355 ;
        RECT 147.395 -130.045 147.725 -129.715 ;
        RECT 147.395 -131.405 147.725 -131.075 ;
        RECT 147.395 -132.765 147.725 -132.435 ;
        RECT 147.395 -134.125 147.725 -133.795 ;
        RECT 147.395 -135.485 147.725 -135.155 ;
        RECT 147.395 -136.845 147.725 -136.515 ;
        RECT 147.395 -138.205 147.725 -137.875 ;
        RECT 147.395 -139.565 147.725 -139.235 ;
        RECT 147.395 -140.925 147.725 -140.595 ;
        RECT 147.395 -142.285 147.725 -141.955 ;
        RECT 147.395 -143.645 147.725 -143.315 ;
        RECT 147.395 -145.005 147.725 -144.675 ;
        RECT 147.395 -146.365 147.725 -146.035 ;
        RECT 147.395 -147.725 147.725 -147.395 ;
        RECT 147.395 -149.085 147.725 -148.755 ;
        RECT 147.395 -150.445 147.725 -150.115 ;
        RECT 147.395 -151.805 147.725 -151.475 ;
        RECT 147.395 -153.165 147.725 -152.835 ;
        RECT 147.395 -154.525 147.725 -154.195 ;
        RECT 147.395 -155.885 147.725 -155.555 ;
        RECT 147.395 -157.245 147.725 -156.915 ;
        RECT 147.395 -158.605 147.725 -158.275 ;
        RECT 147.395 -159.965 147.725 -159.635 ;
        RECT 147.395 -161.325 147.725 -160.995 ;
        RECT 147.395 -162.685 147.725 -162.355 ;
        RECT 147.395 -164.045 147.725 -163.715 ;
        RECT 147.395 -165.405 147.725 -165.075 ;
        RECT 147.395 -166.765 147.725 -166.435 ;
        RECT 147.395 -168.125 147.725 -167.795 ;
        RECT 147.395 -169.485 147.725 -169.155 ;
        RECT 147.395 -170.845 147.725 -170.515 ;
        RECT 147.395 -172.205 147.725 -171.875 ;
        RECT 147.395 -173.565 147.725 -173.235 ;
        RECT 147.395 -174.925 147.725 -174.595 ;
        RECT 147.395 -176.285 147.725 -175.955 ;
        RECT 147.395 -177.645 147.725 -177.315 ;
        RECT 147.395 -183.29 147.725 -182.16 ;
        RECT 147.4 -183.405 147.72 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 148.755 244.04 149.085 245.17 ;
        RECT 148.755 239.875 149.085 240.205 ;
        RECT 148.755 238.515 149.085 238.845 ;
        RECT 148.755 237.155 149.085 237.485 ;
        RECT 148.76 237.155 149.08 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 148.755 -96.045 149.085 -95.715 ;
        RECT 148.755 -97.405 149.085 -97.075 ;
        RECT 148.755 -98.765 149.085 -98.435 ;
        RECT 148.755 -100.125 149.085 -99.795 ;
        RECT 148.755 -101.485 149.085 -101.155 ;
        RECT 148.755 -102.845 149.085 -102.515 ;
        RECT 148.755 -104.205 149.085 -103.875 ;
        RECT 148.755 -105.565 149.085 -105.235 ;
        RECT 148.755 -106.925 149.085 -106.595 ;
        RECT 148.755 -108.285 149.085 -107.955 ;
        RECT 148.755 -109.645 149.085 -109.315 ;
        RECT 148.755 -111.005 149.085 -110.675 ;
        RECT 148.755 -112.365 149.085 -112.035 ;
        RECT 148.755 -113.725 149.085 -113.395 ;
        RECT 148.755 -115.085 149.085 -114.755 ;
        RECT 148.755 -116.445 149.085 -116.115 ;
        RECT 148.755 -117.805 149.085 -117.475 ;
        RECT 148.755 -119.165 149.085 -118.835 ;
        RECT 148.755 -120.525 149.085 -120.195 ;
        RECT 148.755 -121.885 149.085 -121.555 ;
        RECT 148.755 -123.245 149.085 -122.915 ;
        RECT 148.755 -124.605 149.085 -124.275 ;
        RECT 148.755 -125.965 149.085 -125.635 ;
        RECT 148.755 -127.325 149.085 -126.995 ;
        RECT 148.755 -128.685 149.085 -128.355 ;
        RECT 148.755 -130.045 149.085 -129.715 ;
        RECT 148.755 -131.405 149.085 -131.075 ;
        RECT 148.755 -132.765 149.085 -132.435 ;
        RECT 148.755 -134.125 149.085 -133.795 ;
        RECT 148.755 -135.485 149.085 -135.155 ;
        RECT 148.755 -136.845 149.085 -136.515 ;
        RECT 148.755 -138.205 149.085 -137.875 ;
        RECT 148.755 -139.565 149.085 -139.235 ;
        RECT 148.755 -140.925 149.085 -140.595 ;
        RECT 148.755 -142.285 149.085 -141.955 ;
        RECT 148.755 -143.645 149.085 -143.315 ;
        RECT 148.755 -145.005 149.085 -144.675 ;
        RECT 148.755 -146.365 149.085 -146.035 ;
        RECT 148.755 -147.725 149.085 -147.395 ;
        RECT 148.755 -149.085 149.085 -148.755 ;
        RECT 148.755 -150.445 149.085 -150.115 ;
        RECT 148.755 -151.805 149.085 -151.475 ;
        RECT 148.755 -153.165 149.085 -152.835 ;
        RECT 148.755 -154.525 149.085 -154.195 ;
        RECT 148.755 -155.885 149.085 -155.555 ;
        RECT 148.755 -157.245 149.085 -156.915 ;
        RECT 148.755 -158.605 149.085 -158.275 ;
        RECT 148.755 -159.965 149.085 -159.635 ;
        RECT 148.755 -161.325 149.085 -160.995 ;
        RECT 148.755 -162.685 149.085 -162.355 ;
        RECT 148.755 -164.045 149.085 -163.715 ;
        RECT 148.755 -165.405 149.085 -165.075 ;
        RECT 148.755 -166.765 149.085 -166.435 ;
        RECT 148.755 -168.125 149.085 -167.795 ;
        RECT 148.755 -169.485 149.085 -169.155 ;
        RECT 148.755 -170.845 149.085 -170.515 ;
        RECT 148.755 -172.205 149.085 -171.875 ;
        RECT 148.755 -173.565 149.085 -173.235 ;
        RECT 148.755 -174.925 149.085 -174.595 ;
        RECT 148.755 -176.285 149.085 -175.955 ;
        RECT 148.755 -177.645 149.085 -177.315 ;
        RECT 148.755 -183.29 149.085 -182.16 ;
        RECT 148.76 -183.405 149.08 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 149.06 -94.075 149.39 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 150.115 244.04 150.445 245.17 ;
        RECT 150.115 239.875 150.445 240.205 ;
        RECT 150.115 238.515 150.445 238.845 ;
        RECT 150.115 237.155 150.445 237.485 ;
        RECT 150.12 237.155 150.44 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 151.475 244.04 151.805 245.17 ;
        RECT 151.475 239.875 151.805 240.205 ;
        RECT 151.475 238.515 151.805 238.845 ;
        RECT 151.475 237.155 151.805 237.485 ;
        RECT 151.48 237.155 151.8 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 151.475 -0.845 151.805 -0.515 ;
        RECT 151.475 -2.205 151.805 -1.875 ;
        RECT 151.475 -3.565 151.805 -3.235 ;
        RECT 151.48 -3.565 151.8 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 152.835 244.04 153.165 245.17 ;
        RECT 152.835 239.875 153.165 240.205 ;
        RECT 152.835 238.515 153.165 238.845 ;
        RECT 152.835 237.155 153.165 237.485 ;
        RECT 152.84 237.155 153.16 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 152.835 -0.845 153.165 -0.515 ;
        RECT 152.835 -2.205 153.165 -1.875 ;
        RECT 152.835 -3.565 153.165 -3.235 ;
        RECT 152.84 -3.565 153.16 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 154.195 244.04 154.525 245.17 ;
        RECT 154.195 239.875 154.525 240.205 ;
        RECT 154.195 238.515 154.525 238.845 ;
        RECT 154.195 237.155 154.525 237.485 ;
        RECT 154.2 237.155 154.52 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 154.195 -0.845 154.525 -0.515 ;
        RECT 154.195 -2.205 154.525 -1.875 ;
        RECT 154.195 -3.565 154.525 -3.235 ;
        RECT 154.2 -3.565 154.52 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 154.195 -91.965 154.525 -91.635 ;
        RECT 154.195 -93.325 154.525 -92.995 ;
        RECT 154.195 -94.685 154.525 -94.355 ;
        RECT 154.195 -96.045 154.525 -95.715 ;
        RECT 154.195 -97.405 154.525 -97.075 ;
        RECT 154.195 -98.765 154.525 -98.435 ;
        RECT 154.195 -100.125 154.525 -99.795 ;
        RECT 154.195 -101.485 154.525 -101.155 ;
        RECT 154.195 -102.845 154.525 -102.515 ;
        RECT 154.195 -104.205 154.525 -103.875 ;
        RECT 154.195 -105.565 154.525 -105.235 ;
        RECT 154.195 -106.925 154.525 -106.595 ;
        RECT 154.195 -108.285 154.525 -107.955 ;
        RECT 154.195 -109.645 154.525 -109.315 ;
        RECT 154.195 -111.005 154.525 -110.675 ;
        RECT 154.195 -112.365 154.525 -112.035 ;
        RECT 154.195 -113.725 154.525 -113.395 ;
        RECT 154.195 -115.085 154.525 -114.755 ;
        RECT 154.195 -116.445 154.525 -116.115 ;
        RECT 154.195 -117.805 154.525 -117.475 ;
        RECT 154.195 -119.165 154.525 -118.835 ;
        RECT 154.195 -120.525 154.525 -120.195 ;
        RECT 154.195 -121.885 154.525 -121.555 ;
        RECT 154.195 -123.245 154.525 -122.915 ;
        RECT 154.195 -124.605 154.525 -124.275 ;
        RECT 154.195 -125.965 154.525 -125.635 ;
        RECT 154.195 -127.325 154.525 -126.995 ;
        RECT 154.195 -128.685 154.525 -128.355 ;
        RECT 154.195 -130.045 154.525 -129.715 ;
        RECT 154.195 -131.405 154.525 -131.075 ;
        RECT 154.195 -132.765 154.525 -132.435 ;
        RECT 154.195 -134.125 154.525 -133.795 ;
        RECT 154.195 -135.485 154.525 -135.155 ;
        RECT 154.195 -136.845 154.525 -136.515 ;
        RECT 154.195 -138.205 154.525 -137.875 ;
        RECT 154.195 -139.565 154.525 -139.235 ;
        RECT 154.195 -140.925 154.525 -140.595 ;
        RECT 154.195 -142.285 154.525 -141.955 ;
        RECT 154.195 -143.645 154.525 -143.315 ;
        RECT 154.195 -145.005 154.525 -144.675 ;
        RECT 154.195 -146.365 154.525 -146.035 ;
        RECT 154.195 -147.725 154.525 -147.395 ;
        RECT 154.195 -149.085 154.525 -148.755 ;
        RECT 154.195 -150.445 154.525 -150.115 ;
        RECT 154.195 -151.805 154.525 -151.475 ;
        RECT 154.195 -153.165 154.525 -152.835 ;
        RECT 154.195 -154.525 154.525 -154.195 ;
        RECT 154.195 -155.885 154.525 -155.555 ;
        RECT 154.195 -157.245 154.525 -156.915 ;
        RECT 154.195 -158.605 154.525 -158.275 ;
        RECT 154.195 -159.965 154.525 -159.635 ;
        RECT 154.195 -161.325 154.525 -160.995 ;
        RECT 154.195 -162.685 154.525 -162.355 ;
        RECT 154.195 -164.045 154.525 -163.715 ;
        RECT 154.195 -165.405 154.525 -165.075 ;
        RECT 154.195 -166.765 154.525 -166.435 ;
        RECT 154.195 -168.125 154.525 -167.795 ;
        RECT 154.195 -169.485 154.525 -169.155 ;
        RECT 154.195 -170.845 154.525 -170.515 ;
        RECT 154.195 -172.205 154.525 -171.875 ;
        RECT 154.195 -173.565 154.525 -173.235 ;
        RECT 154.195 -174.925 154.525 -174.595 ;
        RECT 154.195 -176.285 154.525 -175.955 ;
        RECT 154.195 -177.645 154.525 -177.315 ;
        RECT 154.195 -183.29 154.525 -182.16 ;
        RECT 154.2 -183.405 154.52 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 155.16 -94.075 155.49 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 155.555 244.04 155.885 245.17 ;
        RECT 155.555 239.875 155.885 240.205 ;
        RECT 155.555 238.515 155.885 238.845 ;
        RECT 155.555 237.155 155.885 237.485 ;
        RECT 155.56 237.155 155.88 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 155.555 -96.045 155.885 -95.715 ;
        RECT 155.555 -97.405 155.885 -97.075 ;
        RECT 155.555 -98.765 155.885 -98.435 ;
        RECT 155.555 -100.125 155.885 -99.795 ;
        RECT 155.555 -101.485 155.885 -101.155 ;
        RECT 155.555 -102.845 155.885 -102.515 ;
        RECT 155.555 -104.205 155.885 -103.875 ;
        RECT 155.555 -105.565 155.885 -105.235 ;
        RECT 155.555 -106.925 155.885 -106.595 ;
        RECT 155.555 -108.285 155.885 -107.955 ;
        RECT 155.555 -109.645 155.885 -109.315 ;
        RECT 155.555 -111.005 155.885 -110.675 ;
        RECT 155.555 -112.365 155.885 -112.035 ;
        RECT 155.555 -113.725 155.885 -113.395 ;
        RECT 155.555 -115.085 155.885 -114.755 ;
        RECT 155.555 -116.445 155.885 -116.115 ;
        RECT 155.555 -117.805 155.885 -117.475 ;
        RECT 155.555 -119.165 155.885 -118.835 ;
        RECT 155.555 -120.525 155.885 -120.195 ;
        RECT 155.555 -121.885 155.885 -121.555 ;
        RECT 155.555 -123.245 155.885 -122.915 ;
        RECT 155.555 -124.605 155.885 -124.275 ;
        RECT 155.555 -125.965 155.885 -125.635 ;
        RECT 155.555 -127.325 155.885 -126.995 ;
        RECT 155.555 -128.685 155.885 -128.355 ;
        RECT 155.555 -130.045 155.885 -129.715 ;
        RECT 155.555 -131.405 155.885 -131.075 ;
        RECT 155.555 -132.765 155.885 -132.435 ;
        RECT 155.555 -134.125 155.885 -133.795 ;
        RECT 155.555 -135.485 155.885 -135.155 ;
        RECT 155.555 -136.845 155.885 -136.515 ;
        RECT 155.555 -138.205 155.885 -137.875 ;
        RECT 155.555 -139.565 155.885 -139.235 ;
        RECT 155.555 -140.925 155.885 -140.595 ;
        RECT 155.555 -142.285 155.885 -141.955 ;
        RECT 155.555 -143.645 155.885 -143.315 ;
        RECT 155.555 -145.005 155.885 -144.675 ;
        RECT 155.555 -146.365 155.885 -146.035 ;
        RECT 155.555 -147.725 155.885 -147.395 ;
        RECT 155.555 -149.085 155.885 -148.755 ;
        RECT 155.555 -150.445 155.885 -150.115 ;
        RECT 155.555 -151.805 155.885 -151.475 ;
        RECT 155.555 -153.165 155.885 -152.835 ;
        RECT 155.555 -154.525 155.885 -154.195 ;
        RECT 155.555 -155.885 155.885 -155.555 ;
        RECT 155.555 -157.245 155.885 -156.915 ;
        RECT 155.555 -158.605 155.885 -158.275 ;
        RECT 155.555 -159.965 155.885 -159.635 ;
        RECT 155.555 -161.325 155.885 -160.995 ;
        RECT 155.555 -162.685 155.885 -162.355 ;
        RECT 155.555 -164.045 155.885 -163.715 ;
        RECT 155.555 -165.405 155.885 -165.075 ;
        RECT 155.555 -166.765 155.885 -166.435 ;
        RECT 155.555 -168.125 155.885 -167.795 ;
        RECT 155.555 -169.485 155.885 -169.155 ;
        RECT 155.555 -170.845 155.885 -170.515 ;
        RECT 155.555 -172.205 155.885 -171.875 ;
        RECT 155.555 -173.565 155.885 -173.235 ;
        RECT 155.555 -174.925 155.885 -174.595 ;
        RECT 155.555 -176.285 155.885 -175.955 ;
        RECT 155.555 -177.645 155.885 -177.315 ;
        RECT 155.555 -183.29 155.885 -182.16 ;
        RECT 155.56 -183.405 155.88 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 156.915 244.04 157.245 245.17 ;
        RECT 156.915 239.875 157.245 240.205 ;
        RECT 156.915 238.515 157.245 238.845 ;
        RECT 156.915 237.155 157.245 237.485 ;
        RECT 156.92 237.155 157.24 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 156.915 -0.845 157.245 -0.515 ;
        RECT 156.915 -2.205 157.245 -1.875 ;
        RECT 156.915 -3.565 157.245 -3.235 ;
        RECT 156.92 -3.565 157.24 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 158.275 244.04 158.605 245.17 ;
        RECT 158.275 239.875 158.605 240.205 ;
        RECT 158.275 238.515 158.605 238.845 ;
        RECT 158.275 237.155 158.605 237.485 ;
        RECT 158.28 237.155 158.6 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 158.275 -0.845 158.605 -0.515 ;
        RECT 158.275 -2.205 158.605 -1.875 ;
        RECT 158.275 -3.565 158.605 -3.235 ;
        RECT 158.28 -3.565 158.6 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 159.635 244.04 159.965 245.17 ;
        RECT 159.635 239.875 159.965 240.205 ;
        RECT 159.635 238.515 159.965 238.845 ;
        RECT 159.635 237.155 159.965 237.485 ;
        RECT 159.64 237.155 159.96 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 159.635 -0.845 159.965 -0.515 ;
        RECT 159.635 -2.205 159.965 -1.875 ;
        RECT 159.635 -3.565 159.965 -3.235 ;
        RECT 159.64 -3.565 159.96 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 159.635 -91.965 159.965 -91.635 ;
        RECT 159.635 -93.325 159.965 -92.995 ;
        RECT 159.635 -94.685 159.965 -94.355 ;
        RECT 159.635 -96.045 159.965 -95.715 ;
        RECT 159.635 -97.405 159.965 -97.075 ;
        RECT 159.635 -98.765 159.965 -98.435 ;
        RECT 159.635 -100.125 159.965 -99.795 ;
        RECT 159.635 -101.485 159.965 -101.155 ;
        RECT 159.635 -102.845 159.965 -102.515 ;
        RECT 159.635 -104.205 159.965 -103.875 ;
        RECT 159.635 -105.565 159.965 -105.235 ;
        RECT 159.635 -106.925 159.965 -106.595 ;
        RECT 159.635 -108.285 159.965 -107.955 ;
        RECT 159.635 -109.645 159.965 -109.315 ;
        RECT 159.635 -111.005 159.965 -110.675 ;
        RECT 159.635 -112.365 159.965 -112.035 ;
        RECT 159.635 -113.725 159.965 -113.395 ;
        RECT 159.635 -115.085 159.965 -114.755 ;
        RECT 159.635 -116.445 159.965 -116.115 ;
        RECT 159.635 -117.805 159.965 -117.475 ;
        RECT 159.635 -119.165 159.965 -118.835 ;
        RECT 159.635 -120.525 159.965 -120.195 ;
        RECT 159.635 -121.885 159.965 -121.555 ;
        RECT 159.635 -123.245 159.965 -122.915 ;
        RECT 159.635 -124.605 159.965 -124.275 ;
        RECT 159.635 -125.965 159.965 -125.635 ;
        RECT 159.635 -127.325 159.965 -126.995 ;
        RECT 159.635 -128.685 159.965 -128.355 ;
        RECT 159.635 -130.045 159.965 -129.715 ;
        RECT 159.635 -131.405 159.965 -131.075 ;
        RECT 159.635 -132.765 159.965 -132.435 ;
        RECT 159.635 -134.125 159.965 -133.795 ;
        RECT 159.635 -135.485 159.965 -135.155 ;
        RECT 159.635 -136.845 159.965 -136.515 ;
        RECT 159.635 -138.205 159.965 -137.875 ;
        RECT 159.635 -139.565 159.965 -139.235 ;
        RECT 159.635 -140.925 159.965 -140.595 ;
        RECT 159.635 -142.285 159.965 -141.955 ;
        RECT 159.635 -143.645 159.965 -143.315 ;
        RECT 159.635 -145.005 159.965 -144.675 ;
        RECT 159.635 -146.365 159.965 -146.035 ;
        RECT 159.635 -147.725 159.965 -147.395 ;
        RECT 159.635 -149.085 159.965 -148.755 ;
        RECT 159.635 -150.445 159.965 -150.115 ;
        RECT 159.635 -151.805 159.965 -151.475 ;
        RECT 159.635 -153.165 159.965 -152.835 ;
        RECT 159.635 -154.525 159.965 -154.195 ;
        RECT 159.635 -155.885 159.965 -155.555 ;
        RECT 159.635 -157.245 159.965 -156.915 ;
        RECT 159.635 -158.605 159.965 -158.275 ;
        RECT 159.635 -159.965 159.965 -159.635 ;
        RECT 159.635 -161.325 159.965 -160.995 ;
        RECT 159.635 -162.685 159.965 -162.355 ;
        RECT 159.635 -164.045 159.965 -163.715 ;
        RECT 159.635 -165.405 159.965 -165.075 ;
        RECT 159.635 -166.765 159.965 -166.435 ;
        RECT 159.635 -168.125 159.965 -167.795 ;
        RECT 159.635 -169.485 159.965 -169.155 ;
        RECT 159.635 -170.845 159.965 -170.515 ;
        RECT 159.635 -172.205 159.965 -171.875 ;
        RECT 159.635 -173.565 159.965 -173.235 ;
        RECT 159.635 -174.925 159.965 -174.595 ;
        RECT 159.635 -176.285 159.965 -175.955 ;
        RECT 159.635 -177.645 159.965 -177.315 ;
        RECT 159.635 -183.29 159.965 -182.16 ;
        RECT 159.64 -183.405 159.96 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 160.995 244.04 161.325 245.17 ;
        RECT 160.995 239.875 161.325 240.205 ;
        RECT 160.995 238.515 161.325 238.845 ;
        RECT 160.995 237.155 161.325 237.485 ;
        RECT 161 237.155 161.32 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 160.995 -96.045 161.325 -95.715 ;
        RECT 160.995 -97.405 161.325 -97.075 ;
        RECT 160.995 -98.765 161.325 -98.435 ;
        RECT 160.995 -100.125 161.325 -99.795 ;
        RECT 160.995 -101.485 161.325 -101.155 ;
        RECT 160.995 -102.845 161.325 -102.515 ;
        RECT 160.995 -104.205 161.325 -103.875 ;
        RECT 160.995 -105.565 161.325 -105.235 ;
        RECT 160.995 -106.925 161.325 -106.595 ;
        RECT 160.995 -108.285 161.325 -107.955 ;
        RECT 160.995 -109.645 161.325 -109.315 ;
        RECT 160.995 -111.005 161.325 -110.675 ;
        RECT 160.995 -112.365 161.325 -112.035 ;
        RECT 160.995 -113.725 161.325 -113.395 ;
        RECT 160.995 -115.085 161.325 -114.755 ;
        RECT 160.995 -116.445 161.325 -116.115 ;
        RECT 160.995 -117.805 161.325 -117.475 ;
        RECT 160.995 -119.165 161.325 -118.835 ;
        RECT 160.995 -120.525 161.325 -120.195 ;
        RECT 160.995 -121.885 161.325 -121.555 ;
        RECT 160.995 -123.245 161.325 -122.915 ;
        RECT 160.995 -124.605 161.325 -124.275 ;
        RECT 160.995 -125.965 161.325 -125.635 ;
        RECT 160.995 -127.325 161.325 -126.995 ;
        RECT 160.995 -128.685 161.325 -128.355 ;
        RECT 160.995 -130.045 161.325 -129.715 ;
        RECT 160.995 -131.405 161.325 -131.075 ;
        RECT 160.995 -132.765 161.325 -132.435 ;
        RECT 160.995 -134.125 161.325 -133.795 ;
        RECT 160.995 -135.485 161.325 -135.155 ;
        RECT 160.995 -136.845 161.325 -136.515 ;
        RECT 160.995 -138.205 161.325 -137.875 ;
        RECT 160.995 -139.565 161.325 -139.235 ;
        RECT 160.995 -140.925 161.325 -140.595 ;
        RECT 160.995 -142.285 161.325 -141.955 ;
        RECT 160.995 -143.645 161.325 -143.315 ;
        RECT 160.995 -145.005 161.325 -144.675 ;
        RECT 160.995 -146.365 161.325 -146.035 ;
        RECT 160.995 -147.725 161.325 -147.395 ;
        RECT 160.995 -149.085 161.325 -148.755 ;
        RECT 160.995 -150.445 161.325 -150.115 ;
        RECT 160.995 -151.805 161.325 -151.475 ;
        RECT 160.995 -153.165 161.325 -152.835 ;
        RECT 160.995 -154.525 161.325 -154.195 ;
        RECT 160.995 -155.885 161.325 -155.555 ;
        RECT 160.995 -157.245 161.325 -156.915 ;
        RECT 160.995 -158.605 161.325 -158.275 ;
        RECT 160.995 -159.965 161.325 -159.635 ;
        RECT 160.995 -161.325 161.325 -160.995 ;
        RECT 160.995 -162.685 161.325 -162.355 ;
        RECT 160.995 -164.045 161.325 -163.715 ;
        RECT 160.995 -165.405 161.325 -165.075 ;
        RECT 160.995 -166.765 161.325 -166.435 ;
        RECT 160.995 -168.125 161.325 -167.795 ;
        RECT 160.995 -169.485 161.325 -169.155 ;
        RECT 160.995 -170.845 161.325 -170.515 ;
        RECT 160.995 -172.205 161.325 -171.875 ;
        RECT 160.995 -173.565 161.325 -173.235 ;
        RECT 160.995 -174.925 161.325 -174.595 ;
        RECT 160.995 -176.285 161.325 -175.955 ;
        RECT 160.995 -177.645 161.325 -177.315 ;
        RECT 160.995 -183.29 161.325 -182.16 ;
        RECT 161 -183.405 161.32 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 161.26 -94.075 161.59 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 162.355 244.04 162.685 245.17 ;
        RECT 162.355 239.875 162.685 240.205 ;
        RECT 162.355 238.515 162.685 238.845 ;
        RECT 162.355 237.155 162.685 237.485 ;
        RECT 162.36 237.155 162.68 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 163.715 244.04 164.045 245.17 ;
        RECT 163.715 239.875 164.045 240.205 ;
        RECT 163.715 238.515 164.045 238.845 ;
        RECT 163.715 237.155 164.045 237.485 ;
        RECT 163.72 237.155 164.04 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 163.715 -0.845 164.045 -0.515 ;
        RECT 163.715 -2.205 164.045 -1.875 ;
        RECT 163.715 -3.565 164.045 -3.235 ;
        RECT 163.72 -3.565 164.04 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 165.075 244.04 165.405 245.17 ;
        RECT 165.075 239.875 165.405 240.205 ;
        RECT 165.075 238.515 165.405 238.845 ;
        RECT 165.075 237.155 165.405 237.485 ;
        RECT 165.08 237.155 165.4 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 165.075 -0.845 165.405 -0.515 ;
        RECT 165.075 -2.205 165.405 -1.875 ;
        RECT 165.075 -3.565 165.405 -3.235 ;
        RECT 165.08 -3.565 165.4 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 165.075 -91.965 165.405 -91.635 ;
        RECT 165.075 -93.325 165.405 -92.995 ;
        RECT 165.075 -94.685 165.405 -94.355 ;
        RECT 165.075 -96.045 165.405 -95.715 ;
        RECT 165.075 -97.405 165.405 -97.075 ;
        RECT 165.075 -98.765 165.405 -98.435 ;
        RECT 165.075 -100.125 165.405 -99.795 ;
        RECT 165.075 -101.485 165.405 -101.155 ;
        RECT 165.075 -102.845 165.405 -102.515 ;
        RECT 165.075 -104.205 165.405 -103.875 ;
        RECT 165.075 -105.565 165.405 -105.235 ;
        RECT 165.075 -106.925 165.405 -106.595 ;
        RECT 165.075 -108.285 165.405 -107.955 ;
        RECT 165.075 -109.645 165.405 -109.315 ;
        RECT 165.075 -111.005 165.405 -110.675 ;
        RECT 165.075 -112.365 165.405 -112.035 ;
        RECT 165.075 -113.725 165.405 -113.395 ;
        RECT 165.075 -115.085 165.405 -114.755 ;
        RECT 165.075 -116.445 165.405 -116.115 ;
        RECT 165.075 -117.805 165.405 -117.475 ;
        RECT 165.075 -119.165 165.405 -118.835 ;
        RECT 165.075 -120.525 165.405 -120.195 ;
        RECT 165.075 -121.885 165.405 -121.555 ;
        RECT 165.075 -123.245 165.405 -122.915 ;
        RECT 165.075 -124.605 165.405 -124.275 ;
        RECT 165.075 -125.965 165.405 -125.635 ;
        RECT 165.075 -127.325 165.405 -126.995 ;
        RECT 165.075 -128.685 165.405 -128.355 ;
        RECT 165.075 -130.045 165.405 -129.715 ;
        RECT 165.075 -131.405 165.405 -131.075 ;
        RECT 165.075 -132.765 165.405 -132.435 ;
        RECT 165.075 -134.125 165.405 -133.795 ;
        RECT 165.075 -135.485 165.405 -135.155 ;
        RECT 165.075 -136.845 165.405 -136.515 ;
        RECT 165.075 -138.205 165.405 -137.875 ;
        RECT 165.075 -139.565 165.405 -139.235 ;
        RECT 165.075 -140.925 165.405 -140.595 ;
        RECT 165.075 -142.285 165.405 -141.955 ;
        RECT 165.075 -143.645 165.405 -143.315 ;
        RECT 165.075 -145.005 165.405 -144.675 ;
        RECT 165.075 -146.365 165.405 -146.035 ;
        RECT 165.075 -147.725 165.405 -147.395 ;
        RECT 165.075 -149.085 165.405 -148.755 ;
        RECT 165.075 -150.445 165.405 -150.115 ;
        RECT 165.075 -151.805 165.405 -151.475 ;
        RECT 165.075 -153.165 165.405 -152.835 ;
        RECT 165.075 -154.525 165.405 -154.195 ;
        RECT 165.075 -155.885 165.405 -155.555 ;
        RECT 165.075 -157.245 165.405 -156.915 ;
        RECT 165.075 -158.605 165.405 -158.275 ;
        RECT 165.075 -159.965 165.405 -159.635 ;
        RECT 165.075 -161.325 165.405 -160.995 ;
        RECT 165.075 -162.685 165.405 -162.355 ;
        RECT 165.075 -164.045 165.405 -163.715 ;
        RECT 165.075 -165.405 165.405 -165.075 ;
        RECT 165.075 -166.765 165.405 -166.435 ;
        RECT 165.075 -168.125 165.405 -167.795 ;
        RECT 165.075 -169.485 165.405 -169.155 ;
        RECT 165.075 -170.845 165.405 -170.515 ;
        RECT 165.075 -172.205 165.405 -171.875 ;
        RECT 165.075 -173.565 165.405 -173.235 ;
        RECT 165.075 -174.925 165.405 -174.595 ;
        RECT 165.075 -176.285 165.405 -175.955 ;
        RECT 165.075 -177.645 165.405 -177.315 ;
        RECT 165.075 -183.29 165.405 -182.16 ;
        RECT 165.08 -183.405 165.4 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 166.435 244.04 166.765 245.17 ;
        RECT 166.435 239.875 166.765 240.205 ;
        RECT 166.435 238.515 166.765 238.845 ;
        RECT 166.435 237.155 166.765 237.485 ;
        RECT 166.44 237.155 166.76 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 166.435 -0.845 166.765 -0.515 ;
        RECT 166.435 -2.205 166.765 -1.875 ;
        RECT 166.435 -3.565 166.765 -3.235 ;
        RECT 166.44 -3.565 166.76 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 166.435 -91.965 166.765 -91.635 ;
        RECT 166.435 -93.325 166.765 -92.995 ;
        RECT 166.435 -94.685 166.765 -94.355 ;
        RECT 166.435 -96.045 166.765 -95.715 ;
        RECT 166.435 -97.405 166.765 -97.075 ;
        RECT 166.435 -98.765 166.765 -98.435 ;
        RECT 166.435 -100.125 166.765 -99.795 ;
        RECT 166.435 -101.485 166.765 -101.155 ;
        RECT 166.435 -102.845 166.765 -102.515 ;
        RECT 166.435 -104.205 166.765 -103.875 ;
        RECT 166.435 -105.565 166.765 -105.235 ;
        RECT 166.435 -106.925 166.765 -106.595 ;
        RECT 166.435 -108.285 166.765 -107.955 ;
        RECT 166.435 -109.645 166.765 -109.315 ;
        RECT 166.435 -111.005 166.765 -110.675 ;
        RECT 166.435 -112.365 166.765 -112.035 ;
        RECT 166.435 -113.725 166.765 -113.395 ;
        RECT 166.435 -115.085 166.765 -114.755 ;
        RECT 166.435 -116.445 166.765 -116.115 ;
        RECT 166.435 -117.805 166.765 -117.475 ;
        RECT 166.435 -119.165 166.765 -118.835 ;
        RECT 166.435 -120.525 166.765 -120.195 ;
        RECT 166.435 -121.885 166.765 -121.555 ;
        RECT 166.435 -123.245 166.765 -122.915 ;
        RECT 166.435 -124.605 166.765 -124.275 ;
        RECT 166.435 -125.965 166.765 -125.635 ;
        RECT 166.435 -127.325 166.765 -126.995 ;
        RECT 166.435 -128.685 166.765 -128.355 ;
        RECT 166.435 -130.045 166.765 -129.715 ;
        RECT 166.435 -131.405 166.765 -131.075 ;
        RECT 166.435 -132.765 166.765 -132.435 ;
        RECT 166.435 -134.125 166.765 -133.795 ;
        RECT 166.435 -135.485 166.765 -135.155 ;
        RECT 166.435 -136.845 166.765 -136.515 ;
        RECT 166.435 -138.205 166.765 -137.875 ;
        RECT 166.435 -139.565 166.765 -139.235 ;
        RECT 166.435 -140.925 166.765 -140.595 ;
        RECT 166.435 -142.285 166.765 -141.955 ;
        RECT 166.435 -143.645 166.765 -143.315 ;
        RECT 166.435 -145.005 166.765 -144.675 ;
        RECT 166.435 -146.365 166.765 -146.035 ;
        RECT 166.435 -147.725 166.765 -147.395 ;
        RECT 166.435 -149.085 166.765 -148.755 ;
        RECT 166.435 -150.445 166.765 -150.115 ;
        RECT 166.435 -151.805 166.765 -151.475 ;
        RECT 166.435 -153.165 166.765 -152.835 ;
        RECT 166.435 -154.525 166.765 -154.195 ;
        RECT 166.435 -155.885 166.765 -155.555 ;
        RECT 166.435 -157.245 166.765 -156.915 ;
        RECT 166.435 -158.605 166.765 -158.275 ;
        RECT 166.435 -159.965 166.765 -159.635 ;
        RECT 166.435 -161.325 166.765 -160.995 ;
        RECT 166.435 -162.685 166.765 -162.355 ;
        RECT 166.435 -164.045 166.765 -163.715 ;
        RECT 166.435 -165.405 166.765 -165.075 ;
        RECT 166.435 -166.765 166.765 -166.435 ;
        RECT 166.435 -168.125 166.765 -167.795 ;
        RECT 166.435 -169.485 166.765 -169.155 ;
        RECT 166.435 -170.845 166.765 -170.515 ;
        RECT 166.435 -172.205 166.765 -171.875 ;
        RECT 166.435 -173.565 166.765 -173.235 ;
        RECT 166.435 -174.925 166.765 -174.595 ;
        RECT 166.435 -176.285 166.765 -175.955 ;
        RECT 166.435 -177.645 166.765 -177.315 ;
        RECT 166.435 -183.29 166.765 -182.16 ;
        RECT 166.44 -183.405 166.76 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 167.36 -94.075 167.69 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 167.795 244.04 168.125 245.17 ;
        RECT 167.795 239.875 168.125 240.205 ;
        RECT 167.795 238.515 168.125 238.845 ;
        RECT 167.795 237.155 168.125 237.485 ;
        RECT 167.8 237.155 168.12 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 167.795 -96.045 168.125 -95.715 ;
        RECT 167.795 -97.405 168.125 -97.075 ;
        RECT 167.795 -98.765 168.125 -98.435 ;
        RECT 167.795 -100.125 168.125 -99.795 ;
        RECT 167.795 -101.485 168.125 -101.155 ;
        RECT 167.795 -102.845 168.125 -102.515 ;
        RECT 167.795 -104.205 168.125 -103.875 ;
        RECT 167.795 -105.565 168.125 -105.235 ;
        RECT 167.795 -106.925 168.125 -106.595 ;
        RECT 167.795 -108.285 168.125 -107.955 ;
        RECT 167.795 -109.645 168.125 -109.315 ;
        RECT 167.795 -111.005 168.125 -110.675 ;
        RECT 167.795 -112.365 168.125 -112.035 ;
        RECT 167.795 -113.725 168.125 -113.395 ;
        RECT 167.795 -115.085 168.125 -114.755 ;
        RECT 167.795 -116.445 168.125 -116.115 ;
        RECT 167.795 -117.805 168.125 -117.475 ;
        RECT 167.795 -119.165 168.125 -118.835 ;
        RECT 167.795 -120.525 168.125 -120.195 ;
        RECT 167.795 -121.885 168.125 -121.555 ;
        RECT 167.795 -123.245 168.125 -122.915 ;
        RECT 167.795 -124.605 168.125 -124.275 ;
        RECT 167.795 -125.965 168.125 -125.635 ;
        RECT 167.795 -127.325 168.125 -126.995 ;
        RECT 167.795 -128.685 168.125 -128.355 ;
        RECT 167.795 -130.045 168.125 -129.715 ;
        RECT 167.795 -131.405 168.125 -131.075 ;
        RECT 167.795 -132.765 168.125 -132.435 ;
        RECT 167.795 -134.125 168.125 -133.795 ;
        RECT 167.795 -135.485 168.125 -135.155 ;
        RECT 167.795 -136.845 168.125 -136.515 ;
        RECT 167.795 -138.205 168.125 -137.875 ;
        RECT 167.795 -139.565 168.125 -139.235 ;
        RECT 167.795 -140.925 168.125 -140.595 ;
        RECT 167.795 -142.285 168.125 -141.955 ;
        RECT 167.795 -143.645 168.125 -143.315 ;
        RECT 167.795 -145.005 168.125 -144.675 ;
        RECT 167.795 -146.365 168.125 -146.035 ;
        RECT 167.795 -147.725 168.125 -147.395 ;
        RECT 167.795 -149.085 168.125 -148.755 ;
        RECT 167.795 -150.445 168.125 -150.115 ;
        RECT 167.795 -151.805 168.125 -151.475 ;
        RECT 167.795 -153.165 168.125 -152.835 ;
        RECT 167.795 -154.525 168.125 -154.195 ;
        RECT 167.795 -155.885 168.125 -155.555 ;
        RECT 167.795 -157.245 168.125 -156.915 ;
        RECT 167.795 -158.605 168.125 -158.275 ;
        RECT 167.795 -159.965 168.125 -159.635 ;
        RECT 167.795 -161.325 168.125 -160.995 ;
        RECT 167.795 -162.685 168.125 -162.355 ;
        RECT 167.795 -164.045 168.125 -163.715 ;
        RECT 167.795 -165.405 168.125 -165.075 ;
        RECT 167.795 -166.765 168.125 -166.435 ;
        RECT 167.795 -168.125 168.125 -167.795 ;
        RECT 167.795 -169.485 168.125 -169.155 ;
        RECT 167.795 -170.845 168.125 -170.515 ;
        RECT 167.795 -172.205 168.125 -171.875 ;
        RECT 167.795 -173.565 168.125 -173.235 ;
        RECT 167.795 -174.925 168.125 -174.595 ;
        RECT 167.795 -176.285 168.125 -175.955 ;
        RECT 167.795 -177.645 168.125 -177.315 ;
        RECT 167.795 -183.29 168.125 -182.16 ;
        RECT 167.8 -183.405 168.12 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 169.155 244.04 169.485 245.17 ;
        RECT 169.155 239.875 169.485 240.205 ;
        RECT 169.155 238.515 169.485 238.845 ;
        RECT 169.155 237.155 169.485 237.485 ;
        RECT 169.16 237.155 169.48 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 169.155 -0.845 169.485 -0.515 ;
        RECT 169.155 -2.205 169.485 -1.875 ;
        RECT 169.155 -3.565 169.485 -3.235 ;
        RECT 169.16 -3.565 169.48 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 170.515 244.04 170.845 245.17 ;
        RECT 170.515 239.875 170.845 240.205 ;
        RECT 170.515 238.515 170.845 238.845 ;
        RECT 170.515 237.155 170.845 237.485 ;
        RECT 170.52 237.155 170.84 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 170.515 -0.845 170.845 -0.515 ;
        RECT 170.515 -2.205 170.845 -1.875 ;
        RECT 170.515 -3.565 170.845 -3.235 ;
        RECT 170.52 -3.565 170.84 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 171.875 244.04 172.205 245.17 ;
        RECT 171.875 239.875 172.205 240.205 ;
        RECT 171.875 238.515 172.205 238.845 ;
        RECT 171.875 237.155 172.205 237.485 ;
        RECT 171.88 237.155 172.2 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 171.875 -0.845 172.205 -0.515 ;
        RECT 171.875 -2.205 172.205 -1.875 ;
        RECT 171.875 -3.565 172.205 -3.235 ;
        RECT 171.88 -3.565 172.2 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 171.875 -157.245 172.205 -156.915 ;
        RECT 171.875 -158.605 172.205 -158.275 ;
        RECT 171.875 -159.965 172.205 -159.635 ;
        RECT 171.875 -161.325 172.205 -160.995 ;
        RECT 171.875 -162.685 172.205 -162.355 ;
        RECT 171.875 -164.045 172.205 -163.715 ;
        RECT 171.875 -165.405 172.205 -165.075 ;
        RECT 171.875 -166.765 172.205 -166.435 ;
        RECT 171.875 -168.125 172.205 -167.795 ;
        RECT 171.875 -169.485 172.205 -169.155 ;
        RECT 171.875 -170.845 172.205 -170.515 ;
        RECT 171.875 -172.205 172.205 -171.875 ;
        RECT 171.875 -173.565 172.205 -173.235 ;
        RECT 171.875 -174.925 172.205 -174.595 ;
        RECT 171.875 -176.285 172.205 -175.955 ;
        RECT 171.875 -177.645 172.205 -177.315 ;
        RECT 171.875 -183.29 172.205 -182.16 ;
        RECT 171.88 -183.405 172.2 -90.96 ;
        RECT 171.875 -91.965 172.205 -91.635 ;
        RECT 171.875 -93.325 172.205 -92.995 ;
        RECT 171.875 -94.685 172.205 -94.355 ;
        RECT 171.875 -96.045 172.205 -95.715 ;
        RECT 171.875 -97.405 172.205 -97.075 ;
        RECT 171.875 -98.765 172.205 -98.435 ;
        RECT 171.875 -100.125 172.205 -99.795 ;
        RECT 171.875 -101.485 172.205 -101.155 ;
        RECT 171.875 -102.845 172.205 -102.515 ;
        RECT 171.875 -104.205 172.205 -103.875 ;
        RECT 171.875 -105.565 172.205 -105.235 ;
        RECT 171.875 -106.925 172.205 -106.595 ;
        RECT 171.875 -108.285 172.205 -107.955 ;
        RECT 171.875 -109.645 172.205 -109.315 ;
        RECT 171.875 -111.005 172.205 -110.675 ;
        RECT 171.875 -112.365 172.205 -112.035 ;
        RECT 171.875 -113.725 172.205 -113.395 ;
        RECT 171.875 -115.085 172.205 -114.755 ;
        RECT 171.875 -116.445 172.205 -116.115 ;
        RECT 171.875 -117.805 172.205 -117.475 ;
        RECT 171.875 -119.165 172.205 -118.835 ;
        RECT 171.875 -120.525 172.205 -120.195 ;
        RECT 171.875 -121.885 172.205 -121.555 ;
        RECT 171.875 -123.245 172.205 -122.915 ;
        RECT 171.875 -124.605 172.205 -124.275 ;
        RECT 171.875 -125.965 172.205 -125.635 ;
        RECT 171.875 -127.325 172.205 -126.995 ;
        RECT 171.875 -128.685 172.205 -128.355 ;
        RECT 171.875 -130.045 172.205 -129.715 ;
        RECT 171.875 -131.405 172.205 -131.075 ;
        RECT 171.875 -132.765 172.205 -132.435 ;
        RECT 171.875 -134.125 172.205 -133.795 ;
        RECT 171.875 -135.485 172.205 -135.155 ;
        RECT 171.875 -136.845 172.205 -136.515 ;
        RECT 171.875 -138.205 172.205 -137.875 ;
        RECT 171.875 -139.565 172.205 -139.235 ;
        RECT 171.875 -140.925 172.205 -140.595 ;
        RECT 171.875 -142.285 172.205 -141.955 ;
        RECT 171.875 -143.645 172.205 -143.315 ;
        RECT 171.875 -145.005 172.205 -144.675 ;
        RECT 171.875 -146.365 172.205 -146.035 ;
        RECT 171.875 -147.725 172.205 -147.395 ;
        RECT 171.875 -149.085 172.205 -148.755 ;
        RECT 171.875 -150.445 172.205 -150.115 ;
        RECT 171.875 -151.805 172.205 -151.475 ;
        RECT 171.875 -153.165 172.205 -152.835 ;
        RECT 171.875 -154.525 172.205 -154.195 ;
        RECT 171.875 -155.885 172.205 -155.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 106.36 -94.075 106.69 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 106.595 244.04 106.925 245.17 ;
        RECT 106.595 239.875 106.925 240.205 ;
        RECT 106.595 238.515 106.925 238.845 ;
        RECT 106.595 237.155 106.925 237.485 ;
        RECT 106.6 237.155 106.92 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 106.595 -96.045 106.925 -95.715 ;
        RECT 106.595 -97.405 106.925 -97.075 ;
        RECT 106.595 -98.765 106.925 -98.435 ;
        RECT 106.595 -100.125 106.925 -99.795 ;
        RECT 106.595 -101.485 106.925 -101.155 ;
        RECT 106.595 -102.845 106.925 -102.515 ;
        RECT 106.595 -104.205 106.925 -103.875 ;
        RECT 106.595 -105.565 106.925 -105.235 ;
        RECT 106.595 -106.925 106.925 -106.595 ;
        RECT 106.595 -108.285 106.925 -107.955 ;
        RECT 106.595 -109.645 106.925 -109.315 ;
        RECT 106.595 -111.005 106.925 -110.675 ;
        RECT 106.595 -112.365 106.925 -112.035 ;
        RECT 106.595 -113.725 106.925 -113.395 ;
        RECT 106.595 -115.085 106.925 -114.755 ;
        RECT 106.595 -116.445 106.925 -116.115 ;
        RECT 106.595 -117.805 106.925 -117.475 ;
        RECT 106.595 -119.165 106.925 -118.835 ;
        RECT 106.595 -120.525 106.925 -120.195 ;
        RECT 106.595 -121.885 106.925 -121.555 ;
        RECT 106.595 -123.245 106.925 -122.915 ;
        RECT 106.595 -124.605 106.925 -124.275 ;
        RECT 106.595 -125.965 106.925 -125.635 ;
        RECT 106.595 -127.325 106.925 -126.995 ;
        RECT 106.595 -128.685 106.925 -128.355 ;
        RECT 106.595 -130.045 106.925 -129.715 ;
        RECT 106.595 -131.405 106.925 -131.075 ;
        RECT 106.595 -132.765 106.925 -132.435 ;
        RECT 106.595 -134.125 106.925 -133.795 ;
        RECT 106.595 -135.485 106.925 -135.155 ;
        RECT 106.595 -136.845 106.925 -136.515 ;
        RECT 106.595 -138.205 106.925 -137.875 ;
        RECT 106.595 -139.565 106.925 -139.235 ;
        RECT 106.595 -140.925 106.925 -140.595 ;
        RECT 106.595 -142.285 106.925 -141.955 ;
        RECT 106.595 -143.645 106.925 -143.315 ;
        RECT 106.595 -145.005 106.925 -144.675 ;
        RECT 106.595 -146.365 106.925 -146.035 ;
        RECT 106.595 -147.725 106.925 -147.395 ;
        RECT 106.595 -149.085 106.925 -148.755 ;
        RECT 106.595 -150.445 106.925 -150.115 ;
        RECT 106.595 -151.805 106.925 -151.475 ;
        RECT 106.595 -153.165 106.925 -152.835 ;
        RECT 106.595 -154.525 106.925 -154.195 ;
        RECT 106.595 -155.885 106.925 -155.555 ;
        RECT 106.595 -157.245 106.925 -156.915 ;
        RECT 106.595 -158.605 106.925 -158.275 ;
        RECT 106.595 -159.965 106.925 -159.635 ;
        RECT 106.595 -161.325 106.925 -160.995 ;
        RECT 106.595 -162.685 106.925 -162.355 ;
        RECT 106.595 -164.045 106.925 -163.715 ;
        RECT 106.595 -165.405 106.925 -165.075 ;
        RECT 106.595 -166.765 106.925 -166.435 ;
        RECT 106.595 -168.125 106.925 -167.795 ;
        RECT 106.595 -169.485 106.925 -169.155 ;
        RECT 106.595 -170.845 106.925 -170.515 ;
        RECT 106.595 -172.205 106.925 -171.875 ;
        RECT 106.595 -173.565 106.925 -173.235 ;
        RECT 106.595 -174.925 106.925 -174.595 ;
        RECT 106.595 -176.285 106.925 -175.955 ;
        RECT 106.595 -177.645 106.925 -177.315 ;
        RECT 106.595 -183.29 106.925 -182.16 ;
        RECT 106.6 -183.405 106.92 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 107.955 244.04 108.285 245.17 ;
        RECT 107.955 239.875 108.285 240.205 ;
        RECT 107.955 238.515 108.285 238.845 ;
        RECT 107.955 237.155 108.285 237.485 ;
        RECT 107.96 237.155 108.28 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 107.955 -0.845 108.285 -0.515 ;
        RECT 107.955 -2.205 108.285 -1.875 ;
        RECT 107.955 -3.565 108.285 -3.235 ;
        RECT 107.96 -3.565 108.28 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 109.315 244.04 109.645 245.17 ;
        RECT 109.315 239.875 109.645 240.205 ;
        RECT 109.315 238.515 109.645 238.845 ;
        RECT 109.315 237.155 109.645 237.485 ;
        RECT 109.32 237.155 109.64 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 109.315 -0.845 109.645 -0.515 ;
        RECT 109.315 -2.205 109.645 -1.875 ;
        RECT 109.315 -3.565 109.645 -3.235 ;
        RECT 109.32 -3.565 109.64 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 110.675 244.04 111.005 245.17 ;
        RECT 110.675 239.875 111.005 240.205 ;
        RECT 110.675 238.515 111.005 238.845 ;
        RECT 110.675 237.155 111.005 237.485 ;
        RECT 110.68 237.155 111 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 110.675 -0.845 111.005 -0.515 ;
        RECT 110.675 -2.205 111.005 -1.875 ;
        RECT 110.675 -3.565 111.005 -3.235 ;
        RECT 110.68 -3.565 111 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 110.675 -91.965 111.005 -91.635 ;
        RECT 110.675 -93.325 111.005 -92.995 ;
        RECT 110.675 -94.685 111.005 -94.355 ;
        RECT 110.675 -96.045 111.005 -95.715 ;
        RECT 110.675 -97.405 111.005 -97.075 ;
        RECT 110.675 -98.765 111.005 -98.435 ;
        RECT 110.675 -100.125 111.005 -99.795 ;
        RECT 110.675 -101.485 111.005 -101.155 ;
        RECT 110.675 -102.845 111.005 -102.515 ;
        RECT 110.675 -104.205 111.005 -103.875 ;
        RECT 110.675 -105.565 111.005 -105.235 ;
        RECT 110.675 -106.925 111.005 -106.595 ;
        RECT 110.675 -108.285 111.005 -107.955 ;
        RECT 110.675 -109.645 111.005 -109.315 ;
        RECT 110.675 -111.005 111.005 -110.675 ;
        RECT 110.675 -112.365 111.005 -112.035 ;
        RECT 110.675 -113.725 111.005 -113.395 ;
        RECT 110.675 -115.085 111.005 -114.755 ;
        RECT 110.675 -116.445 111.005 -116.115 ;
        RECT 110.675 -117.805 111.005 -117.475 ;
        RECT 110.675 -119.165 111.005 -118.835 ;
        RECT 110.675 -120.525 111.005 -120.195 ;
        RECT 110.675 -121.885 111.005 -121.555 ;
        RECT 110.675 -123.245 111.005 -122.915 ;
        RECT 110.675 -124.605 111.005 -124.275 ;
        RECT 110.675 -125.965 111.005 -125.635 ;
        RECT 110.675 -127.325 111.005 -126.995 ;
        RECT 110.675 -128.685 111.005 -128.355 ;
        RECT 110.675 -130.045 111.005 -129.715 ;
        RECT 110.675 -131.405 111.005 -131.075 ;
        RECT 110.675 -132.765 111.005 -132.435 ;
        RECT 110.675 -134.125 111.005 -133.795 ;
        RECT 110.675 -135.485 111.005 -135.155 ;
        RECT 110.675 -136.845 111.005 -136.515 ;
        RECT 110.675 -138.205 111.005 -137.875 ;
        RECT 110.675 -139.565 111.005 -139.235 ;
        RECT 110.675 -140.925 111.005 -140.595 ;
        RECT 110.675 -142.285 111.005 -141.955 ;
        RECT 110.675 -143.645 111.005 -143.315 ;
        RECT 110.675 -145.005 111.005 -144.675 ;
        RECT 110.675 -146.365 111.005 -146.035 ;
        RECT 110.675 -147.725 111.005 -147.395 ;
        RECT 110.675 -149.085 111.005 -148.755 ;
        RECT 110.675 -150.445 111.005 -150.115 ;
        RECT 110.675 -151.805 111.005 -151.475 ;
        RECT 110.675 -153.165 111.005 -152.835 ;
        RECT 110.675 -154.525 111.005 -154.195 ;
        RECT 110.675 -155.885 111.005 -155.555 ;
        RECT 110.675 -157.245 111.005 -156.915 ;
        RECT 110.675 -158.605 111.005 -158.275 ;
        RECT 110.675 -159.965 111.005 -159.635 ;
        RECT 110.675 -161.325 111.005 -160.995 ;
        RECT 110.675 -162.685 111.005 -162.355 ;
        RECT 110.675 -164.045 111.005 -163.715 ;
        RECT 110.675 -165.405 111.005 -165.075 ;
        RECT 110.675 -166.765 111.005 -166.435 ;
        RECT 110.675 -168.125 111.005 -167.795 ;
        RECT 110.675 -169.485 111.005 -169.155 ;
        RECT 110.675 -170.845 111.005 -170.515 ;
        RECT 110.675 -172.205 111.005 -171.875 ;
        RECT 110.675 -173.565 111.005 -173.235 ;
        RECT 110.675 -174.925 111.005 -174.595 ;
        RECT 110.675 -176.285 111.005 -175.955 ;
        RECT 110.675 -177.645 111.005 -177.315 ;
        RECT 110.675 -183.29 111.005 -182.16 ;
        RECT 110.68 -183.405 111 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 112.035 244.04 112.365 245.17 ;
        RECT 112.035 239.875 112.365 240.205 ;
        RECT 112.035 238.515 112.365 238.845 ;
        RECT 112.035 237.155 112.365 237.485 ;
        RECT 112.04 237.155 112.36 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 112.035 -96.045 112.365 -95.715 ;
        RECT 112.035 -97.405 112.365 -97.075 ;
        RECT 112.035 -98.765 112.365 -98.435 ;
        RECT 112.035 -100.125 112.365 -99.795 ;
        RECT 112.035 -101.485 112.365 -101.155 ;
        RECT 112.035 -102.845 112.365 -102.515 ;
        RECT 112.035 -104.205 112.365 -103.875 ;
        RECT 112.035 -105.565 112.365 -105.235 ;
        RECT 112.035 -106.925 112.365 -106.595 ;
        RECT 112.035 -108.285 112.365 -107.955 ;
        RECT 112.035 -109.645 112.365 -109.315 ;
        RECT 112.035 -111.005 112.365 -110.675 ;
        RECT 112.035 -112.365 112.365 -112.035 ;
        RECT 112.035 -113.725 112.365 -113.395 ;
        RECT 112.035 -115.085 112.365 -114.755 ;
        RECT 112.035 -116.445 112.365 -116.115 ;
        RECT 112.035 -117.805 112.365 -117.475 ;
        RECT 112.035 -119.165 112.365 -118.835 ;
        RECT 112.035 -120.525 112.365 -120.195 ;
        RECT 112.035 -121.885 112.365 -121.555 ;
        RECT 112.035 -123.245 112.365 -122.915 ;
        RECT 112.035 -124.605 112.365 -124.275 ;
        RECT 112.035 -125.965 112.365 -125.635 ;
        RECT 112.035 -127.325 112.365 -126.995 ;
        RECT 112.035 -128.685 112.365 -128.355 ;
        RECT 112.035 -130.045 112.365 -129.715 ;
        RECT 112.035 -131.405 112.365 -131.075 ;
        RECT 112.035 -132.765 112.365 -132.435 ;
        RECT 112.035 -134.125 112.365 -133.795 ;
        RECT 112.035 -135.485 112.365 -135.155 ;
        RECT 112.035 -136.845 112.365 -136.515 ;
        RECT 112.035 -138.205 112.365 -137.875 ;
        RECT 112.035 -139.565 112.365 -139.235 ;
        RECT 112.035 -140.925 112.365 -140.595 ;
        RECT 112.035 -142.285 112.365 -141.955 ;
        RECT 112.035 -143.645 112.365 -143.315 ;
        RECT 112.035 -145.005 112.365 -144.675 ;
        RECT 112.035 -146.365 112.365 -146.035 ;
        RECT 112.035 -147.725 112.365 -147.395 ;
        RECT 112.035 -149.085 112.365 -148.755 ;
        RECT 112.035 -150.445 112.365 -150.115 ;
        RECT 112.035 -151.805 112.365 -151.475 ;
        RECT 112.035 -153.165 112.365 -152.835 ;
        RECT 112.035 -154.525 112.365 -154.195 ;
        RECT 112.035 -155.885 112.365 -155.555 ;
        RECT 112.035 -157.245 112.365 -156.915 ;
        RECT 112.035 -158.605 112.365 -158.275 ;
        RECT 112.035 -159.965 112.365 -159.635 ;
        RECT 112.035 -161.325 112.365 -160.995 ;
        RECT 112.035 -162.685 112.365 -162.355 ;
        RECT 112.035 -164.045 112.365 -163.715 ;
        RECT 112.035 -165.405 112.365 -165.075 ;
        RECT 112.035 -166.765 112.365 -166.435 ;
        RECT 112.035 -168.125 112.365 -167.795 ;
        RECT 112.035 -169.485 112.365 -169.155 ;
        RECT 112.035 -170.845 112.365 -170.515 ;
        RECT 112.035 -172.205 112.365 -171.875 ;
        RECT 112.035 -173.565 112.365 -173.235 ;
        RECT 112.035 -174.925 112.365 -174.595 ;
        RECT 112.035 -176.285 112.365 -175.955 ;
        RECT 112.035 -177.645 112.365 -177.315 ;
        RECT 112.035 -183.29 112.365 -182.16 ;
        RECT 112.04 -183.405 112.36 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 112.46 -94.075 112.79 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 113.395 244.04 113.725 245.17 ;
        RECT 113.395 239.875 113.725 240.205 ;
        RECT 113.395 238.515 113.725 238.845 ;
        RECT 113.395 237.155 113.725 237.485 ;
        RECT 113.4 237.155 113.72 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 114.755 244.04 115.085 245.17 ;
        RECT 114.755 239.875 115.085 240.205 ;
        RECT 114.755 238.515 115.085 238.845 ;
        RECT 114.755 237.155 115.085 237.485 ;
        RECT 114.76 237.155 115.08 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 114.755 -0.845 115.085 -0.515 ;
        RECT 114.755 -2.205 115.085 -1.875 ;
        RECT 114.755 -3.565 115.085 -3.235 ;
        RECT 114.76 -3.565 115.08 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 116.115 244.04 116.445 245.17 ;
        RECT 116.115 239.875 116.445 240.205 ;
        RECT 116.115 238.515 116.445 238.845 ;
        RECT 116.115 237.155 116.445 237.485 ;
        RECT 116.12 237.155 116.44 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 116.115 -0.845 116.445 -0.515 ;
        RECT 116.115 -2.205 116.445 -1.875 ;
        RECT 116.115 -3.565 116.445 -3.235 ;
        RECT 116.12 -3.565 116.44 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 117.475 244.04 117.805 245.17 ;
        RECT 117.475 239.875 117.805 240.205 ;
        RECT 117.475 238.515 117.805 238.845 ;
        RECT 117.475 237.155 117.805 237.485 ;
        RECT 117.48 237.155 117.8 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 117.475 -0.845 117.805 -0.515 ;
        RECT 117.475 -2.205 117.805 -1.875 ;
        RECT 117.475 -3.565 117.805 -3.235 ;
        RECT 117.48 -3.565 117.8 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 117.475 -91.965 117.805 -91.635 ;
        RECT 117.475 -93.325 117.805 -92.995 ;
        RECT 117.475 -94.685 117.805 -94.355 ;
        RECT 117.475 -96.045 117.805 -95.715 ;
        RECT 117.475 -97.405 117.805 -97.075 ;
        RECT 117.475 -98.765 117.805 -98.435 ;
        RECT 117.475 -100.125 117.805 -99.795 ;
        RECT 117.475 -101.485 117.805 -101.155 ;
        RECT 117.475 -102.845 117.805 -102.515 ;
        RECT 117.475 -104.205 117.805 -103.875 ;
        RECT 117.475 -105.565 117.805 -105.235 ;
        RECT 117.475 -106.925 117.805 -106.595 ;
        RECT 117.475 -108.285 117.805 -107.955 ;
        RECT 117.475 -109.645 117.805 -109.315 ;
        RECT 117.475 -111.005 117.805 -110.675 ;
        RECT 117.475 -112.365 117.805 -112.035 ;
        RECT 117.475 -113.725 117.805 -113.395 ;
        RECT 117.475 -115.085 117.805 -114.755 ;
        RECT 117.475 -116.445 117.805 -116.115 ;
        RECT 117.475 -117.805 117.805 -117.475 ;
        RECT 117.475 -119.165 117.805 -118.835 ;
        RECT 117.475 -120.525 117.805 -120.195 ;
        RECT 117.475 -121.885 117.805 -121.555 ;
        RECT 117.475 -123.245 117.805 -122.915 ;
        RECT 117.475 -124.605 117.805 -124.275 ;
        RECT 117.475 -125.965 117.805 -125.635 ;
        RECT 117.475 -127.325 117.805 -126.995 ;
        RECT 117.475 -128.685 117.805 -128.355 ;
        RECT 117.475 -130.045 117.805 -129.715 ;
        RECT 117.475 -131.405 117.805 -131.075 ;
        RECT 117.475 -132.765 117.805 -132.435 ;
        RECT 117.475 -134.125 117.805 -133.795 ;
        RECT 117.475 -135.485 117.805 -135.155 ;
        RECT 117.475 -136.845 117.805 -136.515 ;
        RECT 117.475 -138.205 117.805 -137.875 ;
        RECT 117.475 -139.565 117.805 -139.235 ;
        RECT 117.475 -140.925 117.805 -140.595 ;
        RECT 117.475 -142.285 117.805 -141.955 ;
        RECT 117.475 -143.645 117.805 -143.315 ;
        RECT 117.475 -145.005 117.805 -144.675 ;
        RECT 117.475 -146.365 117.805 -146.035 ;
        RECT 117.475 -147.725 117.805 -147.395 ;
        RECT 117.475 -149.085 117.805 -148.755 ;
        RECT 117.475 -150.445 117.805 -150.115 ;
        RECT 117.475 -151.805 117.805 -151.475 ;
        RECT 117.475 -153.165 117.805 -152.835 ;
        RECT 117.475 -154.525 117.805 -154.195 ;
        RECT 117.475 -155.885 117.805 -155.555 ;
        RECT 117.475 -157.245 117.805 -156.915 ;
        RECT 117.475 -158.605 117.805 -158.275 ;
        RECT 117.475 -159.965 117.805 -159.635 ;
        RECT 117.475 -161.325 117.805 -160.995 ;
        RECT 117.475 -162.685 117.805 -162.355 ;
        RECT 117.475 -164.045 117.805 -163.715 ;
        RECT 117.475 -165.405 117.805 -165.075 ;
        RECT 117.475 -166.765 117.805 -166.435 ;
        RECT 117.475 -168.125 117.805 -167.795 ;
        RECT 117.475 -169.485 117.805 -169.155 ;
        RECT 117.475 -170.845 117.805 -170.515 ;
        RECT 117.475 -172.205 117.805 -171.875 ;
        RECT 117.475 -173.565 117.805 -173.235 ;
        RECT 117.475 -174.925 117.805 -174.595 ;
        RECT 117.475 -176.285 117.805 -175.955 ;
        RECT 117.475 -177.645 117.805 -177.315 ;
        RECT 117.475 -183.29 117.805 -182.16 ;
        RECT 117.48 -183.405 117.8 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 118.56 -94.075 118.89 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 118.835 244.04 119.165 245.17 ;
        RECT 118.835 239.875 119.165 240.205 ;
        RECT 118.835 238.515 119.165 238.845 ;
        RECT 118.835 237.155 119.165 237.485 ;
        RECT 118.84 237.155 119.16 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 118.835 -96.045 119.165 -95.715 ;
        RECT 118.835 -97.405 119.165 -97.075 ;
        RECT 118.835 -98.765 119.165 -98.435 ;
        RECT 118.835 -100.125 119.165 -99.795 ;
        RECT 118.835 -101.485 119.165 -101.155 ;
        RECT 118.835 -102.845 119.165 -102.515 ;
        RECT 118.835 -104.205 119.165 -103.875 ;
        RECT 118.835 -105.565 119.165 -105.235 ;
        RECT 118.835 -106.925 119.165 -106.595 ;
        RECT 118.835 -108.285 119.165 -107.955 ;
        RECT 118.835 -109.645 119.165 -109.315 ;
        RECT 118.835 -111.005 119.165 -110.675 ;
        RECT 118.835 -112.365 119.165 -112.035 ;
        RECT 118.835 -113.725 119.165 -113.395 ;
        RECT 118.835 -115.085 119.165 -114.755 ;
        RECT 118.835 -116.445 119.165 -116.115 ;
        RECT 118.835 -117.805 119.165 -117.475 ;
        RECT 118.835 -119.165 119.165 -118.835 ;
        RECT 118.835 -120.525 119.165 -120.195 ;
        RECT 118.835 -121.885 119.165 -121.555 ;
        RECT 118.835 -123.245 119.165 -122.915 ;
        RECT 118.835 -124.605 119.165 -124.275 ;
        RECT 118.835 -125.965 119.165 -125.635 ;
        RECT 118.835 -127.325 119.165 -126.995 ;
        RECT 118.835 -128.685 119.165 -128.355 ;
        RECT 118.835 -130.045 119.165 -129.715 ;
        RECT 118.835 -131.405 119.165 -131.075 ;
        RECT 118.835 -132.765 119.165 -132.435 ;
        RECT 118.835 -134.125 119.165 -133.795 ;
        RECT 118.835 -135.485 119.165 -135.155 ;
        RECT 118.835 -136.845 119.165 -136.515 ;
        RECT 118.835 -138.205 119.165 -137.875 ;
        RECT 118.835 -139.565 119.165 -139.235 ;
        RECT 118.835 -140.925 119.165 -140.595 ;
        RECT 118.835 -142.285 119.165 -141.955 ;
        RECT 118.835 -143.645 119.165 -143.315 ;
        RECT 118.835 -145.005 119.165 -144.675 ;
        RECT 118.835 -146.365 119.165 -146.035 ;
        RECT 118.835 -147.725 119.165 -147.395 ;
        RECT 118.835 -149.085 119.165 -148.755 ;
        RECT 118.835 -150.445 119.165 -150.115 ;
        RECT 118.835 -151.805 119.165 -151.475 ;
        RECT 118.835 -153.165 119.165 -152.835 ;
        RECT 118.835 -154.525 119.165 -154.195 ;
        RECT 118.835 -155.885 119.165 -155.555 ;
        RECT 118.835 -157.245 119.165 -156.915 ;
        RECT 118.835 -158.605 119.165 -158.275 ;
        RECT 118.835 -159.965 119.165 -159.635 ;
        RECT 118.835 -161.325 119.165 -160.995 ;
        RECT 118.835 -162.685 119.165 -162.355 ;
        RECT 118.835 -164.045 119.165 -163.715 ;
        RECT 118.835 -165.405 119.165 -165.075 ;
        RECT 118.835 -166.765 119.165 -166.435 ;
        RECT 118.835 -168.125 119.165 -167.795 ;
        RECT 118.835 -169.485 119.165 -169.155 ;
        RECT 118.835 -170.845 119.165 -170.515 ;
        RECT 118.835 -172.205 119.165 -171.875 ;
        RECT 118.835 -173.565 119.165 -173.235 ;
        RECT 118.835 -174.925 119.165 -174.595 ;
        RECT 118.835 -176.285 119.165 -175.955 ;
        RECT 118.835 -177.645 119.165 -177.315 ;
        RECT 118.835 -183.29 119.165 -182.16 ;
        RECT 118.84 -183.405 119.16 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 120.195 244.04 120.525 245.17 ;
        RECT 120.195 239.875 120.525 240.205 ;
        RECT 120.195 238.515 120.525 238.845 ;
        RECT 120.195 237.155 120.525 237.485 ;
        RECT 120.2 237.155 120.52 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 120.195 -0.845 120.525 -0.515 ;
        RECT 120.195 -2.205 120.525 -1.875 ;
        RECT 120.195 -3.565 120.525 -3.235 ;
        RECT 120.2 -3.565 120.52 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 121.555 244.04 121.885 245.17 ;
        RECT 121.555 239.875 121.885 240.205 ;
        RECT 121.555 238.515 121.885 238.845 ;
        RECT 121.555 237.155 121.885 237.485 ;
        RECT 121.56 237.155 121.88 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 121.555 -0.845 121.885 -0.515 ;
        RECT 121.555 -2.205 121.885 -1.875 ;
        RECT 121.555 -3.565 121.885 -3.235 ;
        RECT 121.56 -3.565 121.88 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 122.915 244.04 123.245 245.17 ;
        RECT 122.915 239.875 123.245 240.205 ;
        RECT 122.915 238.515 123.245 238.845 ;
        RECT 122.915 237.155 123.245 237.485 ;
        RECT 122.92 237.155 123.24 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 122.915 -0.845 123.245 -0.515 ;
        RECT 122.915 -2.205 123.245 -1.875 ;
        RECT 122.915 -3.565 123.245 -3.235 ;
        RECT 122.92 -3.565 123.24 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 122.915 -91.965 123.245 -91.635 ;
        RECT 122.915 -93.325 123.245 -92.995 ;
        RECT 122.915 -94.685 123.245 -94.355 ;
        RECT 122.915 -96.045 123.245 -95.715 ;
        RECT 122.915 -97.405 123.245 -97.075 ;
        RECT 122.915 -98.765 123.245 -98.435 ;
        RECT 122.915 -100.125 123.245 -99.795 ;
        RECT 122.915 -101.485 123.245 -101.155 ;
        RECT 122.915 -102.845 123.245 -102.515 ;
        RECT 122.915 -104.205 123.245 -103.875 ;
        RECT 122.915 -105.565 123.245 -105.235 ;
        RECT 122.915 -106.925 123.245 -106.595 ;
        RECT 122.915 -108.285 123.245 -107.955 ;
        RECT 122.915 -109.645 123.245 -109.315 ;
        RECT 122.915 -111.005 123.245 -110.675 ;
        RECT 122.915 -112.365 123.245 -112.035 ;
        RECT 122.915 -113.725 123.245 -113.395 ;
        RECT 122.915 -115.085 123.245 -114.755 ;
        RECT 122.915 -116.445 123.245 -116.115 ;
        RECT 122.915 -117.805 123.245 -117.475 ;
        RECT 122.915 -119.165 123.245 -118.835 ;
        RECT 122.915 -120.525 123.245 -120.195 ;
        RECT 122.915 -121.885 123.245 -121.555 ;
        RECT 122.915 -123.245 123.245 -122.915 ;
        RECT 122.915 -124.605 123.245 -124.275 ;
        RECT 122.915 -125.965 123.245 -125.635 ;
        RECT 122.915 -127.325 123.245 -126.995 ;
        RECT 122.915 -128.685 123.245 -128.355 ;
        RECT 122.915 -130.045 123.245 -129.715 ;
        RECT 122.915 -131.405 123.245 -131.075 ;
        RECT 122.915 -132.765 123.245 -132.435 ;
        RECT 122.915 -134.125 123.245 -133.795 ;
        RECT 122.915 -135.485 123.245 -135.155 ;
        RECT 122.915 -136.845 123.245 -136.515 ;
        RECT 122.915 -138.205 123.245 -137.875 ;
        RECT 122.915 -139.565 123.245 -139.235 ;
        RECT 122.915 -140.925 123.245 -140.595 ;
        RECT 122.915 -142.285 123.245 -141.955 ;
        RECT 122.915 -143.645 123.245 -143.315 ;
        RECT 122.915 -145.005 123.245 -144.675 ;
        RECT 122.915 -146.365 123.245 -146.035 ;
        RECT 122.915 -147.725 123.245 -147.395 ;
        RECT 122.915 -149.085 123.245 -148.755 ;
        RECT 122.915 -150.445 123.245 -150.115 ;
        RECT 122.915 -151.805 123.245 -151.475 ;
        RECT 122.915 -153.165 123.245 -152.835 ;
        RECT 122.915 -154.525 123.245 -154.195 ;
        RECT 122.915 -155.885 123.245 -155.555 ;
        RECT 122.915 -157.245 123.245 -156.915 ;
        RECT 122.915 -158.605 123.245 -158.275 ;
        RECT 122.915 -159.965 123.245 -159.635 ;
        RECT 122.915 -161.325 123.245 -160.995 ;
        RECT 122.915 -162.685 123.245 -162.355 ;
        RECT 122.915 -164.045 123.245 -163.715 ;
        RECT 122.915 -165.405 123.245 -165.075 ;
        RECT 122.915 -166.765 123.245 -166.435 ;
        RECT 122.915 -168.125 123.245 -167.795 ;
        RECT 122.915 -169.485 123.245 -169.155 ;
        RECT 122.915 -170.845 123.245 -170.515 ;
        RECT 122.915 -172.205 123.245 -171.875 ;
        RECT 122.915 -173.565 123.245 -173.235 ;
        RECT 122.915 -174.925 123.245 -174.595 ;
        RECT 122.915 -176.285 123.245 -175.955 ;
        RECT 122.915 -177.645 123.245 -177.315 ;
        RECT 122.915 -183.29 123.245 -182.16 ;
        RECT 122.92 -183.405 123.24 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 124.275 244.04 124.605 245.17 ;
        RECT 124.275 239.875 124.605 240.205 ;
        RECT 124.275 238.515 124.605 238.845 ;
        RECT 124.275 237.155 124.605 237.485 ;
        RECT 124.28 237.155 124.6 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 124.275 -96.045 124.605 -95.715 ;
        RECT 124.275 -97.405 124.605 -97.075 ;
        RECT 124.275 -98.765 124.605 -98.435 ;
        RECT 124.275 -100.125 124.605 -99.795 ;
        RECT 124.275 -101.485 124.605 -101.155 ;
        RECT 124.275 -102.845 124.605 -102.515 ;
        RECT 124.275 -104.205 124.605 -103.875 ;
        RECT 124.275 -105.565 124.605 -105.235 ;
        RECT 124.275 -106.925 124.605 -106.595 ;
        RECT 124.275 -108.285 124.605 -107.955 ;
        RECT 124.275 -109.645 124.605 -109.315 ;
        RECT 124.275 -111.005 124.605 -110.675 ;
        RECT 124.275 -112.365 124.605 -112.035 ;
        RECT 124.275 -113.725 124.605 -113.395 ;
        RECT 124.275 -115.085 124.605 -114.755 ;
        RECT 124.275 -116.445 124.605 -116.115 ;
        RECT 124.275 -117.805 124.605 -117.475 ;
        RECT 124.275 -119.165 124.605 -118.835 ;
        RECT 124.275 -120.525 124.605 -120.195 ;
        RECT 124.275 -121.885 124.605 -121.555 ;
        RECT 124.275 -123.245 124.605 -122.915 ;
        RECT 124.275 -124.605 124.605 -124.275 ;
        RECT 124.275 -125.965 124.605 -125.635 ;
        RECT 124.275 -127.325 124.605 -126.995 ;
        RECT 124.275 -128.685 124.605 -128.355 ;
        RECT 124.275 -130.045 124.605 -129.715 ;
        RECT 124.275 -131.405 124.605 -131.075 ;
        RECT 124.275 -132.765 124.605 -132.435 ;
        RECT 124.275 -134.125 124.605 -133.795 ;
        RECT 124.275 -135.485 124.605 -135.155 ;
        RECT 124.275 -136.845 124.605 -136.515 ;
        RECT 124.275 -138.205 124.605 -137.875 ;
        RECT 124.275 -139.565 124.605 -139.235 ;
        RECT 124.275 -140.925 124.605 -140.595 ;
        RECT 124.275 -142.285 124.605 -141.955 ;
        RECT 124.275 -143.645 124.605 -143.315 ;
        RECT 124.275 -145.005 124.605 -144.675 ;
        RECT 124.275 -146.365 124.605 -146.035 ;
        RECT 124.275 -147.725 124.605 -147.395 ;
        RECT 124.275 -149.085 124.605 -148.755 ;
        RECT 124.275 -150.445 124.605 -150.115 ;
        RECT 124.275 -151.805 124.605 -151.475 ;
        RECT 124.275 -153.165 124.605 -152.835 ;
        RECT 124.275 -154.525 124.605 -154.195 ;
        RECT 124.275 -155.885 124.605 -155.555 ;
        RECT 124.275 -157.245 124.605 -156.915 ;
        RECT 124.275 -158.605 124.605 -158.275 ;
        RECT 124.275 -159.965 124.605 -159.635 ;
        RECT 124.275 -161.325 124.605 -160.995 ;
        RECT 124.275 -162.685 124.605 -162.355 ;
        RECT 124.275 -164.045 124.605 -163.715 ;
        RECT 124.275 -165.405 124.605 -165.075 ;
        RECT 124.275 -166.765 124.605 -166.435 ;
        RECT 124.275 -168.125 124.605 -167.795 ;
        RECT 124.275 -169.485 124.605 -169.155 ;
        RECT 124.275 -170.845 124.605 -170.515 ;
        RECT 124.275 -172.205 124.605 -171.875 ;
        RECT 124.275 -173.565 124.605 -173.235 ;
        RECT 124.275 -174.925 124.605 -174.595 ;
        RECT 124.275 -176.285 124.605 -175.955 ;
        RECT 124.275 -177.645 124.605 -177.315 ;
        RECT 124.275 -183.29 124.605 -182.16 ;
        RECT 124.28 -183.405 124.6 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 124.66 -94.075 124.99 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 125.635 244.04 125.965 245.17 ;
        RECT 125.635 239.875 125.965 240.205 ;
        RECT 125.635 238.515 125.965 238.845 ;
        RECT 125.635 237.155 125.965 237.485 ;
        RECT 125.64 237.155 125.96 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 126.995 244.04 127.325 245.17 ;
        RECT 126.995 239.875 127.325 240.205 ;
        RECT 126.995 238.515 127.325 238.845 ;
        RECT 126.995 237.155 127.325 237.485 ;
        RECT 127 237.155 127.32 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 126.995 -0.845 127.325 -0.515 ;
        RECT 126.995 -2.205 127.325 -1.875 ;
        RECT 126.995 -3.565 127.325 -3.235 ;
        RECT 127 -3.565 127.32 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 128.355 244.04 128.685 245.17 ;
        RECT 128.355 239.875 128.685 240.205 ;
        RECT 128.355 238.515 128.685 238.845 ;
        RECT 128.355 237.155 128.685 237.485 ;
        RECT 128.36 237.155 128.68 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 128.355 -0.845 128.685 -0.515 ;
        RECT 128.355 -2.205 128.685 -1.875 ;
        RECT 128.355 -3.565 128.685 -3.235 ;
        RECT 128.36 -3.565 128.68 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 128.355 -91.965 128.685 -91.635 ;
        RECT 128.355 -93.325 128.685 -92.995 ;
        RECT 128.355 -94.685 128.685 -94.355 ;
        RECT 128.355 -96.045 128.685 -95.715 ;
        RECT 128.355 -97.405 128.685 -97.075 ;
        RECT 128.355 -98.765 128.685 -98.435 ;
        RECT 128.355 -100.125 128.685 -99.795 ;
        RECT 128.355 -101.485 128.685 -101.155 ;
        RECT 128.355 -102.845 128.685 -102.515 ;
        RECT 128.355 -104.205 128.685 -103.875 ;
        RECT 128.355 -105.565 128.685 -105.235 ;
        RECT 128.355 -106.925 128.685 -106.595 ;
        RECT 128.355 -108.285 128.685 -107.955 ;
        RECT 128.355 -109.645 128.685 -109.315 ;
        RECT 128.355 -111.005 128.685 -110.675 ;
        RECT 128.355 -112.365 128.685 -112.035 ;
        RECT 128.355 -113.725 128.685 -113.395 ;
        RECT 128.355 -115.085 128.685 -114.755 ;
        RECT 128.355 -116.445 128.685 -116.115 ;
        RECT 128.355 -117.805 128.685 -117.475 ;
        RECT 128.355 -119.165 128.685 -118.835 ;
        RECT 128.355 -120.525 128.685 -120.195 ;
        RECT 128.355 -121.885 128.685 -121.555 ;
        RECT 128.355 -123.245 128.685 -122.915 ;
        RECT 128.355 -124.605 128.685 -124.275 ;
        RECT 128.355 -125.965 128.685 -125.635 ;
        RECT 128.355 -127.325 128.685 -126.995 ;
        RECT 128.355 -128.685 128.685 -128.355 ;
        RECT 128.355 -130.045 128.685 -129.715 ;
        RECT 128.355 -131.405 128.685 -131.075 ;
        RECT 128.355 -132.765 128.685 -132.435 ;
        RECT 128.355 -134.125 128.685 -133.795 ;
        RECT 128.355 -135.485 128.685 -135.155 ;
        RECT 128.355 -136.845 128.685 -136.515 ;
        RECT 128.355 -138.205 128.685 -137.875 ;
        RECT 128.355 -139.565 128.685 -139.235 ;
        RECT 128.355 -140.925 128.685 -140.595 ;
        RECT 128.355 -142.285 128.685 -141.955 ;
        RECT 128.355 -143.645 128.685 -143.315 ;
        RECT 128.355 -145.005 128.685 -144.675 ;
        RECT 128.355 -146.365 128.685 -146.035 ;
        RECT 128.355 -147.725 128.685 -147.395 ;
        RECT 128.355 -149.085 128.685 -148.755 ;
        RECT 128.355 -150.445 128.685 -150.115 ;
        RECT 128.355 -151.805 128.685 -151.475 ;
        RECT 128.355 -153.165 128.685 -152.835 ;
        RECT 128.355 -154.525 128.685 -154.195 ;
        RECT 128.355 -155.885 128.685 -155.555 ;
        RECT 128.355 -157.245 128.685 -156.915 ;
        RECT 128.355 -158.605 128.685 -158.275 ;
        RECT 128.355 -159.965 128.685 -159.635 ;
        RECT 128.355 -161.325 128.685 -160.995 ;
        RECT 128.355 -162.685 128.685 -162.355 ;
        RECT 128.355 -164.045 128.685 -163.715 ;
        RECT 128.355 -165.405 128.685 -165.075 ;
        RECT 128.355 -166.765 128.685 -166.435 ;
        RECT 128.355 -168.125 128.685 -167.795 ;
        RECT 128.355 -169.485 128.685 -169.155 ;
        RECT 128.355 -170.845 128.685 -170.515 ;
        RECT 128.355 -172.205 128.685 -171.875 ;
        RECT 128.355 -173.565 128.685 -173.235 ;
        RECT 128.355 -174.925 128.685 -174.595 ;
        RECT 128.355 -176.285 128.685 -175.955 ;
        RECT 128.355 -177.645 128.685 -177.315 ;
        RECT 128.355 -183.29 128.685 -182.16 ;
        RECT 128.36 -183.405 128.68 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.715 244.04 130.045 245.17 ;
        RECT 129.715 239.875 130.045 240.205 ;
        RECT 129.715 238.515 130.045 238.845 ;
        RECT 129.715 237.155 130.045 237.485 ;
        RECT 129.72 237.155 130.04 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.715 -0.845 130.045 -0.515 ;
        RECT 129.715 -2.205 130.045 -1.875 ;
        RECT 129.715 -3.565 130.045 -3.235 ;
        RECT 129.72 -3.565 130.04 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.715 -91.965 130.045 -91.635 ;
        RECT 129.715 -93.325 130.045 -92.995 ;
        RECT 129.715 -94.685 130.045 -94.355 ;
        RECT 129.715 -96.045 130.045 -95.715 ;
        RECT 129.715 -97.405 130.045 -97.075 ;
        RECT 129.715 -98.765 130.045 -98.435 ;
        RECT 129.715 -100.125 130.045 -99.795 ;
        RECT 129.715 -101.485 130.045 -101.155 ;
        RECT 129.715 -102.845 130.045 -102.515 ;
        RECT 129.715 -104.205 130.045 -103.875 ;
        RECT 129.715 -105.565 130.045 -105.235 ;
        RECT 129.715 -106.925 130.045 -106.595 ;
        RECT 129.715 -108.285 130.045 -107.955 ;
        RECT 129.715 -109.645 130.045 -109.315 ;
        RECT 129.715 -111.005 130.045 -110.675 ;
        RECT 129.715 -112.365 130.045 -112.035 ;
        RECT 129.715 -113.725 130.045 -113.395 ;
        RECT 129.715 -115.085 130.045 -114.755 ;
        RECT 129.715 -116.445 130.045 -116.115 ;
        RECT 129.715 -117.805 130.045 -117.475 ;
        RECT 129.715 -119.165 130.045 -118.835 ;
        RECT 129.715 -120.525 130.045 -120.195 ;
        RECT 129.715 -121.885 130.045 -121.555 ;
        RECT 129.715 -123.245 130.045 -122.915 ;
        RECT 129.715 -124.605 130.045 -124.275 ;
        RECT 129.715 -125.965 130.045 -125.635 ;
        RECT 129.715 -127.325 130.045 -126.995 ;
        RECT 129.715 -128.685 130.045 -128.355 ;
        RECT 129.715 -130.045 130.045 -129.715 ;
        RECT 129.715 -131.405 130.045 -131.075 ;
        RECT 129.715 -132.765 130.045 -132.435 ;
        RECT 129.715 -134.125 130.045 -133.795 ;
        RECT 129.715 -135.485 130.045 -135.155 ;
        RECT 129.715 -136.845 130.045 -136.515 ;
        RECT 129.715 -138.205 130.045 -137.875 ;
        RECT 129.715 -139.565 130.045 -139.235 ;
        RECT 129.715 -140.925 130.045 -140.595 ;
        RECT 129.715 -142.285 130.045 -141.955 ;
        RECT 129.715 -143.645 130.045 -143.315 ;
        RECT 129.715 -145.005 130.045 -144.675 ;
        RECT 129.715 -146.365 130.045 -146.035 ;
        RECT 129.715 -147.725 130.045 -147.395 ;
        RECT 129.715 -149.085 130.045 -148.755 ;
        RECT 129.715 -150.445 130.045 -150.115 ;
        RECT 129.715 -151.805 130.045 -151.475 ;
        RECT 129.715 -153.165 130.045 -152.835 ;
        RECT 129.715 -154.525 130.045 -154.195 ;
        RECT 129.715 -155.885 130.045 -155.555 ;
        RECT 129.715 -157.245 130.045 -156.915 ;
        RECT 129.715 -158.605 130.045 -158.275 ;
        RECT 129.715 -159.965 130.045 -159.635 ;
        RECT 129.715 -161.325 130.045 -160.995 ;
        RECT 129.715 -162.685 130.045 -162.355 ;
        RECT 129.715 -164.045 130.045 -163.715 ;
        RECT 129.715 -165.405 130.045 -165.075 ;
        RECT 129.715 -166.765 130.045 -166.435 ;
        RECT 129.715 -168.125 130.045 -167.795 ;
        RECT 129.715 -169.485 130.045 -169.155 ;
        RECT 129.715 -170.845 130.045 -170.515 ;
        RECT 129.715 -172.205 130.045 -171.875 ;
        RECT 129.715 -173.565 130.045 -173.235 ;
        RECT 129.715 -174.925 130.045 -174.595 ;
        RECT 129.715 -176.285 130.045 -175.955 ;
        RECT 129.715 -177.645 130.045 -177.315 ;
        RECT 129.715 -183.29 130.045 -182.16 ;
        RECT 129.72 -183.405 130.04 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 130.76 -94.075 131.09 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 131.075 244.04 131.405 245.17 ;
        RECT 131.075 239.875 131.405 240.205 ;
        RECT 131.075 238.515 131.405 238.845 ;
        RECT 131.075 237.155 131.405 237.485 ;
        RECT 131.08 237.155 131.4 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 131.075 -96.045 131.405 -95.715 ;
        RECT 131.075 -97.405 131.405 -97.075 ;
        RECT 131.075 -98.765 131.405 -98.435 ;
        RECT 131.075 -100.125 131.405 -99.795 ;
        RECT 131.075 -101.485 131.405 -101.155 ;
        RECT 131.075 -102.845 131.405 -102.515 ;
        RECT 131.075 -104.205 131.405 -103.875 ;
        RECT 131.075 -105.565 131.405 -105.235 ;
        RECT 131.075 -106.925 131.405 -106.595 ;
        RECT 131.075 -108.285 131.405 -107.955 ;
        RECT 131.075 -109.645 131.405 -109.315 ;
        RECT 131.075 -111.005 131.405 -110.675 ;
        RECT 131.075 -112.365 131.405 -112.035 ;
        RECT 131.075 -113.725 131.405 -113.395 ;
        RECT 131.075 -115.085 131.405 -114.755 ;
        RECT 131.075 -116.445 131.405 -116.115 ;
        RECT 131.075 -117.805 131.405 -117.475 ;
        RECT 131.075 -119.165 131.405 -118.835 ;
        RECT 131.075 -120.525 131.405 -120.195 ;
        RECT 131.075 -121.885 131.405 -121.555 ;
        RECT 131.075 -123.245 131.405 -122.915 ;
        RECT 131.075 -124.605 131.405 -124.275 ;
        RECT 131.075 -125.965 131.405 -125.635 ;
        RECT 131.075 -127.325 131.405 -126.995 ;
        RECT 131.075 -128.685 131.405 -128.355 ;
        RECT 131.075 -130.045 131.405 -129.715 ;
        RECT 131.075 -131.405 131.405 -131.075 ;
        RECT 131.075 -132.765 131.405 -132.435 ;
        RECT 131.075 -134.125 131.405 -133.795 ;
        RECT 131.075 -135.485 131.405 -135.155 ;
        RECT 131.075 -136.845 131.405 -136.515 ;
        RECT 131.075 -138.205 131.405 -137.875 ;
        RECT 131.075 -139.565 131.405 -139.235 ;
        RECT 131.075 -140.925 131.405 -140.595 ;
        RECT 131.075 -142.285 131.405 -141.955 ;
        RECT 131.075 -143.645 131.405 -143.315 ;
        RECT 131.075 -145.005 131.405 -144.675 ;
        RECT 131.075 -146.365 131.405 -146.035 ;
        RECT 131.075 -147.725 131.405 -147.395 ;
        RECT 131.075 -149.085 131.405 -148.755 ;
        RECT 131.075 -150.445 131.405 -150.115 ;
        RECT 131.075 -151.805 131.405 -151.475 ;
        RECT 131.075 -153.165 131.405 -152.835 ;
        RECT 131.075 -154.525 131.405 -154.195 ;
        RECT 131.075 -155.885 131.405 -155.555 ;
        RECT 131.075 -157.245 131.405 -156.915 ;
        RECT 131.075 -158.605 131.405 -158.275 ;
        RECT 131.075 -159.965 131.405 -159.635 ;
        RECT 131.075 -161.325 131.405 -160.995 ;
        RECT 131.075 -162.685 131.405 -162.355 ;
        RECT 131.075 -164.045 131.405 -163.715 ;
        RECT 131.075 -165.405 131.405 -165.075 ;
        RECT 131.075 -166.765 131.405 -166.435 ;
        RECT 131.075 -168.125 131.405 -167.795 ;
        RECT 131.075 -169.485 131.405 -169.155 ;
        RECT 131.075 -170.845 131.405 -170.515 ;
        RECT 131.075 -172.205 131.405 -171.875 ;
        RECT 131.075 -173.565 131.405 -173.235 ;
        RECT 131.075 -174.925 131.405 -174.595 ;
        RECT 131.075 -176.285 131.405 -175.955 ;
        RECT 131.075 -177.645 131.405 -177.315 ;
        RECT 131.075 -183.29 131.405 -182.16 ;
        RECT 131.08 -183.405 131.4 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 132.435 244.04 132.765 245.17 ;
        RECT 132.435 239.875 132.765 240.205 ;
        RECT 132.435 238.515 132.765 238.845 ;
        RECT 132.435 237.155 132.765 237.485 ;
        RECT 132.44 237.155 132.76 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 132.435 -0.845 132.765 -0.515 ;
        RECT 132.435 -2.205 132.765 -1.875 ;
        RECT 132.435 -3.565 132.765 -3.235 ;
        RECT 132.44 -3.565 132.76 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 133.795 244.04 134.125 245.17 ;
        RECT 133.795 239.875 134.125 240.205 ;
        RECT 133.795 238.515 134.125 238.845 ;
        RECT 133.795 237.155 134.125 237.485 ;
        RECT 133.8 237.155 134.12 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 133.795 -0.845 134.125 -0.515 ;
        RECT 133.795 -2.205 134.125 -1.875 ;
        RECT 133.795 -3.565 134.125 -3.235 ;
        RECT 133.8 -3.565 134.12 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 135.155 244.04 135.485 245.17 ;
        RECT 135.155 239.875 135.485 240.205 ;
        RECT 135.155 238.515 135.485 238.845 ;
        RECT 135.155 237.155 135.485 237.485 ;
        RECT 135.16 237.155 135.48 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 135.155 -0.845 135.485 -0.515 ;
        RECT 135.155 -2.205 135.485 -1.875 ;
        RECT 135.155 -3.565 135.485 -3.235 ;
        RECT 135.16 -3.565 135.48 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 135.155 -91.965 135.485 -91.635 ;
        RECT 135.155 -93.325 135.485 -92.995 ;
        RECT 135.155 -94.685 135.485 -94.355 ;
        RECT 135.155 -96.045 135.485 -95.715 ;
        RECT 135.155 -97.405 135.485 -97.075 ;
        RECT 135.155 -98.765 135.485 -98.435 ;
        RECT 135.155 -100.125 135.485 -99.795 ;
        RECT 135.155 -101.485 135.485 -101.155 ;
        RECT 135.155 -102.845 135.485 -102.515 ;
        RECT 135.155 -104.205 135.485 -103.875 ;
        RECT 135.155 -105.565 135.485 -105.235 ;
        RECT 135.155 -106.925 135.485 -106.595 ;
        RECT 135.155 -108.285 135.485 -107.955 ;
        RECT 135.155 -109.645 135.485 -109.315 ;
        RECT 135.155 -111.005 135.485 -110.675 ;
        RECT 135.155 -112.365 135.485 -112.035 ;
        RECT 135.155 -113.725 135.485 -113.395 ;
        RECT 135.155 -115.085 135.485 -114.755 ;
        RECT 135.155 -116.445 135.485 -116.115 ;
        RECT 135.155 -117.805 135.485 -117.475 ;
        RECT 135.155 -119.165 135.485 -118.835 ;
        RECT 135.155 -120.525 135.485 -120.195 ;
        RECT 135.155 -121.885 135.485 -121.555 ;
        RECT 135.155 -123.245 135.485 -122.915 ;
        RECT 135.155 -124.605 135.485 -124.275 ;
        RECT 135.155 -125.965 135.485 -125.635 ;
        RECT 135.155 -127.325 135.485 -126.995 ;
        RECT 135.155 -128.685 135.485 -128.355 ;
        RECT 135.155 -130.045 135.485 -129.715 ;
        RECT 135.155 -131.405 135.485 -131.075 ;
        RECT 135.155 -132.765 135.485 -132.435 ;
        RECT 135.155 -134.125 135.485 -133.795 ;
        RECT 135.155 -135.485 135.485 -135.155 ;
        RECT 135.155 -136.845 135.485 -136.515 ;
        RECT 135.155 -138.205 135.485 -137.875 ;
        RECT 135.155 -139.565 135.485 -139.235 ;
        RECT 135.155 -140.925 135.485 -140.595 ;
        RECT 135.155 -142.285 135.485 -141.955 ;
        RECT 135.155 -143.645 135.485 -143.315 ;
        RECT 135.155 -145.005 135.485 -144.675 ;
        RECT 135.155 -146.365 135.485 -146.035 ;
        RECT 135.155 -147.725 135.485 -147.395 ;
        RECT 135.155 -149.085 135.485 -148.755 ;
        RECT 135.155 -150.445 135.485 -150.115 ;
        RECT 135.155 -151.805 135.485 -151.475 ;
        RECT 135.155 -153.165 135.485 -152.835 ;
        RECT 135.155 -154.525 135.485 -154.195 ;
        RECT 135.155 -155.885 135.485 -155.555 ;
        RECT 135.155 -157.245 135.485 -156.915 ;
        RECT 135.155 -158.605 135.485 -158.275 ;
        RECT 135.155 -159.965 135.485 -159.635 ;
        RECT 135.155 -161.325 135.485 -160.995 ;
        RECT 135.155 -162.685 135.485 -162.355 ;
        RECT 135.155 -164.045 135.485 -163.715 ;
        RECT 135.155 -165.405 135.485 -165.075 ;
        RECT 135.155 -166.765 135.485 -166.435 ;
        RECT 135.155 -168.125 135.485 -167.795 ;
        RECT 135.155 -169.485 135.485 -169.155 ;
        RECT 135.155 -170.845 135.485 -170.515 ;
        RECT 135.155 -172.205 135.485 -171.875 ;
        RECT 135.155 -173.565 135.485 -173.235 ;
        RECT 135.155 -174.925 135.485 -174.595 ;
        RECT 135.155 -176.285 135.485 -175.955 ;
        RECT 135.155 -177.645 135.485 -177.315 ;
        RECT 135.155 -183.29 135.485 -182.16 ;
        RECT 135.16 -183.405 135.48 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 136.515 244.04 136.845 245.17 ;
        RECT 136.515 239.875 136.845 240.205 ;
        RECT 136.515 238.515 136.845 238.845 ;
        RECT 136.515 237.155 136.845 237.485 ;
        RECT 136.52 237.155 136.84 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 136.515 -96.045 136.845 -95.715 ;
        RECT 136.515 -97.405 136.845 -97.075 ;
        RECT 136.515 -98.765 136.845 -98.435 ;
        RECT 136.515 -100.125 136.845 -99.795 ;
        RECT 136.515 -101.485 136.845 -101.155 ;
        RECT 136.515 -102.845 136.845 -102.515 ;
        RECT 136.515 -104.205 136.845 -103.875 ;
        RECT 136.515 -105.565 136.845 -105.235 ;
        RECT 136.515 -106.925 136.845 -106.595 ;
        RECT 136.515 -108.285 136.845 -107.955 ;
        RECT 136.515 -109.645 136.845 -109.315 ;
        RECT 136.515 -111.005 136.845 -110.675 ;
        RECT 136.515 -112.365 136.845 -112.035 ;
        RECT 136.515 -113.725 136.845 -113.395 ;
        RECT 136.515 -115.085 136.845 -114.755 ;
        RECT 136.515 -116.445 136.845 -116.115 ;
        RECT 136.515 -117.805 136.845 -117.475 ;
        RECT 136.515 -119.165 136.845 -118.835 ;
        RECT 136.515 -120.525 136.845 -120.195 ;
        RECT 136.515 -121.885 136.845 -121.555 ;
        RECT 136.515 -123.245 136.845 -122.915 ;
        RECT 136.515 -124.605 136.845 -124.275 ;
        RECT 136.515 -125.965 136.845 -125.635 ;
        RECT 136.515 -127.325 136.845 -126.995 ;
        RECT 136.515 -128.685 136.845 -128.355 ;
        RECT 136.515 -130.045 136.845 -129.715 ;
        RECT 136.515 -131.405 136.845 -131.075 ;
        RECT 136.515 -132.765 136.845 -132.435 ;
        RECT 136.515 -134.125 136.845 -133.795 ;
        RECT 136.515 -135.485 136.845 -135.155 ;
        RECT 136.515 -136.845 136.845 -136.515 ;
        RECT 136.515 -138.205 136.845 -137.875 ;
        RECT 136.515 -139.565 136.845 -139.235 ;
        RECT 136.515 -140.925 136.845 -140.595 ;
        RECT 136.515 -142.285 136.845 -141.955 ;
        RECT 136.515 -143.645 136.845 -143.315 ;
        RECT 136.515 -145.005 136.845 -144.675 ;
        RECT 136.515 -146.365 136.845 -146.035 ;
        RECT 136.515 -147.725 136.845 -147.395 ;
        RECT 136.515 -149.085 136.845 -148.755 ;
        RECT 136.515 -150.445 136.845 -150.115 ;
        RECT 136.515 -151.805 136.845 -151.475 ;
        RECT 136.515 -153.165 136.845 -152.835 ;
        RECT 136.515 -154.525 136.845 -154.195 ;
        RECT 136.515 -155.885 136.845 -155.555 ;
        RECT 136.515 -157.245 136.845 -156.915 ;
        RECT 136.515 -158.605 136.845 -158.275 ;
        RECT 136.515 -159.965 136.845 -159.635 ;
        RECT 136.515 -161.325 136.845 -160.995 ;
        RECT 136.515 -162.685 136.845 -162.355 ;
        RECT 136.515 -164.045 136.845 -163.715 ;
        RECT 136.515 -165.405 136.845 -165.075 ;
        RECT 136.515 -166.765 136.845 -166.435 ;
        RECT 136.515 -168.125 136.845 -167.795 ;
        RECT 136.515 -169.485 136.845 -169.155 ;
        RECT 136.515 -170.845 136.845 -170.515 ;
        RECT 136.515 -172.205 136.845 -171.875 ;
        RECT 136.515 -173.565 136.845 -173.235 ;
        RECT 136.515 -174.925 136.845 -174.595 ;
        RECT 136.515 -176.285 136.845 -175.955 ;
        RECT 136.515 -177.645 136.845 -177.315 ;
        RECT 136.515 -183.29 136.845 -182.16 ;
        RECT 136.52 -183.405 136.84 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 136.86 -94.075 137.19 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 137.875 237.155 138.205 237.485 ;
        RECT 137.88 237.155 138.2 245.285 ;
        RECT 137.875 244.04 138.205 245.17 ;
        RECT 137.875 239.875 138.205 240.205 ;
        RECT 137.875 238.515 138.205 238.845 ;
    END
    PORT
      LAYER met3 ;
        RECT 75.315 244.04 75.645 245.17 ;
        RECT 75.315 239.875 75.645 240.205 ;
        RECT 75.315 238.515 75.645 238.845 ;
        RECT 75.315 237.155 75.645 237.485 ;
        RECT 75.32 237.155 75.64 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 75.315 -96.045 75.645 -95.715 ;
        RECT 75.315 -97.405 75.645 -97.075 ;
        RECT 75.315 -98.765 75.645 -98.435 ;
        RECT 75.315 -100.125 75.645 -99.795 ;
        RECT 75.315 -101.485 75.645 -101.155 ;
        RECT 75.315 -102.845 75.645 -102.515 ;
        RECT 75.315 -104.205 75.645 -103.875 ;
        RECT 75.315 -105.565 75.645 -105.235 ;
        RECT 75.315 -106.925 75.645 -106.595 ;
        RECT 75.315 -108.285 75.645 -107.955 ;
        RECT 75.315 -109.645 75.645 -109.315 ;
        RECT 75.315 -111.005 75.645 -110.675 ;
        RECT 75.315 -112.365 75.645 -112.035 ;
        RECT 75.315 -113.725 75.645 -113.395 ;
        RECT 75.315 -115.085 75.645 -114.755 ;
        RECT 75.315 -116.445 75.645 -116.115 ;
        RECT 75.315 -117.805 75.645 -117.475 ;
        RECT 75.315 -119.165 75.645 -118.835 ;
        RECT 75.315 -120.525 75.645 -120.195 ;
        RECT 75.315 -121.885 75.645 -121.555 ;
        RECT 75.315 -123.245 75.645 -122.915 ;
        RECT 75.315 -124.605 75.645 -124.275 ;
        RECT 75.315 -125.965 75.645 -125.635 ;
        RECT 75.315 -127.325 75.645 -126.995 ;
        RECT 75.315 -128.685 75.645 -128.355 ;
        RECT 75.315 -130.045 75.645 -129.715 ;
        RECT 75.315 -131.405 75.645 -131.075 ;
        RECT 75.315 -132.765 75.645 -132.435 ;
        RECT 75.315 -134.125 75.645 -133.795 ;
        RECT 75.315 -135.485 75.645 -135.155 ;
        RECT 75.315 -136.845 75.645 -136.515 ;
        RECT 75.315 -138.205 75.645 -137.875 ;
        RECT 75.315 -139.565 75.645 -139.235 ;
        RECT 75.315 -140.925 75.645 -140.595 ;
        RECT 75.315 -142.285 75.645 -141.955 ;
        RECT 75.315 -143.645 75.645 -143.315 ;
        RECT 75.315 -145.005 75.645 -144.675 ;
        RECT 75.315 -146.365 75.645 -146.035 ;
        RECT 75.315 -147.725 75.645 -147.395 ;
        RECT 75.315 -149.085 75.645 -148.755 ;
        RECT 75.315 -150.445 75.645 -150.115 ;
        RECT 75.315 -151.805 75.645 -151.475 ;
        RECT 75.315 -153.165 75.645 -152.835 ;
        RECT 75.315 -154.525 75.645 -154.195 ;
        RECT 75.315 -155.885 75.645 -155.555 ;
        RECT 75.315 -157.245 75.645 -156.915 ;
        RECT 75.315 -158.605 75.645 -158.275 ;
        RECT 75.315 -159.965 75.645 -159.635 ;
        RECT 75.315 -161.325 75.645 -160.995 ;
        RECT 75.315 -162.685 75.645 -162.355 ;
        RECT 75.315 -164.045 75.645 -163.715 ;
        RECT 75.315 -165.405 75.645 -165.075 ;
        RECT 75.315 -166.765 75.645 -166.435 ;
        RECT 75.315 -168.125 75.645 -167.795 ;
        RECT 75.315 -169.485 75.645 -169.155 ;
        RECT 75.315 -170.845 75.645 -170.515 ;
        RECT 75.315 -172.205 75.645 -171.875 ;
        RECT 75.315 -173.565 75.645 -173.235 ;
        RECT 75.315 -174.925 75.645 -174.595 ;
        RECT 75.315 -176.285 75.645 -175.955 ;
        RECT 75.315 -177.645 75.645 -177.315 ;
        RECT 75.315 -183.29 75.645 -182.16 ;
        RECT 75.32 -183.405 75.64 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 75.86 -94.075 76.19 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 76.675 244.04 77.005 245.17 ;
        RECT 76.675 239.875 77.005 240.205 ;
        RECT 76.675 238.515 77.005 238.845 ;
        RECT 76.675 237.155 77.005 237.485 ;
        RECT 76.68 237.155 77 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 78.035 244.04 78.365 245.17 ;
        RECT 78.035 239.875 78.365 240.205 ;
        RECT 78.035 238.515 78.365 238.845 ;
        RECT 78.035 237.155 78.365 237.485 ;
        RECT 78.04 237.155 78.36 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 78.035 -0.845 78.365 -0.515 ;
        RECT 78.035 -2.205 78.365 -1.875 ;
        RECT 78.035 -3.565 78.365 -3.235 ;
        RECT 78.04 -3.565 78.36 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 78.035 -91.965 78.365 -91.635 ;
        RECT 78.035 -93.325 78.365 -92.995 ;
        RECT 78.035 -94.685 78.365 -94.355 ;
        RECT 78.035 -96.045 78.365 -95.715 ;
        RECT 78.035 -97.405 78.365 -97.075 ;
        RECT 78.035 -98.765 78.365 -98.435 ;
        RECT 78.035 -100.125 78.365 -99.795 ;
        RECT 78.035 -101.485 78.365 -101.155 ;
        RECT 78.035 -102.845 78.365 -102.515 ;
        RECT 78.035 -104.205 78.365 -103.875 ;
        RECT 78.035 -105.565 78.365 -105.235 ;
        RECT 78.035 -106.925 78.365 -106.595 ;
        RECT 78.035 -108.285 78.365 -107.955 ;
        RECT 78.035 -109.645 78.365 -109.315 ;
        RECT 78.035 -111.005 78.365 -110.675 ;
        RECT 78.035 -112.365 78.365 -112.035 ;
        RECT 78.035 -113.725 78.365 -113.395 ;
        RECT 78.035 -115.085 78.365 -114.755 ;
        RECT 78.035 -116.445 78.365 -116.115 ;
        RECT 78.035 -117.805 78.365 -117.475 ;
        RECT 78.035 -119.165 78.365 -118.835 ;
        RECT 78.035 -120.525 78.365 -120.195 ;
        RECT 78.035 -121.885 78.365 -121.555 ;
        RECT 78.035 -123.245 78.365 -122.915 ;
        RECT 78.035 -124.605 78.365 -124.275 ;
        RECT 78.035 -125.965 78.365 -125.635 ;
        RECT 78.035 -127.325 78.365 -126.995 ;
        RECT 78.035 -128.685 78.365 -128.355 ;
        RECT 78.035 -130.045 78.365 -129.715 ;
        RECT 78.035 -131.405 78.365 -131.075 ;
        RECT 78.035 -132.765 78.365 -132.435 ;
        RECT 78.035 -134.125 78.365 -133.795 ;
        RECT 78.035 -135.485 78.365 -135.155 ;
        RECT 78.035 -136.845 78.365 -136.515 ;
        RECT 78.035 -138.205 78.365 -137.875 ;
        RECT 78.035 -139.565 78.365 -139.235 ;
        RECT 78.035 -140.925 78.365 -140.595 ;
        RECT 78.035 -142.285 78.365 -141.955 ;
        RECT 78.035 -143.645 78.365 -143.315 ;
        RECT 78.035 -145.005 78.365 -144.675 ;
        RECT 78.035 -146.365 78.365 -146.035 ;
        RECT 78.035 -147.725 78.365 -147.395 ;
        RECT 78.035 -149.085 78.365 -148.755 ;
        RECT 78.035 -150.445 78.365 -150.115 ;
        RECT 78.035 -151.805 78.365 -151.475 ;
        RECT 78.035 -153.165 78.365 -152.835 ;
        RECT 78.035 -154.525 78.365 -154.195 ;
        RECT 78.035 -155.885 78.365 -155.555 ;
        RECT 78.035 -157.245 78.365 -156.915 ;
        RECT 78.035 -158.605 78.365 -158.275 ;
        RECT 78.035 -159.965 78.365 -159.635 ;
        RECT 78.035 -161.325 78.365 -160.995 ;
        RECT 78.035 -162.685 78.365 -162.355 ;
        RECT 78.035 -164.045 78.365 -163.715 ;
        RECT 78.035 -165.405 78.365 -165.075 ;
        RECT 78.035 -166.765 78.365 -166.435 ;
        RECT 78.035 -168.125 78.365 -167.795 ;
        RECT 78.035 -169.485 78.365 -169.155 ;
        RECT 78.035 -170.845 78.365 -170.515 ;
        RECT 78.035 -172.205 78.365 -171.875 ;
        RECT 78.035 -173.565 78.365 -173.235 ;
        RECT 78.035 -174.925 78.365 -174.595 ;
        RECT 78.035 -176.285 78.365 -175.955 ;
        RECT 78.035 -177.645 78.365 -177.315 ;
        RECT 78.035 -183.29 78.365 -182.16 ;
        RECT 78.04 -183.405 78.36 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 79.395 244.04 79.725 245.17 ;
        RECT 79.395 239.875 79.725 240.205 ;
        RECT 79.395 238.515 79.725 238.845 ;
        RECT 79.395 237.155 79.725 237.485 ;
        RECT 79.4 237.155 79.72 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 79.395 -0.845 79.725 -0.515 ;
        RECT 79.395 -2.205 79.725 -1.875 ;
        RECT 79.395 -3.565 79.725 -3.235 ;
        RECT 79.4 -3.565 79.72 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 80.755 244.04 81.085 245.17 ;
        RECT 80.755 239.875 81.085 240.205 ;
        RECT 80.755 238.515 81.085 238.845 ;
        RECT 80.755 237.155 81.085 237.485 ;
        RECT 80.76 237.155 81.08 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 80.755 -0.845 81.085 -0.515 ;
        RECT 80.755 -2.205 81.085 -1.875 ;
        RECT 80.755 -3.565 81.085 -3.235 ;
        RECT 80.76 -3.565 81.08 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 80.755 -91.965 81.085 -91.635 ;
        RECT 80.755 -93.325 81.085 -92.995 ;
        RECT 80.755 -94.685 81.085 -94.355 ;
        RECT 80.755 -96.045 81.085 -95.715 ;
        RECT 80.755 -97.405 81.085 -97.075 ;
        RECT 80.755 -98.765 81.085 -98.435 ;
        RECT 80.755 -100.125 81.085 -99.795 ;
        RECT 80.755 -101.485 81.085 -101.155 ;
        RECT 80.755 -102.845 81.085 -102.515 ;
        RECT 80.755 -104.205 81.085 -103.875 ;
        RECT 80.755 -105.565 81.085 -105.235 ;
        RECT 80.755 -106.925 81.085 -106.595 ;
        RECT 80.755 -108.285 81.085 -107.955 ;
        RECT 80.755 -109.645 81.085 -109.315 ;
        RECT 80.755 -111.005 81.085 -110.675 ;
        RECT 80.755 -112.365 81.085 -112.035 ;
        RECT 80.755 -113.725 81.085 -113.395 ;
        RECT 80.755 -115.085 81.085 -114.755 ;
        RECT 80.755 -116.445 81.085 -116.115 ;
        RECT 80.755 -117.805 81.085 -117.475 ;
        RECT 80.755 -119.165 81.085 -118.835 ;
        RECT 80.755 -120.525 81.085 -120.195 ;
        RECT 80.755 -121.885 81.085 -121.555 ;
        RECT 80.755 -123.245 81.085 -122.915 ;
        RECT 80.755 -124.605 81.085 -124.275 ;
        RECT 80.755 -125.965 81.085 -125.635 ;
        RECT 80.755 -127.325 81.085 -126.995 ;
        RECT 80.755 -128.685 81.085 -128.355 ;
        RECT 80.755 -130.045 81.085 -129.715 ;
        RECT 80.755 -131.405 81.085 -131.075 ;
        RECT 80.755 -132.765 81.085 -132.435 ;
        RECT 80.755 -134.125 81.085 -133.795 ;
        RECT 80.755 -135.485 81.085 -135.155 ;
        RECT 80.755 -136.845 81.085 -136.515 ;
        RECT 80.755 -138.205 81.085 -137.875 ;
        RECT 80.755 -139.565 81.085 -139.235 ;
        RECT 80.755 -140.925 81.085 -140.595 ;
        RECT 80.755 -142.285 81.085 -141.955 ;
        RECT 80.755 -143.645 81.085 -143.315 ;
        RECT 80.755 -145.005 81.085 -144.675 ;
        RECT 80.755 -146.365 81.085 -146.035 ;
        RECT 80.755 -147.725 81.085 -147.395 ;
        RECT 80.755 -149.085 81.085 -148.755 ;
        RECT 80.755 -150.445 81.085 -150.115 ;
        RECT 80.755 -151.805 81.085 -151.475 ;
        RECT 80.755 -153.165 81.085 -152.835 ;
        RECT 80.755 -154.525 81.085 -154.195 ;
        RECT 80.755 -155.885 81.085 -155.555 ;
        RECT 80.755 -157.245 81.085 -156.915 ;
        RECT 80.755 -158.605 81.085 -158.275 ;
        RECT 80.755 -159.965 81.085 -159.635 ;
        RECT 80.755 -161.325 81.085 -160.995 ;
        RECT 80.755 -162.685 81.085 -162.355 ;
        RECT 80.755 -164.045 81.085 -163.715 ;
        RECT 80.755 -165.405 81.085 -165.075 ;
        RECT 80.755 -166.765 81.085 -166.435 ;
        RECT 80.755 -168.125 81.085 -167.795 ;
        RECT 80.755 -169.485 81.085 -169.155 ;
        RECT 80.755 -170.845 81.085 -170.515 ;
        RECT 80.755 -172.205 81.085 -171.875 ;
        RECT 80.755 -173.565 81.085 -173.235 ;
        RECT 80.755 -174.925 81.085 -174.595 ;
        RECT 80.755 -176.285 81.085 -175.955 ;
        RECT 80.755 -177.645 81.085 -177.315 ;
        RECT 80.755 -183.29 81.085 -182.16 ;
        RECT 80.76 -183.405 81.08 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 81.96 -94.075 82.29 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 82.115 244.04 82.445 245.17 ;
        RECT 82.115 239.875 82.445 240.205 ;
        RECT 82.115 238.515 82.445 238.845 ;
        RECT 82.115 237.155 82.445 237.485 ;
        RECT 82.12 237.155 82.44 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 82.115 -96.045 82.445 -95.715 ;
        RECT 82.115 -97.405 82.445 -97.075 ;
        RECT 82.115 -98.765 82.445 -98.435 ;
        RECT 82.115 -100.125 82.445 -99.795 ;
        RECT 82.115 -101.485 82.445 -101.155 ;
        RECT 82.115 -102.845 82.445 -102.515 ;
        RECT 82.115 -104.205 82.445 -103.875 ;
        RECT 82.115 -105.565 82.445 -105.235 ;
        RECT 82.115 -106.925 82.445 -106.595 ;
        RECT 82.115 -108.285 82.445 -107.955 ;
        RECT 82.115 -109.645 82.445 -109.315 ;
        RECT 82.115 -111.005 82.445 -110.675 ;
        RECT 82.115 -112.365 82.445 -112.035 ;
        RECT 82.115 -113.725 82.445 -113.395 ;
        RECT 82.115 -115.085 82.445 -114.755 ;
        RECT 82.115 -116.445 82.445 -116.115 ;
        RECT 82.115 -117.805 82.445 -117.475 ;
        RECT 82.115 -119.165 82.445 -118.835 ;
        RECT 82.115 -120.525 82.445 -120.195 ;
        RECT 82.115 -121.885 82.445 -121.555 ;
        RECT 82.115 -123.245 82.445 -122.915 ;
        RECT 82.115 -124.605 82.445 -124.275 ;
        RECT 82.115 -125.965 82.445 -125.635 ;
        RECT 82.115 -127.325 82.445 -126.995 ;
        RECT 82.115 -128.685 82.445 -128.355 ;
        RECT 82.115 -130.045 82.445 -129.715 ;
        RECT 82.115 -131.405 82.445 -131.075 ;
        RECT 82.115 -132.765 82.445 -132.435 ;
        RECT 82.115 -134.125 82.445 -133.795 ;
        RECT 82.115 -135.485 82.445 -135.155 ;
        RECT 82.115 -136.845 82.445 -136.515 ;
        RECT 82.115 -138.205 82.445 -137.875 ;
        RECT 82.115 -139.565 82.445 -139.235 ;
        RECT 82.115 -140.925 82.445 -140.595 ;
        RECT 82.115 -142.285 82.445 -141.955 ;
        RECT 82.115 -143.645 82.445 -143.315 ;
        RECT 82.115 -145.005 82.445 -144.675 ;
        RECT 82.115 -146.365 82.445 -146.035 ;
        RECT 82.115 -147.725 82.445 -147.395 ;
        RECT 82.115 -149.085 82.445 -148.755 ;
        RECT 82.115 -150.445 82.445 -150.115 ;
        RECT 82.115 -151.805 82.445 -151.475 ;
        RECT 82.115 -153.165 82.445 -152.835 ;
        RECT 82.115 -154.525 82.445 -154.195 ;
        RECT 82.115 -155.885 82.445 -155.555 ;
        RECT 82.115 -157.245 82.445 -156.915 ;
        RECT 82.115 -158.605 82.445 -158.275 ;
        RECT 82.115 -159.965 82.445 -159.635 ;
        RECT 82.115 -161.325 82.445 -160.995 ;
        RECT 82.115 -162.685 82.445 -162.355 ;
        RECT 82.115 -164.045 82.445 -163.715 ;
        RECT 82.115 -165.405 82.445 -165.075 ;
        RECT 82.115 -166.765 82.445 -166.435 ;
        RECT 82.115 -168.125 82.445 -167.795 ;
        RECT 82.115 -169.485 82.445 -169.155 ;
        RECT 82.115 -170.845 82.445 -170.515 ;
        RECT 82.115 -172.205 82.445 -171.875 ;
        RECT 82.115 -173.565 82.445 -173.235 ;
        RECT 82.115 -174.925 82.445 -174.595 ;
        RECT 82.115 -176.285 82.445 -175.955 ;
        RECT 82.115 -177.645 82.445 -177.315 ;
        RECT 82.115 -183.29 82.445 -182.16 ;
        RECT 82.12 -183.405 82.44 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 83.475 244.04 83.805 245.17 ;
        RECT 83.475 239.875 83.805 240.205 ;
        RECT 83.475 238.515 83.805 238.845 ;
        RECT 83.475 237.155 83.805 237.485 ;
        RECT 83.48 237.155 83.8 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 83.475 -0.845 83.805 -0.515 ;
        RECT 83.475 -2.205 83.805 -1.875 ;
        RECT 83.475 -3.565 83.805 -3.235 ;
        RECT 83.48 -3.565 83.8 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 84.835 244.04 85.165 245.17 ;
        RECT 84.835 239.875 85.165 240.205 ;
        RECT 84.835 238.515 85.165 238.845 ;
        RECT 84.835 237.155 85.165 237.485 ;
        RECT 84.84 237.155 85.16 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 84.835 -0.845 85.165 -0.515 ;
        RECT 84.835 -2.205 85.165 -1.875 ;
        RECT 84.835 -3.565 85.165 -3.235 ;
        RECT 84.84 -3.565 85.16 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 86.195 244.04 86.525 245.17 ;
        RECT 86.195 239.875 86.525 240.205 ;
        RECT 86.195 238.515 86.525 238.845 ;
        RECT 86.195 237.155 86.525 237.485 ;
        RECT 86.2 237.155 86.52 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 86.195 -0.845 86.525 -0.515 ;
        RECT 86.195 -2.205 86.525 -1.875 ;
        RECT 86.195 -3.565 86.525 -3.235 ;
        RECT 86.2 -3.565 86.52 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 86.195 -91.965 86.525 -91.635 ;
        RECT 86.195 -93.325 86.525 -92.995 ;
        RECT 86.195 -94.685 86.525 -94.355 ;
        RECT 86.195 -96.045 86.525 -95.715 ;
        RECT 86.195 -97.405 86.525 -97.075 ;
        RECT 86.195 -98.765 86.525 -98.435 ;
        RECT 86.195 -100.125 86.525 -99.795 ;
        RECT 86.195 -101.485 86.525 -101.155 ;
        RECT 86.195 -102.845 86.525 -102.515 ;
        RECT 86.195 -104.205 86.525 -103.875 ;
        RECT 86.195 -105.565 86.525 -105.235 ;
        RECT 86.195 -106.925 86.525 -106.595 ;
        RECT 86.195 -108.285 86.525 -107.955 ;
        RECT 86.195 -109.645 86.525 -109.315 ;
        RECT 86.195 -111.005 86.525 -110.675 ;
        RECT 86.195 -112.365 86.525 -112.035 ;
        RECT 86.195 -113.725 86.525 -113.395 ;
        RECT 86.195 -115.085 86.525 -114.755 ;
        RECT 86.195 -116.445 86.525 -116.115 ;
        RECT 86.195 -117.805 86.525 -117.475 ;
        RECT 86.195 -119.165 86.525 -118.835 ;
        RECT 86.195 -120.525 86.525 -120.195 ;
        RECT 86.195 -121.885 86.525 -121.555 ;
        RECT 86.195 -123.245 86.525 -122.915 ;
        RECT 86.195 -124.605 86.525 -124.275 ;
        RECT 86.195 -125.965 86.525 -125.635 ;
        RECT 86.195 -127.325 86.525 -126.995 ;
        RECT 86.195 -128.685 86.525 -128.355 ;
        RECT 86.195 -130.045 86.525 -129.715 ;
        RECT 86.195 -131.405 86.525 -131.075 ;
        RECT 86.195 -132.765 86.525 -132.435 ;
        RECT 86.195 -134.125 86.525 -133.795 ;
        RECT 86.195 -135.485 86.525 -135.155 ;
        RECT 86.195 -136.845 86.525 -136.515 ;
        RECT 86.195 -138.205 86.525 -137.875 ;
        RECT 86.195 -139.565 86.525 -139.235 ;
        RECT 86.195 -140.925 86.525 -140.595 ;
        RECT 86.195 -142.285 86.525 -141.955 ;
        RECT 86.195 -143.645 86.525 -143.315 ;
        RECT 86.195 -145.005 86.525 -144.675 ;
        RECT 86.195 -146.365 86.525 -146.035 ;
        RECT 86.195 -147.725 86.525 -147.395 ;
        RECT 86.195 -149.085 86.525 -148.755 ;
        RECT 86.195 -150.445 86.525 -150.115 ;
        RECT 86.195 -151.805 86.525 -151.475 ;
        RECT 86.195 -153.165 86.525 -152.835 ;
        RECT 86.195 -154.525 86.525 -154.195 ;
        RECT 86.195 -155.885 86.525 -155.555 ;
        RECT 86.195 -157.245 86.525 -156.915 ;
        RECT 86.195 -158.605 86.525 -158.275 ;
        RECT 86.195 -159.965 86.525 -159.635 ;
        RECT 86.195 -161.325 86.525 -160.995 ;
        RECT 86.195 -162.685 86.525 -162.355 ;
        RECT 86.195 -164.045 86.525 -163.715 ;
        RECT 86.195 -165.405 86.525 -165.075 ;
        RECT 86.195 -166.765 86.525 -166.435 ;
        RECT 86.195 -168.125 86.525 -167.795 ;
        RECT 86.195 -169.485 86.525 -169.155 ;
        RECT 86.195 -170.845 86.525 -170.515 ;
        RECT 86.195 -172.205 86.525 -171.875 ;
        RECT 86.195 -173.565 86.525 -173.235 ;
        RECT 86.195 -174.925 86.525 -174.595 ;
        RECT 86.195 -176.285 86.525 -175.955 ;
        RECT 86.195 -177.645 86.525 -177.315 ;
        RECT 86.195 -183.29 86.525 -182.16 ;
        RECT 86.2 -183.405 86.52 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 87.555 244.04 87.885 245.17 ;
        RECT 87.555 239.875 87.885 240.205 ;
        RECT 87.555 238.515 87.885 238.845 ;
        RECT 87.555 237.155 87.885 237.485 ;
        RECT 87.56 237.155 87.88 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 87.555 -96.045 87.885 -95.715 ;
        RECT 87.555 -97.405 87.885 -97.075 ;
        RECT 87.555 -98.765 87.885 -98.435 ;
        RECT 87.555 -100.125 87.885 -99.795 ;
        RECT 87.555 -101.485 87.885 -101.155 ;
        RECT 87.555 -102.845 87.885 -102.515 ;
        RECT 87.555 -104.205 87.885 -103.875 ;
        RECT 87.555 -105.565 87.885 -105.235 ;
        RECT 87.555 -106.925 87.885 -106.595 ;
        RECT 87.555 -108.285 87.885 -107.955 ;
        RECT 87.555 -109.645 87.885 -109.315 ;
        RECT 87.555 -111.005 87.885 -110.675 ;
        RECT 87.555 -112.365 87.885 -112.035 ;
        RECT 87.555 -113.725 87.885 -113.395 ;
        RECT 87.555 -115.085 87.885 -114.755 ;
        RECT 87.555 -116.445 87.885 -116.115 ;
        RECT 87.555 -117.805 87.885 -117.475 ;
        RECT 87.555 -119.165 87.885 -118.835 ;
        RECT 87.555 -120.525 87.885 -120.195 ;
        RECT 87.555 -121.885 87.885 -121.555 ;
        RECT 87.555 -123.245 87.885 -122.915 ;
        RECT 87.555 -124.605 87.885 -124.275 ;
        RECT 87.555 -125.965 87.885 -125.635 ;
        RECT 87.555 -127.325 87.885 -126.995 ;
        RECT 87.555 -128.685 87.885 -128.355 ;
        RECT 87.555 -130.045 87.885 -129.715 ;
        RECT 87.555 -131.405 87.885 -131.075 ;
        RECT 87.555 -132.765 87.885 -132.435 ;
        RECT 87.555 -134.125 87.885 -133.795 ;
        RECT 87.555 -135.485 87.885 -135.155 ;
        RECT 87.555 -136.845 87.885 -136.515 ;
        RECT 87.555 -138.205 87.885 -137.875 ;
        RECT 87.555 -139.565 87.885 -139.235 ;
        RECT 87.555 -140.925 87.885 -140.595 ;
        RECT 87.555 -142.285 87.885 -141.955 ;
        RECT 87.555 -143.645 87.885 -143.315 ;
        RECT 87.555 -145.005 87.885 -144.675 ;
        RECT 87.555 -146.365 87.885 -146.035 ;
        RECT 87.555 -147.725 87.885 -147.395 ;
        RECT 87.555 -149.085 87.885 -148.755 ;
        RECT 87.555 -150.445 87.885 -150.115 ;
        RECT 87.555 -151.805 87.885 -151.475 ;
        RECT 87.555 -153.165 87.885 -152.835 ;
        RECT 87.555 -154.525 87.885 -154.195 ;
        RECT 87.555 -155.885 87.885 -155.555 ;
        RECT 87.555 -157.245 87.885 -156.915 ;
        RECT 87.555 -158.605 87.885 -158.275 ;
        RECT 87.555 -159.965 87.885 -159.635 ;
        RECT 87.555 -161.325 87.885 -160.995 ;
        RECT 87.555 -162.685 87.885 -162.355 ;
        RECT 87.555 -164.045 87.885 -163.715 ;
        RECT 87.555 -165.405 87.885 -165.075 ;
        RECT 87.555 -166.765 87.885 -166.435 ;
        RECT 87.555 -168.125 87.885 -167.795 ;
        RECT 87.555 -169.485 87.885 -169.155 ;
        RECT 87.555 -170.845 87.885 -170.515 ;
        RECT 87.555 -172.205 87.885 -171.875 ;
        RECT 87.555 -173.565 87.885 -173.235 ;
        RECT 87.555 -174.925 87.885 -174.595 ;
        RECT 87.555 -176.285 87.885 -175.955 ;
        RECT 87.555 -177.645 87.885 -177.315 ;
        RECT 87.555 -183.29 87.885 -182.16 ;
        RECT 87.56 -183.405 87.88 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 88.06 -94.075 88.39 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 88.915 244.04 89.245 245.17 ;
        RECT 88.915 239.875 89.245 240.205 ;
        RECT 88.915 238.515 89.245 238.845 ;
        RECT 88.915 237.155 89.245 237.485 ;
        RECT 88.92 237.155 89.24 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 90.275 244.04 90.605 245.17 ;
        RECT 90.275 239.875 90.605 240.205 ;
        RECT 90.275 238.515 90.605 238.845 ;
        RECT 90.275 237.155 90.605 237.485 ;
        RECT 90.28 237.155 90.6 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 90.275 -0.845 90.605 -0.515 ;
        RECT 90.275 -2.205 90.605 -1.875 ;
        RECT 90.275 -3.565 90.605 -3.235 ;
        RECT 90.28 -3.565 90.6 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 90.275 -91.965 90.605 -91.635 ;
        RECT 90.275 -93.325 90.605 -92.995 ;
        RECT 90.275 -94.685 90.605 -94.355 ;
        RECT 90.275 -96.045 90.605 -95.715 ;
        RECT 90.275 -97.405 90.605 -97.075 ;
        RECT 90.275 -98.765 90.605 -98.435 ;
        RECT 90.275 -100.125 90.605 -99.795 ;
        RECT 90.275 -101.485 90.605 -101.155 ;
        RECT 90.275 -102.845 90.605 -102.515 ;
        RECT 90.275 -104.205 90.605 -103.875 ;
        RECT 90.275 -105.565 90.605 -105.235 ;
        RECT 90.275 -106.925 90.605 -106.595 ;
        RECT 90.275 -108.285 90.605 -107.955 ;
        RECT 90.275 -109.645 90.605 -109.315 ;
        RECT 90.275 -111.005 90.605 -110.675 ;
        RECT 90.275 -112.365 90.605 -112.035 ;
        RECT 90.275 -113.725 90.605 -113.395 ;
        RECT 90.275 -115.085 90.605 -114.755 ;
        RECT 90.275 -116.445 90.605 -116.115 ;
        RECT 90.275 -117.805 90.605 -117.475 ;
        RECT 90.275 -119.165 90.605 -118.835 ;
        RECT 90.275 -120.525 90.605 -120.195 ;
        RECT 90.275 -121.885 90.605 -121.555 ;
        RECT 90.275 -123.245 90.605 -122.915 ;
        RECT 90.275 -124.605 90.605 -124.275 ;
        RECT 90.275 -125.965 90.605 -125.635 ;
        RECT 90.275 -127.325 90.605 -126.995 ;
        RECT 90.275 -128.685 90.605 -128.355 ;
        RECT 90.275 -130.045 90.605 -129.715 ;
        RECT 90.275 -131.405 90.605 -131.075 ;
        RECT 90.275 -132.765 90.605 -132.435 ;
        RECT 90.275 -134.125 90.605 -133.795 ;
        RECT 90.275 -135.485 90.605 -135.155 ;
        RECT 90.275 -136.845 90.605 -136.515 ;
        RECT 90.275 -138.205 90.605 -137.875 ;
        RECT 90.275 -139.565 90.605 -139.235 ;
        RECT 90.275 -140.925 90.605 -140.595 ;
        RECT 90.275 -142.285 90.605 -141.955 ;
        RECT 90.275 -143.645 90.605 -143.315 ;
        RECT 90.275 -145.005 90.605 -144.675 ;
        RECT 90.275 -146.365 90.605 -146.035 ;
        RECT 90.275 -147.725 90.605 -147.395 ;
        RECT 90.275 -149.085 90.605 -148.755 ;
        RECT 90.275 -150.445 90.605 -150.115 ;
        RECT 90.275 -151.805 90.605 -151.475 ;
        RECT 90.275 -153.165 90.605 -152.835 ;
        RECT 90.275 -154.525 90.605 -154.195 ;
        RECT 90.275 -155.885 90.605 -155.555 ;
        RECT 90.275 -157.245 90.605 -156.915 ;
        RECT 90.275 -158.605 90.605 -158.275 ;
        RECT 90.275 -159.965 90.605 -159.635 ;
        RECT 90.275 -161.325 90.605 -160.995 ;
        RECT 90.275 -162.685 90.605 -162.355 ;
        RECT 90.275 -164.045 90.605 -163.715 ;
        RECT 90.275 -165.405 90.605 -165.075 ;
        RECT 90.275 -166.765 90.605 -166.435 ;
        RECT 90.275 -168.125 90.605 -167.795 ;
        RECT 90.275 -169.485 90.605 -169.155 ;
        RECT 90.275 -170.845 90.605 -170.515 ;
        RECT 90.275 -172.205 90.605 -171.875 ;
        RECT 90.275 -173.565 90.605 -173.235 ;
        RECT 90.275 -174.925 90.605 -174.595 ;
        RECT 90.275 -176.285 90.605 -175.955 ;
        RECT 90.275 -177.645 90.605 -177.315 ;
        RECT 90.275 -183.29 90.605 -182.16 ;
        RECT 90.28 -183.405 90.6 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 91.635 244.04 91.965 245.17 ;
        RECT 91.635 239.875 91.965 240.205 ;
        RECT 91.635 238.515 91.965 238.845 ;
        RECT 91.635 237.155 91.965 237.485 ;
        RECT 91.64 237.155 91.96 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 91.635 -0.845 91.965 -0.515 ;
        RECT 91.635 -2.205 91.965 -1.875 ;
        RECT 91.635 -3.565 91.965 -3.235 ;
        RECT 91.64 -3.565 91.96 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 92.995 244.04 93.325 245.17 ;
        RECT 92.995 239.875 93.325 240.205 ;
        RECT 92.995 238.515 93.325 238.845 ;
        RECT 92.995 237.155 93.325 237.485 ;
        RECT 93 237.155 93.32 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 92.995 -0.845 93.325 -0.515 ;
        RECT 92.995 -2.205 93.325 -1.875 ;
        RECT 92.995 -3.565 93.325 -3.235 ;
        RECT 93 -3.565 93.32 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 92.995 -91.965 93.325 -91.635 ;
        RECT 92.995 -93.325 93.325 -92.995 ;
        RECT 92.995 -94.685 93.325 -94.355 ;
        RECT 92.995 -96.045 93.325 -95.715 ;
        RECT 92.995 -97.405 93.325 -97.075 ;
        RECT 92.995 -98.765 93.325 -98.435 ;
        RECT 92.995 -100.125 93.325 -99.795 ;
        RECT 92.995 -101.485 93.325 -101.155 ;
        RECT 92.995 -102.845 93.325 -102.515 ;
        RECT 92.995 -104.205 93.325 -103.875 ;
        RECT 92.995 -105.565 93.325 -105.235 ;
        RECT 92.995 -106.925 93.325 -106.595 ;
        RECT 92.995 -108.285 93.325 -107.955 ;
        RECT 92.995 -109.645 93.325 -109.315 ;
        RECT 92.995 -111.005 93.325 -110.675 ;
        RECT 92.995 -112.365 93.325 -112.035 ;
        RECT 92.995 -113.725 93.325 -113.395 ;
        RECT 92.995 -115.085 93.325 -114.755 ;
        RECT 92.995 -116.445 93.325 -116.115 ;
        RECT 92.995 -117.805 93.325 -117.475 ;
        RECT 92.995 -119.165 93.325 -118.835 ;
        RECT 92.995 -120.525 93.325 -120.195 ;
        RECT 92.995 -121.885 93.325 -121.555 ;
        RECT 92.995 -123.245 93.325 -122.915 ;
        RECT 92.995 -124.605 93.325 -124.275 ;
        RECT 92.995 -125.965 93.325 -125.635 ;
        RECT 92.995 -127.325 93.325 -126.995 ;
        RECT 92.995 -128.685 93.325 -128.355 ;
        RECT 92.995 -130.045 93.325 -129.715 ;
        RECT 92.995 -131.405 93.325 -131.075 ;
        RECT 92.995 -132.765 93.325 -132.435 ;
        RECT 92.995 -134.125 93.325 -133.795 ;
        RECT 92.995 -135.485 93.325 -135.155 ;
        RECT 92.995 -136.845 93.325 -136.515 ;
        RECT 92.995 -138.205 93.325 -137.875 ;
        RECT 92.995 -139.565 93.325 -139.235 ;
        RECT 92.995 -140.925 93.325 -140.595 ;
        RECT 92.995 -142.285 93.325 -141.955 ;
        RECT 92.995 -143.645 93.325 -143.315 ;
        RECT 92.995 -145.005 93.325 -144.675 ;
        RECT 92.995 -146.365 93.325 -146.035 ;
        RECT 92.995 -147.725 93.325 -147.395 ;
        RECT 92.995 -149.085 93.325 -148.755 ;
        RECT 92.995 -150.445 93.325 -150.115 ;
        RECT 92.995 -151.805 93.325 -151.475 ;
        RECT 92.995 -153.165 93.325 -152.835 ;
        RECT 92.995 -154.525 93.325 -154.195 ;
        RECT 92.995 -155.885 93.325 -155.555 ;
        RECT 92.995 -157.245 93.325 -156.915 ;
        RECT 92.995 -158.605 93.325 -158.275 ;
        RECT 92.995 -159.965 93.325 -159.635 ;
        RECT 92.995 -161.325 93.325 -160.995 ;
        RECT 92.995 -162.685 93.325 -162.355 ;
        RECT 92.995 -164.045 93.325 -163.715 ;
        RECT 92.995 -165.405 93.325 -165.075 ;
        RECT 92.995 -166.765 93.325 -166.435 ;
        RECT 92.995 -168.125 93.325 -167.795 ;
        RECT 92.995 -169.485 93.325 -169.155 ;
        RECT 92.995 -170.845 93.325 -170.515 ;
        RECT 92.995 -172.205 93.325 -171.875 ;
        RECT 92.995 -173.565 93.325 -173.235 ;
        RECT 92.995 -174.925 93.325 -174.595 ;
        RECT 92.995 -176.285 93.325 -175.955 ;
        RECT 92.995 -177.645 93.325 -177.315 ;
        RECT 92.995 -183.29 93.325 -182.16 ;
        RECT 93 -183.405 93.32 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 94.16 -94.075 94.49 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 94.355 244.04 94.685 245.17 ;
        RECT 94.355 239.875 94.685 240.205 ;
        RECT 94.355 238.515 94.685 238.845 ;
        RECT 94.355 237.155 94.685 237.485 ;
        RECT 94.36 237.155 94.68 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 94.355 -96.045 94.685 -95.715 ;
        RECT 94.355 -97.405 94.685 -97.075 ;
        RECT 94.355 -98.765 94.685 -98.435 ;
        RECT 94.355 -100.125 94.685 -99.795 ;
        RECT 94.355 -101.485 94.685 -101.155 ;
        RECT 94.355 -102.845 94.685 -102.515 ;
        RECT 94.355 -104.205 94.685 -103.875 ;
        RECT 94.355 -105.565 94.685 -105.235 ;
        RECT 94.355 -106.925 94.685 -106.595 ;
        RECT 94.355 -108.285 94.685 -107.955 ;
        RECT 94.355 -109.645 94.685 -109.315 ;
        RECT 94.355 -111.005 94.685 -110.675 ;
        RECT 94.355 -112.365 94.685 -112.035 ;
        RECT 94.355 -113.725 94.685 -113.395 ;
        RECT 94.355 -115.085 94.685 -114.755 ;
        RECT 94.355 -116.445 94.685 -116.115 ;
        RECT 94.355 -117.805 94.685 -117.475 ;
        RECT 94.355 -119.165 94.685 -118.835 ;
        RECT 94.355 -120.525 94.685 -120.195 ;
        RECT 94.355 -121.885 94.685 -121.555 ;
        RECT 94.355 -123.245 94.685 -122.915 ;
        RECT 94.355 -124.605 94.685 -124.275 ;
        RECT 94.355 -125.965 94.685 -125.635 ;
        RECT 94.355 -127.325 94.685 -126.995 ;
        RECT 94.355 -128.685 94.685 -128.355 ;
        RECT 94.355 -130.045 94.685 -129.715 ;
        RECT 94.355 -131.405 94.685 -131.075 ;
        RECT 94.355 -132.765 94.685 -132.435 ;
        RECT 94.355 -134.125 94.685 -133.795 ;
        RECT 94.355 -135.485 94.685 -135.155 ;
        RECT 94.355 -136.845 94.685 -136.515 ;
        RECT 94.355 -138.205 94.685 -137.875 ;
        RECT 94.355 -139.565 94.685 -139.235 ;
        RECT 94.355 -140.925 94.685 -140.595 ;
        RECT 94.355 -142.285 94.685 -141.955 ;
        RECT 94.355 -143.645 94.685 -143.315 ;
        RECT 94.355 -145.005 94.685 -144.675 ;
        RECT 94.355 -146.365 94.685 -146.035 ;
        RECT 94.355 -147.725 94.685 -147.395 ;
        RECT 94.355 -149.085 94.685 -148.755 ;
        RECT 94.355 -150.445 94.685 -150.115 ;
        RECT 94.355 -151.805 94.685 -151.475 ;
        RECT 94.355 -153.165 94.685 -152.835 ;
        RECT 94.355 -154.525 94.685 -154.195 ;
        RECT 94.355 -155.885 94.685 -155.555 ;
        RECT 94.355 -157.245 94.685 -156.915 ;
        RECT 94.355 -158.605 94.685 -158.275 ;
        RECT 94.355 -159.965 94.685 -159.635 ;
        RECT 94.355 -161.325 94.685 -160.995 ;
        RECT 94.355 -162.685 94.685 -162.355 ;
        RECT 94.355 -164.045 94.685 -163.715 ;
        RECT 94.355 -165.405 94.685 -165.075 ;
        RECT 94.355 -166.765 94.685 -166.435 ;
        RECT 94.355 -168.125 94.685 -167.795 ;
        RECT 94.355 -169.485 94.685 -169.155 ;
        RECT 94.355 -170.845 94.685 -170.515 ;
        RECT 94.355 -172.205 94.685 -171.875 ;
        RECT 94.355 -173.565 94.685 -173.235 ;
        RECT 94.355 -174.925 94.685 -174.595 ;
        RECT 94.355 -176.285 94.685 -175.955 ;
        RECT 94.355 -177.645 94.685 -177.315 ;
        RECT 94.355 -183.29 94.685 -182.16 ;
        RECT 94.36 -183.405 94.68 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 95.715 244.04 96.045 245.17 ;
        RECT 95.715 239.875 96.045 240.205 ;
        RECT 95.715 238.515 96.045 238.845 ;
        RECT 95.715 237.155 96.045 237.485 ;
        RECT 95.72 237.155 96.04 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 95.715 -0.845 96.045 -0.515 ;
        RECT 95.715 -2.205 96.045 -1.875 ;
        RECT 95.715 -3.565 96.045 -3.235 ;
        RECT 95.72 -3.565 96.04 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 97.075 244.04 97.405 245.17 ;
        RECT 97.075 239.875 97.405 240.205 ;
        RECT 97.075 238.515 97.405 238.845 ;
        RECT 97.075 237.155 97.405 237.485 ;
        RECT 97.08 237.155 97.4 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 97.075 -0.845 97.405 -0.515 ;
        RECT 97.075 -2.205 97.405 -1.875 ;
        RECT 97.075 -3.565 97.405 -3.235 ;
        RECT 97.08 -3.565 97.4 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 98.435 244.04 98.765 245.17 ;
        RECT 98.435 239.875 98.765 240.205 ;
        RECT 98.435 238.515 98.765 238.845 ;
        RECT 98.435 237.155 98.765 237.485 ;
        RECT 98.44 237.155 98.76 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 98.435 -0.845 98.765 -0.515 ;
        RECT 98.435 -2.205 98.765 -1.875 ;
        RECT 98.435 -3.565 98.765 -3.235 ;
        RECT 98.44 -3.565 98.76 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 98.435 -91.965 98.765 -91.635 ;
        RECT 98.435 -93.325 98.765 -92.995 ;
        RECT 98.435 -94.685 98.765 -94.355 ;
        RECT 98.435 -96.045 98.765 -95.715 ;
        RECT 98.435 -97.405 98.765 -97.075 ;
        RECT 98.435 -98.765 98.765 -98.435 ;
        RECT 98.435 -100.125 98.765 -99.795 ;
        RECT 98.435 -101.485 98.765 -101.155 ;
        RECT 98.435 -102.845 98.765 -102.515 ;
        RECT 98.435 -104.205 98.765 -103.875 ;
        RECT 98.435 -105.565 98.765 -105.235 ;
        RECT 98.435 -106.925 98.765 -106.595 ;
        RECT 98.435 -108.285 98.765 -107.955 ;
        RECT 98.435 -109.645 98.765 -109.315 ;
        RECT 98.435 -111.005 98.765 -110.675 ;
        RECT 98.435 -112.365 98.765 -112.035 ;
        RECT 98.435 -113.725 98.765 -113.395 ;
        RECT 98.435 -115.085 98.765 -114.755 ;
        RECT 98.435 -116.445 98.765 -116.115 ;
        RECT 98.435 -117.805 98.765 -117.475 ;
        RECT 98.435 -119.165 98.765 -118.835 ;
        RECT 98.435 -120.525 98.765 -120.195 ;
        RECT 98.435 -121.885 98.765 -121.555 ;
        RECT 98.435 -123.245 98.765 -122.915 ;
        RECT 98.435 -124.605 98.765 -124.275 ;
        RECT 98.435 -125.965 98.765 -125.635 ;
        RECT 98.435 -127.325 98.765 -126.995 ;
        RECT 98.435 -128.685 98.765 -128.355 ;
        RECT 98.435 -130.045 98.765 -129.715 ;
        RECT 98.435 -131.405 98.765 -131.075 ;
        RECT 98.435 -132.765 98.765 -132.435 ;
        RECT 98.435 -134.125 98.765 -133.795 ;
        RECT 98.435 -135.485 98.765 -135.155 ;
        RECT 98.435 -136.845 98.765 -136.515 ;
        RECT 98.435 -138.205 98.765 -137.875 ;
        RECT 98.435 -139.565 98.765 -139.235 ;
        RECT 98.435 -140.925 98.765 -140.595 ;
        RECT 98.435 -142.285 98.765 -141.955 ;
        RECT 98.435 -143.645 98.765 -143.315 ;
        RECT 98.435 -145.005 98.765 -144.675 ;
        RECT 98.435 -146.365 98.765 -146.035 ;
        RECT 98.435 -147.725 98.765 -147.395 ;
        RECT 98.435 -149.085 98.765 -148.755 ;
        RECT 98.435 -150.445 98.765 -150.115 ;
        RECT 98.435 -151.805 98.765 -151.475 ;
        RECT 98.435 -153.165 98.765 -152.835 ;
        RECT 98.435 -154.525 98.765 -154.195 ;
        RECT 98.435 -155.885 98.765 -155.555 ;
        RECT 98.435 -157.245 98.765 -156.915 ;
        RECT 98.435 -158.605 98.765 -158.275 ;
        RECT 98.435 -159.965 98.765 -159.635 ;
        RECT 98.435 -161.325 98.765 -160.995 ;
        RECT 98.435 -162.685 98.765 -162.355 ;
        RECT 98.435 -164.045 98.765 -163.715 ;
        RECT 98.435 -165.405 98.765 -165.075 ;
        RECT 98.435 -166.765 98.765 -166.435 ;
        RECT 98.435 -168.125 98.765 -167.795 ;
        RECT 98.435 -169.485 98.765 -169.155 ;
        RECT 98.435 -170.845 98.765 -170.515 ;
        RECT 98.435 -172.205 98.765 -171.875 ;
        RECT 98.435 -173.565 98.765 -173.235 ;
        RECT 98.435 -174.925 98.765 -174.595 ;
        RECT 98.435 -176.285 98.765 -175.955 ;
        RECT 98.435 -177.645 98.765 -177.315 ;
        RECT 98.435 -183.29 98.765 -182.16 ;
        RECT 98.44 -183.405 98.76 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 99.795 244.04 100.125 245.17 ;
        RECT 99.795 239.875 100.125 240.205 ;
        RECT 99.795 238.515 100.125 238.845 ;
        RECT 99.795 237.155 100.125 237.485 ;
        RECT 99.8 237.155 100.12 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 99.795 -96.045 100.125 -95.715 ;
        RECT 99.795 -97.405 100.125 -97.075 ;
        RECT 99.795 -98.765 100.125 -98.435 ;
        RECT 99.795 -100.125 100.125 -99.795 ;
        RECT 99.795 -101.485 100.125 -101.155 ;
        RECT 99.795 -102.845 100.125 -102.515 ;
        RECT 99.795 -104.205 100.125 -103.875 ;
        RECT 99.795 -105.565 100.125 -105.235 ;
        RECT 99.795 -106.925 100.125 -106.595 ;
        RECT 99.795 -108.285 100.125 -107.955 ;
        RECT 99.795 -109.645 100.125 -109.315 ;
        RECT 99.795 -111.005 100.125 -110.675 ;
        RECT 99.795 -112.365 100.125 -112.035 ;
        RECT 99.795 -113.725 100.125 -113.395 ;
        RECT 99.795 -115.085 100.125 -114.755 ;
        RECT 99.795 -116.445 100.125 -116.115 ;
        RECT 99.795 -117.805 100.125 -117.475 ;
        RECT 99.795 -119.165 100.125 -118.835 ;
        RECT 99.795 -120.525 100.125 -120.195 ;
        RECT 99.795 -121.885 100.125 -121.555 ;
        RECT 99.795 -123.245 100.125 -122.915 ;
        RECT 99.795 -124.605 100.125 -124.275 ;
        RECT 99.795 -125.965 100.125 -125.635 ;
        RECT 99.795 -127.325 100.125 -126.995 ;
        RECT 99.795 -128.685 100.125 -128.355 ;
        RECT 99.795 -130.045 100.125 -129.715 ;
        RECT 99.795 -131.405 100.125 -131.075 ;
        RECT 99.795 -132.765 100.125 -132.435 ;
        RECT 99.795 -134.125 100.125 -133.795 ;
        RECT 99.795 -135.485 100.125 -135.155 ;
        RECT 99.795 -136.845 100.125 -136.515 ;
        RECT 99.795 -138.205 100.125 -137.875 ;
        RECT 99.795 -139.565 100.125 -139.235 ;
        RECT 99.795 -140.925 100.125 -140.595 ;
        RECT 99.795 -142.285 100.125 -141.955 ;
        RECT 99.795 -143.645 100.125 -143.315 ;
        RECT 99.795 -145.005 100.125 -144.675 ;
        RECT 99.795 -146.365 100.125 -146.035 ;
        RECT 99.795 -147.725 100.125 -147.395 ;
        RECT 99.795 -149.085 100.125 -148.755 ;
        RECT 99.795 -150.445 100.125 -150.115 ;
        RECT 99.795 -151.805 100.125 -151.475 ;
        RECT 99.795 -153.165 100.125 -152.835 ;
        RECT 99.795 -154.525 100.125 -154.195 ;
        RECT 99.795 -155.885 100.125 -155.555 ;
        RECT 99.795 -157.245 100.125 -156.915 ;
        RECT 99.795 -158.605 100.125 -158.275 ;
        RECT 99.795 -159.965 100.125 -159.635 ;
        RECT 99.795 -161.325 100.125 -160.995 ;
        RECT 99.795 -162.685 100.125 -162.355 ;
        RECT 99.795 -164.045 100.125 -163.715 ;
        RECT 99.795 -165.405 100.125 -165.075 ;
        RECT 99.795 -166.765 100.125 -166.435 ;
        RECT 99.795 -168.125 100.125 -167.795 ;
        RECT 99.795 -169.485 100.125 -169.155 ;
        RECT 99.795 -170.845 100.125 -170.515 ;
        RECT 99.795 -172.205 100.125 -171.875 ;
        RECT 99.795 -173.565 100.125 -173.235 ;
        RECT 99.795 -174.925 100.125 -174.595 ;
        RECT 99.795 -176.285 100.125 -175.955 ;
        RECT 99.795 -177.645 100.125 -177.315 ;
        RECT 99.795 -183.29 100.125 -182.16 ;
        RECT 99.8 -183.405 100.12 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 100.26 -94.075 100.59 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 101.155 244.04 101.485 245.17 ;
        RECT 101.155 239.875 101.485 240.205 ;
        RECT 101.155 238.515 101.485 238.845 ;
        RECT 101.155 237.155 101.485 237.485 ;
        RECT 101.16 237.155 101.48 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 102.515 244.04 102.845 245.17 ;
        RECT 102.515 239.875 102.845 240.205 ;
        RECT 102.515 238.515 102.845 238.845 ;
        RECT 102.515 237.155 102.845 237.485 ;
        RECT 102.52 237.155 102.84 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 102.515 -0.845 102.845 -0.515 ;
        RECT 102.515 -2.205 102.845 -1.875 ;
        RECT 102.515 -3.565 102.845 -3.235 ;
        RECT 102.52 -3.565 102.84 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 102.515 -91.965 102.845 -91.635 ;
        RECT 102.515 -93.325 102.845 -92.995 ;
        RECT 102.515 -94.685 102.845 -94.355 ;
        RECT 102.515 -96.045 102.845 -95.715 ;
        RECT 102.515 -97.405 102.845 -97.075 ;
        RECT 102.515 -98.765 102.845 -98.435 ;
        RECT 102.515 -100.125 102.845 -99.795 ;
        RECT 102.515 -101.485 102.845 -101.155 ;
        RECT 102.515 -102.845 102.845 -102.515 ;
        RECT 102.515 -104.205 102.845 -103.875 ;
        RECT 102.515 -105.565 102.845 -105.235 ;
        RECT 102.515 -106.925 102.845 -106.595 ;
        RECT 102.515 -108.285 102.845 -107.955 ;
        RECT 102.515 -109.645 102.845 -109.315 ;
        RECT 102.515 -111.005 102.845 -110.675 ;
        RECT 102.515 -112.365 102.845 -112.035 ;
        RECT 102.515 -113.725 102.845 -113.395 ;
        RECT 102.515 -115.085 102.845 -114.755 ;
        RECT 102.515 -116.445 102.845 -116.115 ;
        RECT 102.515 -117.805 102.845 -117.475 ;
        RECT 102.515 -119.165 102.845 -118.835 ;
        RECT 102.515 -120.525 102.845 -120.195 ;
        RECT 102.515 -121.885 102.845 -121.555 ;
        RECT 102.515 -123.245 102.845 -122.915 ;
        RECT 102.515 -124.605 102.845 -124.275 ;
        RECT 102.515 -125.965 102.845 -125.635 ;
        RECT 102.515 -127.325 102.845 -126.995 ;
        RECT 102.515 -128.685 102.845 -128.355 ;
        RECT 102.515 -130.045 102.845 -129.715 ;
        RECT 102.515 -131.405 102.845 -131.075 ;
        RECT 102.515 -132.765 102.845 -132.435 ;
        RECT 102.515 -134.125 102.845 -133.795 ;
        RECT 102.515 -135.485 102.845 -135.155 ;
        RECT 102.515 -136.845 102.845 -136.515 ;
        RECT 102.515 -138.205 102.845 -137.875 ;
        RECT 102.515 -139.565 102.845 -139.235 ;
        RECT 102.515 -140.925 102.845 -140.595 ;
        RECT 102.515 -142.285 102.845 -141.955 ;
        RECT 102.515 -143.645 102.845 -143.315 ;
        RECT 102.515 -145.005 102.845 -144.675 ;
        RECT 102.515 -146.365 102.845 -146.035 ;
        RECT 102.515 -147.725 102.845 -147.395 ;
        RECT 102.515 -149.085 102.845 -148.755 ;
        RECT 102.515 -150.445 102.845 -150.115 ;
        RECT 102.515 -151.805 102.845 -151.475 ;
        RECT 102.515 -153.165 102.845 -152.835 ;
        RECT 102.515 -154.525 102.845 -154.195 ;
        RECT 102.515 -155.885 102.845 -155.555 ;
        RECT 102.515 -157.245 102.845 -156.915 ;
        RECT 102.515 -158.605 102.845 -158.275 ;
        RECT 102.515 -159.965 102.845 -159.635 ;
        RECT 102.515 -161.325 102.845 -160.995 ;
        RECT 102.515 -162.685 102.845 -162.355 ;
        RECT 102.515 -164.045 102.845 -163.715 ;
        RECT 102.515 -165.405 102.845 -165.075 ;
        RECT 102.515 -166.765 102.845 -166.435 ;
        RECT 102.515 -168.125 102.845 -167.795 ;
        RECT 102.515 -169.485 102.845 -169.155 ;
        RECT 102.515 -170.845 102.845 -170.515 ;
        RECT 102.515 -172.205 102.845 -171.875 ;
        RECT 102.515 -173.565 102.845 -173.235 ;
        RECT 102.515 -174.925 102.845 -174.595 ;
        RECT 102.515 -176.285 102.845 -175.955 ;
        RECT 102.515 -177.645 102.845 -177.315 ;
        RECT 102.515 -183.29 102.845 -182.16 ;
        RECT 102.52 -183.405 102.84 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 103.875 244.04 104.205 245.17 ;
        RECT 103.875 239.875 104.205 240.205 ;
        RECT 103.875 238.515 104.205 238.845 ;
        RECT 103.875 237.155 104.205 237.485 ;
        RECT 103.88 237.155 104.2 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 103.875 -0.845 104.205 -0.515 ;
        RECT 103.875 -2.205 104.205 -1.875 ;
        RECT 103.875 -3.565 104.205 -3.235 ;
        RECT 103.88 -3.565 104.2 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 105.235 244.04 105.565 245.17 ;
        RECT 105.235 239.875 105.565 240.205 ;
        RECT 105.235 238.515 105.565 238.845 ;
        RECT 105.235 237.155 105.565 237.485 ;
        RECT 105.24 237.155 105.56 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 105.235 -0.845 105.565 -0.515 ;
        RECT 105.235 -2.205 105.565 -1.875 ;
        RECT 105.235 -3.565 105.565 -3.235 ;
        RECT 105.24 -3.565 105.56 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 105.235 -150.445 105.565 -150.115 ;
        RECT 105.235 -151.805 105.565 -151.475 ;
        RECT 105.235 -153.165 105.565 -152.835 ;
        RECT 105.235 -154.525 105.565 -154.195 ;
        RECT 105.235 -155.885 105.565 -155.555 ;
        RECT 105.235 -157.245 105.565 -156.915 ;
        RECT 105.235 -158.605 105.565 -158.275 ;
        RECT 105.235 -159.965 105.565 -159.635 ;
        RECT 105.235 -161.325 105.565 -160.995 ;
        RECT 105.235 -162.685 105.565 -162.355 ;
        RECT 105.235 -164.045 105.565 -163.715 ;
        RECT 105.235 -165.405 105.565 -165.075 ;
        RECT 105.235 -166.765 105.565 -166.435 ;
        RECT 105.235 -168.125 105.565 -167.795 ;
        RECT 105.235 -169.485 105.565 -169.155 ;
        RECT 105.235 -170.845 105.565 -170.515 ;
        RECT 105.235 -172.205 105.565 -171.875 ;
        RECT 105.235 -173.565 105.565 -173.235 ;
        RECT 105.235 -174.925 105.565 -174.595 ;
        RECT 105.235 -176.285 105.565 -175.955 ;
        RECT 105.235 -177.645 105.565 -177.315 ;
        RECT 105.235 -183.29 105.565 -182.16 ;
        RECT 105.24 -183.405 105.56 -90.96 ;
        RECT 105.235 -91.965 105.565 -91.635 ;
        RECT 105.235 -93.325 105.565 -92.995 ;
        RECT 105.235 -94.685 105.565 -94.355 ;
        RECT 105.235 -96.045 105.565 -95.715 ;
        RECT 105.235 -97.405 105.565 -97.075 ;
        RECT 105.235 -98.765 105.565 -98.435 ;
        RECT 105.235 -100.125 105.565 -99.795 ;
        RECT 105.235 -101.485 105.565 -101.155 ;
        RECT 105.235 -102.845 105.565 -102.515 ;
        RECT 105.235 -104.205 105.565 -103.875 ;
        RECT 105.235 -105.565 105.565 -105.235 ;
        RECT 105.235 -106.925 105.565 -106.595 ;
        RECT 105.235 -108.285 105.565 -107.955 ;
        RECT 105.235 -109.645 105.565 -109.315 ;
        RECT 105.235 -111.005 105.565 -110.675 ;
        RECT 105.235 -112.365 105.565 -112.035 ;
        RECT 105.235 -113.725 105.565 -113.395 ;
        RECT 105.235 -115.085 105.565 -114.755 ;
        RECT 105.235 -116.445 105.565 -116.115 ;
        RECT 105.235 -117.805 105.565 -117.475 ;
        RECT 105.235 -119.165 105.565 -118.835 ;
        RECT 105.235 -120.525 105.565 -120.195 ;
        RECT 105.235 -121.885 105.565 -121.555 ;
        RECT 105.235 -123.245 105.565 -122.915 ;
        RECT 105.235 -124.605 105.565 -124.275 ;
        RECT 105.235 -125.965 105.565 -125.635 ;
        RECT 105.235 -127.325 105.565 -126.995 ;
        RECT 105.235 -128.685 105.565 -128.355 ;
        RECT 105.235 -130.045 105.565 -129.715 ;
        RECT 105.235 -131.405 105.565 -131.075 ;
        RECT 105.235 -132.765 105.565 -132.435 ;
        RECT 105.235 -134.125 105.565 -133.795 ;
        RECT 105.235 -135.485 105.565 -135.155 ;
        RECT 105.235 -136.845 105.565 -136.515 ;
        RECT 105.235 -138.205 105.565 -137.875 ;
        RECT 105.235 -139.565 105.565 -139.235 ;
        RECT 105.235 -140.925 105.565 -140.595 ;
        RECT 105.235 -142.285 105.565 -141.955 ;
        RECT 105.235 -143.645 105.565 -143.315 ;
        RECT 105.235 -145.005 105.565 -144.675 ;
        RECT 105.235 -146.365 105.565 -146.035 ;
        RECT 105.235 -147.725 105.565 -147.395 ;
        RECT 105.235 -149.085 105.565 -148.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.035 -91.965 44.365 -91.635 ;
        RECT 44.035 -93.325 44.365 -92.995 ;
        RECT 44.035 -94.685 44.365 -94.355 ;
        RECT 44.035 -96.045 44.365 -95.715 ;
        RECT 44.035 -97.405 44.365 -97.075 ;
        RECT 44.035 -98.765 44.365 -98.435 ;
        RECT 44.035 -100.125 44.365 -99.795 ;
        RECT 44.035 -101.485 44.365 -101.155 ;
        RECT 44.035 -102.845 44.365 -102.515 ;
        RECT 44.035 -104.205 44.365 -103.875 ;
        RECT 44.035 -105.565 44.365 -105.235 ;
        RECT 44.035 -106.925 44.365 -106.595 ;
        RECT 44.035 -108.285 44.365 -107.955 ;
        RECT 44.035 -109.645 44.365 -109.315 ;
        RECT 44.035 -111.005 44.365 -110.675 ;
        RECT 44.035 -112.365 44.365 -112.035 ;
        RECT 44.035 -113.725 44.365 -113.395 ;
        RECT 44.035 -115.085 44.365 -114.755 ;
        RECT 44.035 -116.445 44.365 -116.115 ;
        RECT 44.035 -117.805 44.365 -117.475 ;
        RECT 44.035 -119.165 44.365 -118.835 ;
        RECT 44.035 -120.525 44.365 -120.195 ;
        RECT 44.035 -121.885 44.365 -121.555 ;
        RECT 44.035 -123.245 44.365 -122.915 ;
        RECT 44.035 -124.605 44.365 -124.275 ;
        RECT 44.035 -125.965 44.365 -125.635 ;
        RECT 44.035 -127.325 44.365 -126.995 ;
        RECT 44.035 -128.685 44.365 -128.355 ;
        RECT 44.035 -130.045 44.365 -129.715 ;
        RECT 44.035 -131.405 44.365 -131.075 ;
        RECT 44.035 -132.765 44.365 -132.435 ;
        RECT 44.035 -134.125 44.365 -133.795 ;
        RECT 44.035 -135.485 44.365 -135.155 ;
        RECT 44.035 -136.845 44.365 -136.515 ;
        RECT 44.035 -138.205 44.365 -137.875 ;
        RECT 44.035 -139.565 44.365 -139.235 ;
        RECT 44.035 -140.925 44.365 -140.595 ;
        RECT 44.035 -142.285 44.365 -141.955 ;
        RECT 44.035 -143.645 44.365 -143.315 ;
        RECT 44.035 -145.005 44.365 -144.675 ;
        RECT 44.035 -146.365 44.365 -146.035 ;
        RECT 44.035 -147.725 44.365 -147.395 ;
        RECT 44.035 -149.085 44.365 -148.755 ;
        RECT 44.035 -150.445 44.365 -150.115 ;
        RECT 44.035 -151.805 44.365 -151.475 ;
        RECT 44.035 -153.165 44.365 -152.835 ;
        RECT 44.035 -154.525 44.365 -154.195 ;
        RECT 44.035 -155.885 44.365 -155.555 ;
        RECT 44.035 -157.245 44.365 -156.915 ;
        RECT 44.035 -158.605 44.365 -158.275 ;
        RECT 44.035 -159.965 44.365 -159.635 ;
        RECT 44.035 -161.325 44.365 -160.995 ;
        RECT 44.035 -162.685 44.365 -162.355 ;
        RECT 44.035 -164.045 44.365 -163.715 ;
        RECT 44.035 -165.405 44.365 -165.075 ;
        RECT 44.035 -166.765 44.365 -166.435 ;
        RECT 44.035 -168.125 44.365 -167.795 ;
        RECT 44.035 -169.485 44.365 -169.155 ;
        RECT 44.035 -170.845 44.365 -170.515 ;
        RECT 44.035 -172.205 44.365 -171.875 ;
        RECT 44.035 -173.565 44.365 -173.235 ;
        RECT 44.035 -174.925 44.365 -174.595 ;
        RECT 44.035 -176.285 44.365 -175.955 ;
        RECT 44.035 -177.645 44.365 -177.315 ;
        RECT 44.035 -183.29 44.365 -182.16 ;
        RECT 44.04 -183.405 44.36 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.36 -94.075 45.69 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.395 244.04 45.725 245.17 ;
        RECT 45.395 239.875 45.725 240.205 ;
        RECT 45.395 238.515 45.725 238.845 ;
        RECT 45.395 237.155 45.725 237.485 ;
        RECT 45.4 237.155 45.72 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.395 -96.045 45.725 -95.715 ;
        RECT 45.395 -97.405 45.725 -97.075 ;
        RECT 45.395 -98.765 45.725 -98.435 ;
        RECT 45.395 -100.125 45.725 -99.795 ;
        RECT 45.395 -101.485 45.725 -101.155 ;
        RECT 45.395 -102.845 45.725 -102.515 ;
        RECT 45.395 -104.205 45.725 -103.875 ;
        RECT 45.395 -105.565 45.725 -105.235 ;
        RECT 45.395 -106.925 45.725 -106.595 ;
        RECT 45.395 -108.285 45.725 -107.955 ;
        RECT 45.395 -109.645 45.725 -109.315 ;
        RECT 45.395 -111.005 45.725 -110.675 ;
        RECT 45.395 -112.365 45.725 -112.035 ;
        RECT 45.395 -113.725 45.725 -113.395 ;
        RECT 45.395 -115.085 45.725 -114.755 ;
        RECT 45.395 -116.445 45.725 -116.115 ;
        RECT 45.395 -117.805 45.725 -117.475 ;
        RECT 45.395 -119.165 45.725 -118.835 ;
        RECT 45.395 -120.525 45.725 -120.195 ;
        RECT 45.395 -121.885 45.725 -121.555 ;
        RECT 45.395 -123.245 45.725 -122.915 ;
        RECT 45.395 -124.605 45.725 -124.275 ;
        RECT 45.395 -125.965 45.725 -125.635 ;
        RECT 45.395 -127.325 45.725 -126.995 ;
        RECT 45.395 -128.685 45.725 -128.355 ;
        RECT 45.395 -130.045 45.725 -129.715 ;
        RECT 45.395 -131.405 45.725 -131.075 ;
        RECT 45.395 -132.765 45.725 -132.435 ;
        RECT 45.395 -134.125 45.725 -133.795 ;
        RECT 45.395 -135.485 45.725 -135.155 ;
        RECT 45.395 -136.845 45.725 -136.515 ;
        RECT 45.395 -138.205 45.725 -137.875 ;
        RECT 45.395 -139.565 45.725 -139.235 ;
        RECT 45.395 -140.925 45.725 -140.595 ;
        RECT 45.395 -142.285 45.725 -141.955 ;
        RECT 45.395 -143.645 45.725 -143.315 ;
        RECT 45.395 -145.005 45.725 -144.675 ;
        RECT 45.395 -146.365 45.725 -146.035 ;
        RECT 45.395 -147.725 45.725 -147.395 ;
        RECT 45.395 -149.085 45.725 -148.755 ;
        RECT 45.395 -150.445 45.725 -150.115 ;
        RECT 45.395 -151.805 45.725 -151.475 ;
        RECT 45.395 -153.165 45.725 -152.835 ;
        RECT 45.395 -154.525 45.725 -154.195 ;
        RECT 45.395 -155.885 45.725 -155.555 ;
        RECT 45.395 -157.245 45.725 -156.915 ;
        RECT 45.395 -158.605 45.725 -158.275 ;
        RECT 45.395 -159.965 45.725 -159.635 ;
        RECT 45.395 -161.325 45.725 -160.995 ;
        RECT 45.395 -162.685 45.725 -162.355 ;
        RECT 45.395 -164.045 45.725 -163.715 ;
        RECT 45.395 -165.405 45.725 -165.075 ;
        RECT 45.395 -166.765 45.725 -166.435 ;
        RECT 45.395 -168.125 45.725 -167.795 ;
        RECT 45.395 -169.485 45.725 -169.155 ;
        RECT 45.395 -170.845 45.725 -170.515 ;
        RECT 45.395 -172.205 45.725 -171.875 ;
        RECT 45.395 -173.565 45.725 -173.235 ;
        RECT 45.395 -174.925 45.725 -174.595 ;
        RECT 45.395 -176.285 45.725 -175.955 ;
        RECT 45.395 -177.645 45.725 -177.315 ;
        RECT 45.395 -183.29 45.725 -182.16 ;
        RECT 45.4 -183.405 45.72 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.755 244.04 47.085 245.17 ;
        RECT 46.755 239.875 47.085 240.205 ;
        RECT 46.755 238.515 47.085 238.845 ;
        RECT 46.755 237.155 47.085 237.485 ;
        RECT 46.76 237.155 47.08 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.755 -0.845 47.085 -0.515 ;
        RECT 46.755 -2.205 47.085 -1.875 ;
        RECT 46.755 -3.565 47.085 -3.235 ;
        RECT 46.76 -3.565 47.08 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.115 244.04 48.445 245.17 ;
        RECT 48.115 239.875 48.445 240.205 ;
        RECT 48.115 238.515 48.445 238.845 ;
        RECT 48.115 237.155 48.445 237.485 ;
        RECT 48.12 237.155 48.44 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.115 -0.845 48.445 -0.515 ;
        RECT 48.115 -2.205 48.445 -1.875 ;
        RECT 48.115 -3.565 48.445 -3.235 ;
        RECT 48.12 -3.565 48.44 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.475 244.04 49.805 245.17 ;
        RECT 49.475 239.875 49.805 240.205 ;
        RECT 49.475 238.515 49.805 238.845 ;
        RECT 49.475 237.155 49.805 237.485 ;
        RECT 49.48 237.155 49.8 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.475 -0.845 49.805 -0.515 ;
        RECT 49.475 -2.205 49.805 -1.875 ;
        RECT 49.475 -3.565 49.805 -3.235 ;
        RECT 49.48 -3.565 49.8 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.475 -91.965 49.805 -91.635 ;
        RECT 49.475 -93.325 49.805 -92.995 ;
        RECT 49.475 -94.685 49.805 -94.355 ;
        RECT 49.475 -96.045 49.805 -95.715 ;
        RECT 49.475 -97.405 49.805 -97.075 ;
        RECT 49.475 -98.765 49.805 -98.435 ;
        RECT 49.475 -100.125 49.805 -99.795 ;
        RECT 49.475 -101.485 49.805 -101.155 ;
        RECT 49.475 -102.845 49.805 -102.515 ;
        RECT 49.475 -104.205 49.805 -103.875 ;
        RECT 49.475 -105.565 49.805 -105.235 ;
        RECT 49.475 -106.925 49.805 -106.595 ;
        RECT 49.475 -108.285 49.805 -107.955 ;
        RECT 49.475 -109.645 49.805 -109.315 ;
        RECT 49.475 -111.005 49.805 -110.675 ;
        RECT 49.475 -112.365 49.805 -112.035 ;
        RECT 49.475 -113.725 49.805 -113.395 ;
        RECT 49.475 -115.085 49.805 -114.755 ;
        RECT 49.475 -116.445 49.805 -116.115 ;
        RECT 49.475 -117.805 49.805 -117.475 ;
        RECT 49.475 -119.165 49.805 -118.835 ;
        RECT 49.475 -120.525 49.805 -120.195 ;
        RECT 49.475 -121.885 49.805 -121.555 ;
        RECT 49.475 -123.245 49.805 -122.915 ;
        RECT 49.475 -124.605 49.805 -124.275 ;
        RECT 49.475 -125.965 49.805 -125.635 ;
        RECT 49.475 -127.325 49.805 -126.995 ;
        RECT 49.475 -128.685 49.805 -128.355 ;
        RECT 49.475 -130.045 49.805 -129.715 ;
        RECT 49.475 -131.405 49.805 -131.075 ;
        RECT 49.475 -132.765 49.805 -132.435 ;
        RECT 49.475 -134.125 49.805 -133.795 ;
        RECT 49.475 -135.485 49.805 -135.155 ;
        RECT 49.475 -136.845 49.805 -136.515 ;
        RECT 49.475 -138.205 49.805 -137.875 ;
        RECT 49.475 -139.565 49.805 -139.235 ;
        RECT 49.475 -140.925 49.805 -140.595 ;
        RECT 49.475 -142.285 49.805 -141.955 ;
        RECT 49.475 -143.645 49.805 -143.315 ;
        RECT 49.475 -145.005 49.805 -144.675 ;
        RECT 49.475 -146.365 49.805 -146.035 ;
        RECT 49.475 -147.725 49.805 -147.395 ;
        RECT 49.475 -149.085 49.805 -148.755 ;
        RECT 49.475 -150.445 49.805 -150.115 ;
        RECT 49.475 -151.805 49.805 -151.475 ;
        RECT 49.475 -153.165 49.805 -152.835 ;
        RECT 49.475 -154.525 49.805 -154.195 ;
        RECT 49.475 -155.885 49.805 -155.555 ;
        RECT 49.475 -157.245 49.805 -156.915 ;
        RECT 49.475 -158.605 49.805 -158.275 ;
        RECT 49.475 -159.965 49.805 -159.635 ;
        RECT 49.475 -161.325 49.805 -160.995 ;
        RECT 49.475 -162.685 49.805 -162.355 ;
        RECT 49.475 -164.045 49.805 -163.715 ;
        RECT 49.475 -165.405 49.805 -165.075 ;
        RECT 49.475 -166.765 49.805 -166.435 ;
        RECT 49.475 -168.125 49.805 -167.795 ;
        RECT 49.475 -169.485 49.805 -169.155 ;
        RECT 49.475 -170.845 49.805 -170.515 ;
        RECT 49.475 -172.205 49.805 -171.875 ;
        RECT 49.475 -173.565 49.805 -173.235 ;
        RECT 49.475 -174.925 49.805 -174.595 ;
        RECT 49.475 -176.285 49.805 -175.955 ;
        RECT 49.475 -177.645 49.805 -177.315 ;
        RECT 49.475 -183.29 49.805 -182.16 ;
        RECT 49.48 -183.405 49.8 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.835 244.04 51.165 245.17 ;
        RECT 50.835 239.875 51.165 240.205 ;
        RECT 50.835 238.515 51.165 238.845 ;
        RECT 50.835 237.155 51.165 237.485 ;
        RECT 50.84 237.155 51.16 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.835 -96.045 51.165 -95.715 ;
        RECT 50.835 -97.405 51.165 -97.075 ;
        RECT 50.835 -98.765 51.165 -98.435 ;
        RECT 50.835 -100.125 51.165 -99.795 ;
        RECT 50.835 -101.485 51.165 -101.155 ;
        RECT 50.835 -102.845 51.165 -102.515 ;
        RECT 50.835 -104.205 51.165 -103.875 ;
        RECT 50.835 -105.565 51.165 -105.235 ;
        RECT 50.835 -106.925 51.165 -106.595 ;
        RECT 50.835 -108.285 51.165 -107.955 ;
        RECT 50.835 -109.645 51.165 -109.315 ;
        RECT 50.835 -111.005 51.165 -110.675 ;
        RECT 50.835 -112.365 51.165 -112.035 ;
        RECT 50.835 -113.725 51.165 -113.395 ;
        RECT 50.835 -115.085 51.165 -114.755 ;
        RECT 50.835 -116.445 51.165 -116.115 ;
        RECT 50.835 -117.805 51.165 -117.475 ;
        RECT 50.835 -119.165 51.165 -118.835 ;
        RECT 50.835 -120.525 51.165 -120.195 ;
        RECT 50.835 -121.885 51.165 -121.555 ;
        RECT 50.835 -123.245 51.165 -122.915 ;
        RECT 50.835 -124.605 51.165 -124.275 ;
        RECT 50.835 -125.965 51.165 -125.635 ;
        RECT 50.835 -127.325 51.165 -126.995 ;
        RECT 50.835 -128.685 51.165 -128.355 ;
        RECT 50.835 -130.045 51.165 -129.715 ;
        RECT 50.835 -131.405 51.165 -131.075 ;
        RECT 50.835 -132.765 51.165 -132.435 ;
        RECT 50.835 -134.125 51.165 -133.795 ;
        RECT 50.835 -135.485 51.165 -135.155 ;
        RECT 50.835 -136.845 51.165 -136.515 ;
        RECT 50.835 -138.205 51.165 -137.875 ;
        RECT 50.835 -139.565 51.165 -139.235 ;
        RECT 50.835 -140.925 51.165 -140.595 ;
        RECT 50.835 -142.285 51.165 -141.955 ;
        RECT 50.835 -143.645 51.165 -143.315 ;
        RECT 50.835 -145.005 51.165 -144.675 ;
        RECT 50.835 -146.365 51.165 -146.035 ;
        RECT 50.835 -147.725 51.165 -147.395 ;
        RECT 50.835 -149.085 51.165 -148.755 ;
        RECT 50.835 -150.445 51.165 -150.115 ;
        RECT 50.835 -151.805 51.165 -151.475 ;
        RECT 50.835 -153.165 51.165 -152.835 ;
        RECT 50.835 -154.525 51.165 -154.195 ;
        RECT 50.835 -155.885 51.165 -155.555 ;
        RECT 50.835 -157.245 51.165 -156.915 ;
        RECT 50.835 -158.605 51.165 -158.275 ;
        RECT 50.835 -159.965 51.165 -159.635 ;
        RECT 50.835 -161.325 51.165 -160.995 ;
        RECT 50.835 -162.685 51.165 -162.355 ;
        RECT 50.835 -164.045 51.165 -163.715 ;
        RECT 50.835 -165.405 51.165 -165.075 ;
        RECT 50.835 -166.765 51.165 -166.435 ;
        RECT 50.835 -168.125 51.165 -167.795 ;
        RECT 50.835 -169.485 51.165 -169.155 ;
        RECT 50.835 -170.845 51.165 -170.515 ;
        RECT 50.835 -172.205 51.165 -171.875 ;
        RECT 50.835 -173.565 51.165 -173.235 ;
        RECT 50.835 -174.925 51.165 -174.595 ;
        RECT 50.835 -176.285 51.165 -175.955 ;
        RECT 50.835 -177.645 51.165 -177.315 ;
        RECT 50.835 -183.29 51.165 -182.16 ;
        RECT 50.84 -183.405 51.16 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.46 -94.075 51.79 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.195 244.04 52.525 245.17 ;
        RECT 52.195 239.875 52.525 240.205 ;
        RECT 52.195 238.515 52.525 238.845 ;
        RECT 52.195 237.155 52.525 237.485 ;
        RECT 52.2 237.155 52.52 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.555 244.04 53.885 245.17 ;
        RECT 53.555 239.875 53.885 240.205 ;
        RECT 53.555 238.515 53.885 238.845 ;
        RECT 53.555 237.155 53.885 237.485 ;
        RECT 53.56 237.155 53.88 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.555 -0.845 53.885 -0.515 ;
        RECT 53.555 -2.205 53.885 -1.875 ;
        RECT 53.555 -3.565 53.885 -3.235 ;
        RECT 53.56 -3.565 53.88 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.555 -91.965 53.885 -91.635 ;
        RECT 53.555 -93.325 53.885 -92.995 ;
        RECT 53.555 -94.685 53.885 -94.355 ;
        RECT 53.555 -96.045 53.885 -95.715 ;
        RECT 53.555 -97.405 53.885 -97.075 ;
        RECT 53.555 -98.765 53.885 -98.435 ;
        RECT 53.555 -100.125 53.885 -99.795 ;
        RECT 53.555 -101.485 53.885 -101.155 ;
        RECT 53.555 -102.845 53.885 -102.515 ;
        RECT 53.555 -104.205 53.885 -103.875 ;
        RECT 53.555 -105.565 53.885 -105.235 ;
        RECT 53.555 -106.925 53.885 -106.595 ;
        RECT 53.555 -108.285 53.885 -107.955 ;
        RECT 53.555 -109.645 53.885 -109.315 ;
        RECT 53.555 -111.005 53.885 -110.675 ;
        RECT 53.555 -112.365 53.885 -112.035 ;
        RECT 53.555 -113.725 53.885 -113.395 ;
        RECT 53.555 -115.085 53.885 -114.755 ;
        RECT 53.555 -116.445 53.885 -116.115 ;
        RECT 53.555 -117.805 53.885 -117.475 ;
        RECT 53.555 -119.165 53.885 -118.835 ;
        RECT 53.555 -120.525 53.885 -120.195 ;
        RECT 53.555 -121.885 53.885 -121.555 ;
        RECT 53.555 -123.245 53.885 -122.915 ;
        RECT 53.555 -124.605 53.885 -124.275 ;
        RECT 53.555 -125.965 53.885 -125.635 ;
        RECT 53.555 -127.325 53.885 -126.995 ;
        RECT 53.555 -128.685 53.885 -128.355 ;
        RECT 53.555 -130.045 53.885 -129.715 ;
        RECT 53.555 -131.405 53.885 -131.075 ;
        RECT 53.555 -132.765 53.885 -132.435 ;
        RECT 53.555 -134.125 53.885 -133.795 ;
        RECT 53.555 -135.485 53.885 -135.155 ;
        RECT 53.555 -136.845 53.885 -136.515 ;
        RECT 53.555 -138.205 53.885 -137.875 ;
        RECT 53.555 -139.565 53.885 -139.235 ;
        RECT 53.555 -140.925 53.885 -140.595 ;
        RECT 53.555 -142.285 53.885 -141.955 ;
        RECT 53.555 -143.645 53.885 -143.315 ;
        RECT 53.555 -145.005 53.885 -144.675 ;
        RECT 53.555 -146.365 53.885 -146.035 ;
        RECT 53.555 -147.725 53.885 -147.395 ;
        RECT 53.555 -149.085 53.885 -148.755 ;
        RECT 53.555 -150.445 53.885 -150.115 ;
        RECT 53.555 -151.805 53.885 -151.475 ;
        RECT 53.555 -153.165 53.885 -152.835 ;
        RECT 53.555 -154.525 53.885 -154.195 ;
        RECT 53.555 -155.885 53.885 -155.555 ;
        RECT 53.555 -157.245 53.885 -156.915 ;
        RECT 53.555 -158.605 53.885 -158.275 ;
        RECT 53.555 -159.965 53.885 -159.635 ;
        RECT 53.555 -161.325 53.885 -160.995 ;
        RECT 53.555 -162.685 53.885 -162.355 ;
        RECT 53.555 -164.045 53.885 -163.715 ;
        RECT 53.555 -165.405 53.885 -165.075 ;
        RECT 53.555 -166.765 53.885 -166.435 ;
        RECT 53.555 -168.125 53.885 -167.795 ;
        RECT 53.555 -169.485 53.885 -169.155 ;
        RECT 53.555 -170.845 53.885 -170.515 ;
        RECT 53.555 -172.205 53.885 -171.875 ;
        RECT 53.555 -173.565 53.885 -173.235 ;
        RECT 53.555 -174.925 53.885 -174.595 ;
        RECT 53.555 -176.285 53.885 -175.955 ;
        RECT 53.555 -177.645 53.885 -177.315 ;
        RECT 53.555 -183.29 53.885 -182.16 ;
        RECT 53.56 -183.405 53.88 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.915 244.04 55.245 245.17 ;
        RECT 54.915 239.875 55.245 240.205 ;
        RECT 54.915 238.515 55.245 238.845 ;
        RECT 54.915 237.155 55.245 237.485 ;
        RECT 54.92 237.155 55.24 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.915 -0.845 55.245 -0.515 ;
        RECT 54.915 -2.205 55.245 -1.875 ;
        RECT 54.915 -3.565 55.245 -3.235 ;
        RECT 54.92 -3.565 55.24 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.275 244.04 56.605 245.17 ;
        RECT 56.275 239.875 56.605 240.205 ;
        RECT 56.275 238.515 56.605 238.845 ;
        RECT 56.275 237.155 56.605 237.485 ;
        RECT 56.28 237.155 56.6 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.275 -0.845 56.605 -0.515 ;
        RECT 56.275 -2.205 56.605 -1.875 ;
        RECT 56.275 -3.565 56.605 -3.235 ;
        RECT 56.28 -3.565 56.6 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.275 -91.965 56.605 -91.635 ;
        RECT 56.275 -93.325 56.605 -92.995 ;
        RECT 56.275 -94.685 56.605 -94.355 ;
        RECT 56.275 -96.045 56.605 -95.715 ;
        RECT 56.275 -97.405 56.605 -97.075 ;
        RECT 56.275 -98.765 56.605 -98.435 ;
        RECT 56.275 -100.125 56.605 -99.795 ;
        RECT 56.275 -101.485 56.605 -101.155 ;
        RECT 56.275 -102.845 56.605 -102.515 ;
        RECT 56.275 -104.205 56.605 -103.875 ;
        RECT 56.275 -105.565 56.605 -105.235 ;
        RECT 56.275 -106.925 56.605 -106.595 ;
        RECT 56.275 -108.285 56.605 -107.955 ;
        RECT 56.275 -109.645 56.605 -109.315 ;
        RECT 56.275 -111.005 56.605 -110.675 ;
        RECT 56.275 -112.365 56.605 -112.035 ;
        RECT 56.275 -113.725 56.605 -113.395 ;
        RECT 56.275 -115.085 56.605 -114.755 ;
        RECT 56.275 -116.445 56.605 -116.115 ;
        RECT 56.275 -117.805 56.605 -117.475 ;
        RECT 56.275 -119.165 56.605 -118.835 ;
        RECT 56.275 -120.525 56.605 -120.195 ;
        RECT 56.275 -121.885 56.605 -121.555 ;
        RECT 56.275 -123.245 56.605 -122.915 ;
        RECT 56.275 -124.605 56.605 -124.275 ;
        RECT 56.275 -125.965 56.605 -125.635 ;
        RECT 56.275 -127.325 56.605 -126.995 ;
        RECT 56.275 -128.685 56.605 -128.355 ;
        RECT 56.275 -130.045 56.605 -129.715 ;
        RECT 56.275 -131.405 56.605 -131.075 ;
        RECT 56.275 -132.765 56.605 -132.435 ;
        RECT 56.275 -134.125 56.605 -133.795 ;
        RECT 56.275 -135.485 56.605 -135.155 ;
        RECT 56.275 -136.845 56.605 -136.515 ;
        RECT 56.275 -138.205 56.605 -137.875 ;
        RECT 56.275 -139.565 56.605 -139.235 ;
        RECT 56.275 -140.925 56.605 -140.595 ;
        RECT 56.275 -142.285 56.605 -141.955 ;
        RECT 56.275 -143.645 56.605 -143.315 ;
        RECT 56.275 -145.005 56.605 -144.675 ;
        RECT 56.275 -146.365 56.605 -146.035 ;
        RECT 56.275 -147.725 56.605 -147.395 ;
        RECT 56.275 -149.085 56.605 -148.755 ;
        RECT 56.275 -150.445 56.605 -150.115 ;
        RECT 56.275 -151.805 56.605 -151.475 ;
        RECT 56.275 -153.165 56.605 -152.835 ;
        RECT 56.275 -154.525 56.605 -154.195 ;
        RECT 56.275 -155.885 56.605 -155.555 ;
        RECT 56.275 -157.245 56.605 -156.915 ;
        RECT 56.275 -158.605 56.605 -158.275 ;
        RECT 56.275 -159.965 56.605 -159.635 ;
        RECT 56.275 -161.325 56.605 -160.995 ;
        RECT 56.275 -162.685 56.605 -162.355 ;
        RECT 56.275 -164.045 56.605 -163.715 ;
        RECT 56.275 -165.405 56.605 -165.075 ;
        RECT 56.275 -166.765 56.605 -166.435 ;
        RECT 56.275 -168.125 56.605 -167.795 ;
        RECT 56.275 -169.485 56.605 -169.155 ;
        RECT 56.275 -170.845 56.605 -170.515 ;
        RECT 56.275 -172.205 56.605 -171.875 ;
        RECT 56.275 -173.565 56.605 -173.235 ;
        RECT 56.275 -174.925 56.605 -174.595 ;
        RECT 56.275 -176.285 56.605 -175.955 ;
        RECT 56.275 -177.645 56.605 -177.315 ;
        RECT 56.275 -183.29 56.605 -182.16 ;
        RECT 56.28 -183.405 56.6 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.56 -94.075 57.89 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.635 244.04 57.965 245.17 ;
        RECT 57.635 239.875 57.965 240.205 ;
        RECT 57.635 238.515 57.965 238.845 ;
        RECT 57.635 237.155 57.965 237.485 ;
        RECT 57.64 237.155 57.96 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.635 -96.045 57.965 -95.715 ;
        RECT 57.635 -97.405 57.965 -97.075 ;
        RECT 57.635 -98.765 57.965 -98.435 ;
        RECT 57.635 -100.125 57.965 -99.795 ;
        RECT 57.635 -101.485 57.965 -101.155 ;
        RECT 57.635 -102.845 57.965 -102.515 ;
        RECT 57.635 -104.205 57.965 -103.875 ;
        RECT 57.635 -105.565 57.965 -105.235 ;
        RECT 57.635 -106.925 57.965 -106.595 ;
        RECT 57.635 -108.285 57.965 -107.955 ;
        RECT 57.635 -109.645 57.965 -109.315 ;
        RECT 57.635 -111.005 57.965 -110.675 ;
        RECT 57.635 -112.365 57.965 -112.035 ;
        RECT 57.635 -113.725 57.965 -113.395 ;
        RECT 57.635 -115.085 57.965 -114.755 ;
        RECT 57.635 -116.445 57.965 -116.115 ;
        RECT 57.635 -117.805 57.965 -117.475 ;
        RECT 57.635 -119.165 57.965 -118.835 ;
        RECT 57.635 -120.525 57.965 -120.195 ;
        RECT 57.635 -121.885 57.965 -121.555 ;
        RECT 57.635 -123.245 57.965 -122.915 ;
        RECT 57.635 -124.605 57.965 -124.275 ;
        RECT 57.635 -125.965 57.965 -125.635 ;
        RECT 57.635 -127.325 57.965 -126.995 ;
        RECT 57.635 -128.685 57.965 -128.355 ;
        RECT 57.635 -130.045 57.965 -129.715 ;
        RECT 57.635 -131.405 57.965 -131.075 ;
        RECT 57.635 -132.765 57.965 -132.435 ;
        RECT 57.635 -134.125 57.965 -133.795 ;
        RECT 57.635 -135.485 57.965 -135.155 ;
        RECT 57.635 -136.845 57.965 -136.515 ;
        RECT 57.635 -138.205 57.965 -137.875 ;
        RECT 57.635 -139.565 57.965 -139.235 ;
        RECT 57.635 -140.925 57.965 -140.595 ;
        RECT 57.635 -142.285 57.965 -141.955 ;
        RECT 57.635 -143.645 57.965 -143.315 ;
        RECT 57.635 -145.005 57.965 -144.675 ;
        RECT 57.635 -146.365 57.965 -146.035 ;
        RECT 57.635 -147.725 57.965 -147.395 ;
        RECT 57.635 -149.085 57.965 -148.755 ;
        RECT 57.635 -150.445 57.965 -150.115 ;
        RECT 57.635 -151.805 57.965 -151.475 ;
        RECT 57.635 -153.165 57.965 -152.835 ;
        RECT 57.635 -154.525 57.965 -154.195 ;
        RECT 57.635 -155.885 57.965 -155.555 ;
        RECT 57.635 -157.245 57.965 -156.915 ;
        RECT 57.635 -158.605 57.965 -158.275 ;
        RECT 57.635 -159.965 57.965 -159.635 ;
        RECT 57.635 -161.325 57.965 -160.995 ;
        RECT 57.635 -162.685 57.965 -162.355 ;
        RECT 57.635 -164.045 57.965 -163.715 ;
        RECT 57.635 -165.405 57.965 -165.075 ;
        RECT 57.635 -166.765 57.965 -166.435 ;
        RECT 57.635 -168.125 57.965 -167.795 ;
        RECT 57.635 -169.485 57.965 -169.155 ;
        RECT 57.635 -170.845 57.965 -170.515 ;
        RECT 57.635 -172.205 57.965 -171.875 ;
        RECT 57.635 -173.565 57.965 -173.235 ;
        RECT 57.635 -174.925 57.965 -174.595 ;
        RECT 57.635 -176.285 57.965 -175.955 ;
        RECT 57.635 -177.645 57.965 -177.315 ;
        RECT 57.635 -183.29 57.965 -182.16 ;
        RECT 57.64 -183.405 57.96 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.995 244.04 59.325 245.17 ;
        RECT 58.995 239.875 59.325 240.205 ;
        RECT 58.995 238.515 59.325 238.845 ;
        RECT 58.995 237.155 59.325 237.485 ;
        RECT 59 237.155 59.32 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.995 -0.845 59.325 -0.515 ;
        RECT 58.995 -2.205 59.325 -1.875 ;
        RECT 58.995 -3.565 59.325 -3.235 ;
        RECT 59 -3.565 59.32 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.355 244.04 60.685 245.17 ;
        RECT 60.355 239.875 60.685 240.205 ;
        RECT 60.355 238.515 60.685 238.845 ;
        RECT 60.355 237.155 60.685 237.485 ;
        RECT 60.36 237.155 60.68 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.355 -0.845 60.685 -0.515 ;
        RECT 60.355 -2.205 60.685 -1.875 ;
        RECT 60.355 -3.565 60.685 -3.235 ;
        RECT 60.36 -3.565 60.68 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.715 244.04 62.045 245.17 ;
        RECT 61.715 239.875 62.045 240.205 ;
        RECT 61.715 238.515 62.045 238.845 ;
        RECT 61.715 237.155 62.045 237.485 ;
        RECT 61.72 237.155 62.04 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.715 -0.845 62.045 -0.515 ;
        RECT 61.715 -2.205 62.045 -1.875 ;
        RECT 61.715 -3.565 62.045 -3.235 ;
        RECT 61.72 -3.565 62.04 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.715 -91.965 62.045 -91.635 ;
        RECT 61.715 -93.325 62.045 -92.995 ;
        RECT 61.715 -94.685 62.045 -94.355 ;
        RECT 61.715 -96.045 62.045 -95.715 ;
        RECT 61.715 -97.405 62.045 -97.075 ;
        RECT 61.715 -98.765 62.045 -98.435 ;
        RECT 61.715 -100.125 62.045 -99.795 ;
        RECT 61.715 -101.485 62.045 -101.155 ;
        RECT 61.715 -102.845 62.045 -102.515 ;
        RECT 61.715 -104.205 62.045 -103.875 ;
        RECT 61.715 -105.565 62.045 -105.235 ;
        RECT 61.715 -106.925 62.045 -106.595 ;
        RECT 61.715 -108.285 62.045 -107.955 ;
        RECT 61.715 -109.645 62.045 -109.315 ;
        RECT 61.715 -111.005 62.045 -110.675 ;
        RECT 61.715 -112.365 62.045 -112.035 ;
        RECT 61.715 -113.725 62.045 -113.395 ;
        RECT 61.715 -115.085 62.045 -114.755 ;
        RECT 61.715 -116.445 62.045 -116.115 ;
        RECT 61.715 -117.805 62.045 -117.475 ;
        RECT 61.715 -119.165 62.045 -118.835 ;
        RECT 61.715 -120.525 62.045 -120.195 ;
        RECT 61.715 -121.885 62.045 -121.555 ;
        RECT 61.715 -123.245 62.045 -122.915 ;
        RECT 61.715 -124.605 62.045 -124.275 ;
        RECT 61.715 -125.965 62.045 -125.635 ;
        RECT 61.715 -127.325 62.045 -126.995 ;
        RECT 61.715 -128.685 62.045 -128.355 ;
        RECT 61.715 -130.045 62.045 -129.715 ;
        RECT 61.715 -131.405 62.045 -131.075 ;
        RECT 61.715 -132.765 62.045 -132.435 ;
        RECT 61.715 -134.125 62.045 -133.795 ;
        RECT 61.715 -135.485 62.045 -135.155 ;
        RECT 61.715 -136.845 62.045 -136.515 ;
        RECT 61.715 -138.205 62.045 -137.875 ;
        RECT 61.715 -139.565 62.045 -139.235 ;
        RECT 61.715 -140.925 62.045 -140.595 ;
        RECT 61.715 -142.285 62.045 -141.955 ;
        RECT 61.715 -143.645 62.045 -143.315 ;
        RECT 61.715 -145.005 62.045 -144.675 ;
        RECT 61.715 -146.365 62.045 -146.035 ;
        RECT 61.715 -147.725 62.045 -147.395 ;
        RECT 61.715 -149.085 62.045 -148.755 ;
        RECT 61.715 -150.445 62.045 -150.115 ;
        RECT 61.715 -151.805 62.045 -151.475 ;
        RECT 61.715 -153.165 62.045 -152.835 ;
        RECT 61.715 -154.525 62.045 -154.195 ;
        RECT 61.715 -155.885 62.045 -155.555 ;
        RECT 61.715 -157.245 62.045 -156.915 ;
        RECT 61.715 -158.605 62.045 -158.275 ;
        RECT 61.715 -159.965 62.045 -159.635 ;
        RECT 61.715 -161.325 62.045 -160.995 ;
        RECT 61.715 -162.685 62.045 -162.355 ;
        RECT 61.715 -164.045 62.045 -163.715 ;
        RECT 61.715 -165.405 62.045 -165.075 ;
        RECT 61.715 -166.765 62.045 -166.435 ;
        RECT 61.715 -168.125 62.045 -167.795 ;
        RECT 61.715 -169.485 62.045 -169.155 ;
        RECT 61.715 -170.845 62.045 -170.515 ;
        RECT 61.715 -172.205 62.045 -171.875 ;
        RECT 61.715 -173.565 62.045 -173.235 ;
        RECT 61.715 -174.925 62.045 -174.595 ;
        RECT 61.715 -176.285 62.045 -175.955 ;
        RECT 61.715 -177.645 62.045 -177.315 ;
        RECT 61.715 -183.29 62.045 -182.16 ;
        RECT 61.72 -183.405 62.04 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.075 244.04 63.405 245.17 ;
        RECT 63.075 239.875 63.405 240.205 ;
        RECT 63.075 238.515 63.405 238.845 ;
        RECT 63.075 237.155 63.405 237.485 ;
        RECT 63.08 237.155 63.4 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.075 -96.045 63.405 -95.715 ;
        RECT 63.075 -97.405 63.405 -97.075 ;
        RECT 63.075 -98.765 63.405 -98.435 ;
        RECT 63.075 -100.125 63.405 -99.795 ;
        RECT 63.075 -101.485 63.405 -101.155 ;
        RECT 63.075 -102.845 63.405 -102.515 ;
        RECT 63.075 -104.205 63.405 -103.875 ;
        RECT 63.075 -105.565 63.405 -105.235 ;
        RECT 63.075 -106.925 63.405 -106.595 ;
        RECT 63.075 -108.285 63.405 -107.955 ;
        RECT 63.075 -109.645 63.405 -109.315 ;
        RECT 63.075 -111.005 63.405 -110.675 ;
        RECT 63.075 -112.365 63.405 -112.035 ;
        RECT 63.075 -113.725 63.405 -113.395 ;
        RECT 63.075 -115.085 63.405 -114.755 ;
        RECT 63.075 -116.445 63.405 -116.115 ;
        RECT 63.075 -117.805 63.405 -117.475 ;
        RECT 63.075 -119.165 63.405 -118.835 ;
        RECT 63.075 -120.525 63.405 -120.195 ;
        RECT 63.075 -121.885 63.405 -121.555 ;
        RECT 63.075 -123.245 63.405 -122.915 ;
        RECT 63.075 -124.605 63.405 -124.275 ;
        RECT 63.075 -125.965 63.405 -125.635 ;
        RECT 63.075 -127.325 63.405 -126.995 ;
        RECT 63.075 -128.685 63.405 -128.355 ;
        RECT 63.075 -130.045 63.405 -129.715 ;
        RECT 63.075 -131.405 63.405 -131.075 ;
        RECT 63.075 -132.765 63.405 -132.435 ;
        RECT 63.075 -134.125 63.405 -133.795 ;
        RECT 63.075 -135.485 63.405 -135.155 ;
        RECT 63.075 -136.845 63.405 -136.515 ;
        RECT 63.075 -138.205 63.405 -137.875 ;
        RECT 63.075 -139.565 63.405 -139.235 ;
        RECT 63.075 -140.925 63.405 -140.595 ;
        RECT 63.075 -142.285 63.405 -141.955 ;
        RECT 63.075 -143.645 63.405 -143.315 ;
        RECT 63.075 -145.005 63.405 -144.675 ;
        RECT 63.075 -146.365 63.405 -146.035 ;
        RECT 63.075 -147.725 63.405 -147.395 ;
        RECT 63.075 -149.085 63.405 -148.755 ;
        RECT 63.075 -150.445 63.405 -150.115 ;
        RECT 63.075 -151.805 63.405 -151.475 ;
        RECT 63.075 -153.165 63.405 -152.835 ;
        RECT 63.075 -154.525 63.405 -154.195 ;
        RECT 63.075 -155.885 63.405 -155.555 ;
        RECT 63.075 -157.245 63.405 -156.915 ;
        RECT 63.075 -158.605 63.405 -158.275 ;
        RECT 63.075 -159.965 63.405 -159.635 ;
        RECT 63.075 -161.325 63.405 -160.995 ;
        RECT 63.075 -162.685 63.405 -162.355 ;
        RECT 63.075 -164.045 63.405 -163.715 ;
        RECT 63.075 -165.405 63.405 -165.075 ;
        RECT 63.075 -166.765 63.405 -166.435 ;
        RECT 63.075 -168.125 63.405 -167.795 ;
        RECT 63.075 -169.485 63.405 -169.155 ;
        RECT 63.075 -170.845 63.405 -170.515 ;
        RECT 63.075 -172.205 63.405 -171.875 ;
        RECT 63.075 -173.565 63.405 -173.235 ;
        RECT 63.075 -174.925 63.405 -174.595 ;
        RECT 63.075 -176.285 63.405 -175.955 ;
        RECT 63.075 -177.645 63.405 -177.315 ;
        RECT 63.075 -183.29 63.405 -182.16 ;
        RECT 63.08 -183.405 63.4 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.66 -94.075 63.99 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.435 244.04 64.765 245.17 ;
        RECT 64.435 239.875 64.765 240.205 ;
        RECT 64.435 238.515 64.765 238.845 ;
        RECT 64.435 237.155 64.765 237.485 ;
        RECT 64.44 237.155 64.76 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.795 244.04 66.125 245.17 ;
        RECT 65.795 239.875 66.125 240.205 ;
        RECT 65.795 238.515 66.125 238.845 ;
        RECT 65.795 237.155 66.125 237.485 ;
        RECT 65.8 237.155 66.12 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.795 -0.845 66.125 -0.515 ;
        RECT 65.795 -2.205 66.125 -1.875 ;
        RECT 65.795 -3.565 66.125 -3.235 ;
        RECT 65.8 -3.565 66.12 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.795 -91.965 66.125 -91.635 ;
        RECT 65.795 -93.325 66.125 -92.995 ;
        RECT 65.795 -94.685 66.125 -94.355 ;
        RECT 65.795 -96.045 66.125 -95.715 ;
        RECT 65.795 -97.405 66.125 -97.075 ;
        RECT 65.795 -98.765 66.125 -98.435 ;
        RECT 65.795 -100.125 66.125 -99.795 ;
        RECT 65.795 -101.485 66.125 -101.155 ;
        RECT 65.795 -102.845 66.125 -102.515 ;
        RECT 65.795 -104.205 66.125 -103.875 ;
        RECT 65.795 -105.565 66.125 -105.235 ;
        RECT 65.795 -106.925 66.125 -106.595 ;
        RECT 65.795 -108.285 66.125 -107.955 ;
        RECT 65.795 -109.645 66.125 -109.315 ;
        RECT 65.795 -111.005 66.125 -110.675 ;
        RECT 65.795 -112.365 66.125 -112.035 ;
        RECT 65.795 -113.725 66.125 -113.395 ;
        RECT 65.795 -115.085 66.125 -114.755 ;
        RECT 65.795 -116.445 66.125 -116.115 ;
        RECT 65.795 -117.805 66.125 -117.475 ;
        RECT 65.795 -119.165 66.125 -118.835 ;
        RECT 65.795 -120.525 66.125 -120.195 ;
        RECT 65.795 -121.885 66.125 -121.555 ;
        RECT 65.795 -123.245 66.125 -122.915 ;
        RECT 65.795 -124.605 66.125 -124.275 ;
        RECT 65.795 -125.965 66.125 -125.635 ;
        RECT 65.795 -127.325 66.125 -126.995 ;
        RECT 65.795 -128.685 66.125 -128.355 ;
        RECT 65.795 -130.045 66.125 -129.715 ;
        RECT 65.795 -131.405 66.125 -131.075 ;
        RECT 65.795 -132.765 66.125 -132.435 ;
        RECT 65.795 -134.125 66.125 -133.795 ;
        RECT 65.795 -135.485 66.125 -135.155 ;
        RECT 65.795 -136.845 66.125 -136.515 ;
        RECT 65.795 -138.205 66.125 -137.875 ;
        RECT 65.795 -139.565 66.125 -139.235 ;
        RECT 65.795 -140.925 66.125 -140.595 ;
        RECT 65.795 -142.285 66.125 -141.955 ;
        RECT 65.795 -143.645 66.125 -143.315 ;
        RECT 65.795 -145.005 66.125 -144.675 ;
        RECT 65.795 -146.365 66.125 -146.035 ;
        RECT 65.795 -147.725 66.125 -147.395 ;
        RECT 65.795 -149.085 66.125 -148.755 ;
        RECT 65.795 -150.445 66.125 -150.115 ;
        RECT 65.795 -151.805 66.125 -151.475 ;
        RECT 65.795 -153.165 66.125 -152.835 ;
        RECT 65.795 -154.525 66.125 -154.195 ;
        RECT 65.795 -155.885 66.125 -155.555 ;
        RECT 65.795 -157.245 66.125 -156.915 ;
        RECT 65.795 -158.605 66.125 -158.275 ;
        RECT 65.795 -159.965 66.125 -159.635 ;
        RECT 65.795 -161.325 66.125 -160.995 ;
        RECT 65.795 -162.685 66.125 -162.355 ;
        RECT 65.795 -164.045 66.125 -163.715 ;
        RECT 65.795 -165.405 66.125 -165.075 ;
        RECT 65.795 -166.765 66.125 -166.435 ;
        RECT 65.795 -168.125 66.125 -167.795 ;
        RECT 65.795 -169.485 66.125 -169.155 ;
        RECT 65.795 -170.845 66.125 -170.515 ;
        RECT 65.795 -172.205 66.125 -171.875 ;
        RECT 65.795 -173.565 66.125 -173.235 ;
        RECT 65.795 -174.925 66.125 -174.595 ;
        RECT 65.795 -176.285 66.125 -175.955 ;
        RECT 65.795 -177.645 66.125 -177.315 ;
        RECT 65.795 -183.29 66.125 -182.16 ;
        RECT 65.8 -183.405 66.12 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.155 244.04 67.485 245.17 ;
        RECT 67.155 239.875 67.485 240.205 ;
        RECT 67.155 238.515 67.485 238.845 ;
        RECT 67.155 237.155 67.485 237.485 ;
        RECT 67.16 237.155 67.48 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.155 -0.845 67.485 -0.515 ;
        RECT 67.155 -2.205 67.485 -1.875 ;
        RECT 67.155 -3.565 67.485 -3.235 ;
        RECT 67.16 -3.565 67.48 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.515 244.04 68.845 245.17 ;
        RECT 68.515 239.875 68.845 240.205 ;
        RECT 68.515 238.515 68.845 238.845 ;
        RECT 68.515 237.155 68.845 237.485 ;
        RECT 68.52 237.155 68.84 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.515 -0.845 68.845 -0.515 ;
        RECT 68.515 -2.205 68.845 -1.875 ;
        RECT 68.515 -3.565 68.845 -3.235 ;
        RECT 68.52 -3.565 68.84 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.515 -91.965 68.845 -91.635 ;
        RECT 68.515 -93.325 68.845 -92.995 ;
        RECT 68.515 -94.685 68.845 -94.355 ;
        RECT 68.515 -96.045 68.845 -95.715 ;
        RECT 68.515 -97.405 68.845 -97.075 ;
        RECT 68.515 -98.765 68.845 -98.435 ;
        RECT 68.515 -100.125 68.845 -99.795 ;
        RECT 68.515 -101.485 68.845 -101.155 ;
        RECT 68.515 -102.845 68.845 -102.515 ;
        RECT 68.515 -104.205 68.845 -103.875 ;
        RECT 68.515 -105.565 68.845 -105.235 ;
        RECT 68.515 -106.925 68.845 -106.595 ;
        RECT 68.515 -108.285 68.845 -107.955 ;
        RECT 68.515 -109.645 68.845 -109.315 ;
        RECT 68.515 -111.005 68.845 -110.675 ;
        RECT 68.515 -112.365 68.845 -112.035 ;
        RECT 68.515 -113.725 68.845 -113.395 ;
        RECT 68.515 -115.085 68.845 -114.755 ;
        RECT 68.515 -116.445 68.845 -116.115 ;
        RECT 68.515 -117.805 68.845 -117.475 ;
        RECT 68.515 -119.165 68.845 -118.835 ;
        RECT 68.515 -120.525 68.845 -120.195 ;
        RECT 68.515 -121.885 68.845 -121.555 ;
        RECT 68.515 -123.245 68.845 -122.915 ;
        RECT 68.515 -124.605 68.845 -124.275 ;
        RECT 68.515 -125.965 68.845 -125.635 ;
        RECT 68.515 -127.325 68.845 -126.995 ;
        RECT 68.515 -128.685 68.845 -128.355 ;
        RECT 68.515 -130.045 68.845 -129.715 ;
        RECT 68.515 -131.405 68.845 -131.075 ;
        RECT 68.515 -132.765 68.845 -132.435 ;
        RECT 68.515 -134.125 68.845 -133.795 ;
        RECT 68.515 -135.485 68.845 -135.155 ;
        RECT 68.515 -136.845 68.845 -136.515 ;
        RECT 68.515 -138.205 68.845 -137.875 ;
        RECT 68.515 -139.565 68.845 -139.235 ;
        RECT 68.515 -140.925 68.845 -140.595 ;
        RECT 68.515 -142.285 68.845 -141.955 ;
        RECT 68.515 -143.645 68.845 -143.315 ;
        RECT 68.515 -145.005 68.845 -144.675 ;
        RECT 68.515 -146.365 68.845 -146.035 ;
        RECT 68.515 -147.725 68.845 -147.395 ;
        RECT 68.515 -149.085 68.845 -148.755 ;
        RECT 68.515 -150.445 68.845 -150.115 ;
        RECT 68.515 -151.805 68.845 -151.475 ;
        RECT 68.515 -153.165 68.845 -152.835 ;
        RECT 68.515 -154.525 68.845 -154.195 ;
        RECT 68.515 -155.885 68.845 -155.555 ;
        RECT 68.515 -157.245 68.845 -156.915 ;
        RECT 68.515 -158.605 68.845 -158.275 ;
        RECT 68.515 -159.965 68.845 -159.635 ;
        RECT 68.515 -161.325 68.845 -160.995 ;
        RECT 68.515 -162.685 68.845 -162.355 ;
        RECT 68.515 -164.045 68.845 -163.715 ;
        RECT 68.515 -165.405 68.845 -165.075 ;
        RECT 68.515 -166.765 68.845 -166.435 ;
        RECT 68.515 -168.125 68.845 -167.795 ;
        RECT 68.515 -169.485 68.845 -169.155 ;
        RECT 68.515 -170.845 68.845 -170.515 ;
        RECT 68.515 -172.205 68.845 -171.875 ;
        RECT 68.515 -173.565 68.845 -173.235 ;
        RECT 68.515 -174.925 68.845 -174.595 ;
        RECT 68.515 -176.285 68.845 -175.955 ;
        RECT 68.515 -177.645 68.845 -177.315 ;
        RECT 68.515 -183.29 68.845 -182.16 ;
        RECT 68.52 -183.405 68.84 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.76 -94.075 70.09 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.875 244.04 70.205 245.17 ;
        RECT 69.875 239.875 70.205 240.205 ;
        RECT 69.875 238.515 70.205 238.845 ;
        RECT 69.875 237.155 70.205 237.485 ;
        RECT 69.88 237.155 70.2 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.875 -96.045 70.205 -95.715 ;
        RECT 69.875 -97.405 70.205 -97.075 ;
        RECT 69.875 -98.765 70.205 -98.435 ;
        RECT 69.875 -100.125 70.205 -99.795 ;
        RECT 69.875 -101.485 70.205 -101.155 ;
        RECT 69.875 -102.845 70.205 -102.515 ;
        RECT 69.875 -104.205 70.205 -103.875 ;
        RECT 69.875 -105.565 70.205 -105.235 ;
        RECT 69.875 -106.925 70.205 -106.595 ;
        RECT 69.875 -108.285 70.205 -107.955 ;
        RECT 69.875 -109.645 70.205 -109.315 ;
        RECT 69.875 -111.005 70.205 -110.675 ;
        RECT 69.875 -112.365 70.205 -112.035 ;
        RECT 69.875 -113.725 70.205 -113.395 ;
        RECT 69.875 -115.085 70.205 -114.755 ;
        RECT 69.875 -116.445 70.205 -116.115 ;
        RECT 69.875 -117.805 70.205 -117.475 ;
        RECT 69.875 -119.165 70.205 -118.835 ;
        RECT 69.875 -120.525 70.205 -120.195 ;
        RECT 69.875 -121.885 70.205 -121.555 ;
        RECT 69.875 -123.245 70.205 -122.915 ;
        RECT 69.875 -124.605 70.205 -124.275 ;
        RECT 69.875 -125.965 70.205 -125.635 ;
        RECT 69.875 -127.325 70.205 -126.995 ;
        RECT 69.875 -128.685 70.205 -128.355 ;
        RECT 69.875 -130.045 70.205 -129.715 ;
        RECT 69.875 -131.405 70.205 -131.075 ;
        RECT 69.875 -132.765 70.205 -132.435 ;
        RECT 69.875 -134.125 70.205 -133.795 ;
        RECT 69.875 -135.485 70.205 -135.155 ;
        RECT 69.875 -136.845 70.205 -136.515 ;
        RECT 69.875 -138.205 70.205 -137.875 ;
        RECT 69.875 -139.565 70.205 -139.235 ;
        RECT 69.875 -140.925 70.205 -140.595 ;
        RECT 69.875 -142.285 70.205 -141.955 ;
        RECT 69.875 -143.645 70.205 -143.315 ;
        RECT 69.875 -145.005 70.205 -144.675 ;
        RECT 69.875 -146.365 70.205 -146.035 ;
        RECT 69.875 -147.725 70.205 -147.395 ;
        RECT 69.875 -149.085 70.205 -148.755 ;
        RECT 69.875 -150.445 70.205 -150.115 ;
        RECT 69.875 -151.805 70.205 -151.475 ;
        RECT 69.875 -153.165 70.205 -152.835 ;
        RECT 69.875 -154.525 70.205 -154.195 ;
        RECT 69.875 -155.885 70.205 -155.555 ;
        RECT 69.875 -157.245 70.205 -156.915 ;
        RECT 69.875 -158.605 70.205 -158.275 ;
        RECT 69.875 -159.965 70.205 -159.635 ;
        RECT 69.875 -161.325 70.205 -160.995 ;
        RECT 69.875 -162.685 70.205 -162.355 ;
        RECT 69.875 -164.045 70.205 -163.715 ;
        RECT 69.875 -165.405 70.205 -165.075 ;
        RECT 69.875 -166.765 70.205 -166.435 ;
        RECT 69.875 -168.125 70.205 -167.795 ;
        RECT 69.875 -169.485 70.205 -169.155 ;
        RECT 69.875 -170.845 70.205 -170.515 ;
        RECT 69.875 -172.205 70.205 -171.875 ;
        RECT 69.875 -173.565 70.205 -173.235 ;
        RECT 69.875 -174.925 70.205 -174.595 ;
        RECT 69.875 -176.285 70.205 -175.955 ;
        RECT 69.875 -177.645 70.205 -177.315 ;
        RECT 69.875 -183.29 70.205 -182.16 ;
        RECT 69.88 -183.405 70.2 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.235 244.04 71.565 245.17 ;
        RECT 71.235 239.875 71.565 240.205 ;
        RECT 71.235 238.515 71.565 238.845 ;
        RECT 71.235 237.155 71.565 237.485 ;
        RECT 71.24 237.155 71.56 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.235 -0.845 71.565 -0.515 ;
        RECT 71.235 -2.205 71.565 -1.875 ;
        RECT 71.235 -3.565 71.565 -3.235 ;
        RECT 71.24 -3.565 71.56 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.595 244.04 72.925 245.17 ;
        RECT 72.595 239.875 72.925 240.205 ;
        RECT 72.595 238.515 72.925 238.845 ;
        RECT 72.595 237.155 72.925 237.485 ;
        RECT 72.6 237.155 72.92 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.595 -0.845 72.925 -0.515 ;
        RECT 72.595 -2.205 72.925 -1.875 ;
        RECT 72.595 -3.565 72.925 -3.235 ;
        RECT 72.6 -3.565 72.92 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.955 244.04 74.285 245.17 ;
        RECT 73.955 239.875 74.285 240.205 ;
        RECT 73.955 238.515 74.285 238.845 ;
        RECT 73.955 237.155 74.285 237.485 ;
        RECT 73.96 237.155 74.28 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.955 -0.845 74.285 -0.515 ;
        RECT 73.955 -2.205 74.285 -1.875 ;
        RECT 73.955 -3.565 74.285 -3.235 ;
        RECT 73.96 -3.565 74.28 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.955 -119.165 74.285 -118.835 ;
        RECT 73.955 -120.525 74.285 -120.195 ;
        RECT 73.955 -121.885 74.285 -121.555 ;
        RECT 73.955 -123.245 74.285 -122.915 ;
        RECT 73.955 -124.605 74.285 -124.275 ;
        RECT 73.955 -125.965 74.285 -125.635 ;
        RECT 73.955 -127.325 74.285 -126.995 ;
        RECT 73.955 -128.685 74.285 -128.355 ;
        RECT 73.955 -130.045 74.285 -129.715 ;
        RECT 73.955 -131.405 74.285 -131.075 ;
        RECT 73.955 -132.765 74.285 -132.435 ;
        RECT 73.955 -134.125 74.285 -133.795 ;
        RECT 73.955 -135.485 74.285 -135.155 ;
        RECT 73.955 -136.845 74.285 -136.515 ;
        RECT 73.955 -138.205 74.285 -137.875 ;
        RECT 73.955 -139.565 74.285 -139.235 ;
        RECT 73.955 -140.925 74.285 -140.595 ;
        RECT 73.955 -142.285 74.285 -141.955 ;
        RECT 73.955 -143.645 74.285 -143.315 ;
        RECT 73.955 -145.005 74.285 -144.675 ;
        RECT 73.955 -146.365 74.285 -146.035 ;
        RECT 73.955 -147.725 74.285 -147.395 ;
        RECT 73.955 -149.085 74.285 -148.755 ;
        RECT 73.955 -150.445 74.285 -150.115 ;
        RECT 73.955 -151.805 74.285 -151.475 ;
        RECT 73.955 -153.165 74.285 -152.835 ;
        RECT 73.955 -154.525 74.285 -154.195 ;
        RECT 73.955 -155.885 74.285 -155.555 ;
        RECT 73.955 -157.245 74.285 -156.915 ;
        RECT 73.955 -158.605 74.285 -158.275 ;
        RECT 73.955 -159.965 74.285 -159.635 ;
        RECT 73.955 -161.325 74.285 -160.995 ;
        RECT 73.955 -162.685 74.285 -162.355 ;
        RECT 73.955 -164.045 74.285 -163.715 ;
        RECT 73.955 -165.405 74.285 -165.075 ;
        RECT 73.955 -166.765 74.285 -166.435 ;
        RECT 73.955 -168.125 74.285 -167.795 ;
        RECT 73.955 -169.485 74.285 -169.155 ;
        RECT 73.955 -170.845 74.285 -170.515 ;
        RECT 73.955 -172.205 74.285 -171.875 ;
        RECT 73.955 -173.565 74.285 -173.235 ;
        RECT 73.955 -174.925 74.285 -174.595 ;
        RECT 73.955 -176.285 74.285 -175.955 ;
        RECT 73.955 -177.645 74.285 -177.315 ;
        RECT 73.955 -183.29 74.285 -182.16 ;
        RECT 73.96 -183.405 74.28 -90.96 ;
        RECT 73.955 -91.965 74.285 -91.635 ;
        RECT 73.955 -93.325 74.285 -92.995 ;
        RECT 73.955 -94.685 74.285 -94.355 ;
        RECT 73.955 -96.045 74.285 -95.715 ;
        RECT 73.955 -97.405 74.285 -97.075 ;
        RECT 73.955 -98.765 74.285 -98.435 ;
        RECT 73.955 -100.125 74.285 -99.795 ;
        RECT 73.955 -101.485 74.285 -101.155 ;
        RECT 73.955 -102.845 74.285 -102.515 ;
        RECT 73.955 -104.205 74.285 -103.875 ;
        RECT 73.955 -105.565 74.285 -105.235 ;
        RECT 73.955 -106.925 74.285 -106.595 ;
        RECT 73.955 -108.285 74.285 -107.955 ;
        RECT 73.955 -109.645 74.285 -109.315 ;
        RECT 73.955 -111.005 74.285 -110.675 ;
        RECT 73.955 -112.365 74.285 -112.035 ;
        RECT 73.955 -113.725 74.285 -113.395 ;
        RECT 73.955 -115.085 74.285 -114.755 ;
        RECT 73.955 -116.445 74.285 -116.115 ;
        RECT 73.955 -117.805 74.285 -117.475 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.76 -94.075 9.09 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.035 244.04 10.365 245.17 ;
        RECT 10.035 239.875 10.365 240.205 ;
        RECT 10.035 238.515 10.365 238.845 ;
        RECT 10.035 237.155 10.365 237.485 ;
        RECT 10.04 237.155 10.36 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.395 244.04 11.725 245.17 ;
        RECT 11.395 239.875 11.725 240.205 ;
        RECT 11.395 238.515 11.725 238.845 ;
        RECT 11.395 237.155 11.725 237.485 ;
        RECT 11.4 237.155 11.72 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.395 -0.845 11.725 -0.515 ;
        RECT 11.395 -2.205 11.725 -1.875 ;
        RECT 11.395 -3.565 11.725 -3.235 ;
        RECT 11.4 -3.565 11.72 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.755 244.04 13.085 245.17 ;
        RECT 12.755 239.875 13.085 240.205 ;
        RECT 12.755 238.515 13.085 238.845 ;
        RECT 12.755 237.155 13.085 237.485 ;
        RECT 12.76 237.155 13.08 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.755 -0.845 13.085 -0.515 ;
        RECT 12.755 -2.205 13.085 -1.875 ;
        RECT 12.755 -3.565 13.085 -3.235 ;
        RECT 12.76 -3.565 13.08 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.755 -91.965 13.085 -91.635 ;
        RECT 12.755 -93.325 13.085 -92.995 ;
        RECT 12.755 -94.685 13.085 -94.355 ;
        RECT 12.755 -96.045 13.085 -95.715 ;
        RECT 12.755 -97.405 13.085 -97.075 ;
        RECT 12.755 -98.765 13.085 -98.435 ;
        RECT 12.755 -100.125 13.085 -99.795 ;
        RECT 12.755 -101.485 13.085 -101.155 ;
        RECT 12.755 -102.845 13.085 -102.515 ;
        RECT 12.755 -104.205 13.085 -103.875 ;
        RECT 12.755 -105.565 13.085 -105.235 ;
        RECT 12.755 -106.925 13.085 -106.595 ;
        RECT 12.755 -108.285 13.085 -107.955 ;
        RECT 12.755 -109.645 13.085 -109.315 ;
        RECT 12.755 -111.005 13.085 -110.675 ;
        RECT 12.755 -112.365 13.085 -112.035 ;
        RECT 12.755 -113.725 13.085 -113.395 ;
        RECT 12.755 -115.085 13.085 -114.755 ;
        RECT 12.755 -116.445 13.085 -116.115 ;
        RECT 12.755 -117.805 13.085 -117.475 ;
        RECT 12.755 -119.165 13.085 -118.835 ;
        RECT 12.755 -120.525 13.085 -120.195 ;
        RECT 12.755 -121.885 13.085 -121.555 ;
        RECT 12.755 -123.245 13.085 -122.915 ;
        RECT 12.755 -124.605 13.085 -124.275 ;
        RECT 12.755 -125.965 13.085 -125.635 ;
        RECT 12.755 -127.325 13.085 -126.995 ;
        RECT 12.755 -128.685 13.085 -128.355 ;
        RECT 12.755 -130.045 13.085 -129.715 ;
        RECT 12.755 -131.405 13.085 -131.075 ;
        RECT 12.755 -132.765 13.085 -132.435 ;
        RECT 12.755 -134.125 13.085 -133.795 ;
        RECT 12.755 -135.485 13.085 -135.155 ;
        RECT 12.755 -136.845 13.085 -136.515 ;
        RECT 12.755 -138.205 13.085 -137.875 ;
        RECT 12.755 -139.565 13.085 -139.235 ;
        RECT 12.755 -140.925 13.085 -140.595 ;
        RECT 12.755 -142.285 13.085 -141.955 ;
        RECT 12.755 -143.645 13.085 -143.315 ;
        RECT 12.755 -145.005 13.085 -144.675 ;
        RECT 12.755 -146.365 13.085 -146.035 ;
        RECT 12.755 -147.725 13.085 -147.395 ;
        RECT 12.755 -149.085 13.085 -148.755 ;
        RECT 12.755 -150.445 13.085 -150.115 ;
        RECT 12.755 -151.805 13.085 -151.475 ;
        RECT 12.755 -153.165 13.085 -152.835 ;
        RECT 12.755 -154.525 13.085 -154.195 ;
        RECT 12.755 -155.885 13.085 -155.555 ;
        RECT 12.755 -157.245 13.085 -156.915 ;
        RECT 12.755 -158.605 13.085 -158.275 ;
        RECT 12.755 -159.965 13.085 -159.635 ;
        RECT 12.755 -161.325 13.085 -160.995 ;
        RECT 12.755 -162.685 13.085 -162.355 ;
        RECT 12.755 -164.045 13.085 -163.715 ;
        RECT 12.755 -165.405 13.085 -165.075 ;
        RECT 12.755 -166.765 13.085 -166.435 ;
        RECT 12.755 -168.125 13.085 -167.795 ;
        RECT 12.755 -169.485 13.085 -169.155 ;
        RECT 12.755 -170.845 13.085 -170.515 ;
        RECT 12.755 -172.205 13.085 -171.875 ;
        RECT 12.755 -173.565 13.085 -173.235 ;
        RECT 12.755 -174.925 13.085 -174.595 ;
        RECT 12.755 -176.285 13.085 -175.955 ;
        RECT 12.755 -177.645 13.085 -177.315 ;
        RECT 12.755 -183.29 13.085 -182.16 ;
        RECT 12.76 -183.405 13.08 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.115 244.04 14.445 245.17 ;
        RECT 14.115 239.875 14.445 240.205 ;
        RECT 14.115 238.515 14.445 238.845 ;
        RECT 14.115 237.155 14.445 237.485 ;
        RECT 14.12 237.155 14.44 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.115 -0.845 14.445 -0.515 ;
        RECT 14.115 -2.205 14.445 -1.875 ;
        RECT 14.115 -3.565 14.445 -3.235 ;
        RECT 14.12 -3.565 14.44 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.115 -91.965 14.445 -91.635 ;
        RECT 14.115 -93.325 14.445 -92.995 ;
        RECT 14.115 -94.685 14.445 -94.355 ;
        RECT 14.115 -96.045 14.445 -95.715 ;
        RECT 14.115 -97.405 14.445 -97.075 ;
        RECT 14.115 -98.765 14.445 -98.435 ;
        RECT 14.115 -100.125 14.445 -99.795 ;
        RECT 14.115 -101.485 14.445 -101.155 ;
        RECT 14.115 -102.845 14.445 -102.515 ;
        RECT 14.115 -104.205 14.445 -103.875 ;
        RECT 14.115 -105.565 14.445 -105.235 ;
        RECT 14.115 -106.925 14.445 -106.595 ;
        RECT 14.115 -108.285 14.445 -107.955 ;
        RECT 14.115 -109.645 14.445 -109.315 ;
        RECT 14.115 -111.005 14.445 -110.675 ;
        RECT 14.115 -112.365 14.445 -112.035 ;
        RECT 14.115 -113.725 14.445 -113.395 ;
        RECT 14.115 -115.085 14.445 -114.755 ;
        RECT 14.115 -116.445 14.445 -116.115 ;
        RECT 14.115 -117.805 14.445 -117.475 ;
        RECT 14.115 -119.165 14.445 -118.835 ;
        RECT 14.115 -120.525 14.445 -120.195 ;
        RECT 14.115 -121.885 14.445 -121.555 ;
        RECT 14.115 -123.245 14.445 -122.915 ;
        RECT 14.115 -124.605 14.445 -124.275 ;
        RECT 14.115 -125.965 14.445 -125.635 ;
        RECT 14.115 -127.325 14.445 -126.995 ;
        RECT 14.115 -128.685 14.445 -128.355 ;
        RECT 14.115 -130.045 14.445 -129.715 ;
        RECT 14.115 -131.405 14.445 -131.075 ;
        RECT 14.115 -132.765 14.445 -132.435 ;
        RECT 14.115 -134.125 14.445 -133.795 ;
        RECT 14.115 -135.485 14.445 -135.155 ;
        RECT 14.115 -136.845 14.445 -136.515 ;
        RECT 14.115 -138.205 14.445 -137.875 ;
        RECT 14.115 -139.565 14.445 -139.235 ;
        RECT 14.115 -140.925 14.445 -140.595 ;
        RECT 14.115 -142.285 14.445 -141.955 ;
        RECT 14.115 -143.645 14.445 -143.315 ;
        RECT 14.115 -145.005 14.445 -144.675 ;
        RECT 14.115 -146.365 14.445 -146.035 ;
        RECT 14.115 -147.725 14.445 -147.395 ;
        RECT 14.115 -149.085 14.445 -148.755 ;
        RECT 14.115 -150.445 14.445 -150.115 ;
        RECT 14.115 -151.805 14.445 -151.475 ;
        RECT 14.115 -153.165 14.445 -152.835 ;
        RECT 14.115 -154.525 14.445 -154.195 ;
        RECT 14.115 -155.885 14.445 -155.555 ;
        RECT 14.115 -157.245 14.445 -156.915 ;
        RECT 14.115 -158.605 14.445 -158.275 ;
        RECT 14.115 -159.965 14.445 -159.635 ;
        RECT 14.115 -161.325 14.445 -160.995 ;
        RECT 14.115 -162.685 14.445 -162.355 ;
        RECT 14.115 -164.045 14.445 -163.715 ;
        RECT 14.115 -165.405 14.445 -165.075 ;
        RECT 14.115 -166.765 14.445 -166.435 ;
        RECT 14.115 -168.125 14.445 -167.795 ;
        RECT 14.115 -169.485 14.445 -169.155 ;
        RECT 14.115 -170.845 14.445 -170.515 ;
        RECT 14.115 -172.205 14.445 -171.875 ;
        RECT 14.115 -173.565 14.445 -173.235 ;
        RECT 14.115 -174.925 14.445 -174.595 ;
        RECT 14.115 -176.285 14.445 -175.955 ;
        RECT 14.115 -177.645 14.445 -177.315 ;
        RECT 14.115 -183.29 14.445 -182.16 ;
        RECT 14.12 -183.405 14.44 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.86 -94.075 15.19 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.475 244.04 15.805 245.17 ;
        RECT 15.475 239.875 15.805 240.205 ;
        RECT 15.475 238.515 15.805 238.845 ;
        RECT 15.475 237.155 15.805 237.485 ;
        RECT 15.48 237.155 15.8 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.475 -96.045 15.805 -95.715 ;
        RECT 15.475 -97.405 15.805 -97.075 ;
        RECT 15.475 -98.765 15.805 -98.435 ;
        RECT 15.475 -100.125 15.805 -99.795 ;
        RECT 15.475 -101.485 15.805 -101.155 ;
        RECT 15.475 -102.845 15.805 -102.515 ;
        RECT 15.475 -104.205 15.805 -103.875 ;
        RECT 15.475 -105.565 15.805 -105.235 ;
        RECT 15.475 -106.925 15.805 -106.595 ;
        RECT 15.475 -108.285 15.805 -107.955 ;
        RECT 15.475 -109.645 15.805 -109.315 ;
        RECT 15.475 -111.005 15.805 -110.675 ;
        RECT 15.475 -112.365 15.805 -112.035 ;
        RECT 15.475 -113.725 15.805 -113.395 ;
        RECT 15.475 -115.085 15.805 -114.755 ;
        RECT 15.475 -116.445 15.805 -116.115 ;
        RECT 15.475 -117.805 15.805 -117.475 ;
        RECT 15.475 -119.165 15.805 -118.835 ;
        RECT 15.475 -120.525 15.805 -120.195 ;
        RECT 15.475 -121.885 15.805 -121.555 ;
        RECT 15.475 -123.245 15.805 -122.915 ;
        RECT 15.475 -124.605 15.805 -124.275 ;
        RECT 15.475 -125.965 15.805 -125.635 ;
        RECT 15.475 -127.325 15.805 -126.995 ;
        RECT 15.475 -128.685 15.805 -128.355 ;
        RECT 15.475 -130.045 15.805 -129.715 ;
        RECT 15.475 -131.405 15.805 -131.075 ;
        RECT 15.475 -132.765 15.805 -132.435 ;
        RECT 15.475 -134.125 15.805 -133.795 ;
        RECT 15.475 -135.485 15.805 -135.155 ;
        RECT 15.475 -136.845 15.805 -136.515 ;
        RECT 15.475 -138.205 15.805 -137.875 ;
        RECT 15.475 -139.565 15.805 -139.235 ;
        RECT 15.475 -140.925 15.805 -140.595 ;
        RECT 15.475 -142.285 15.805 -141.955 ;
        RECT 15.475 -143.645 15.805 -143.315 ;
        RECT 15.475 -145.005 15.805 -144.675 ;
        RECT 15.475 -146.365 15.805 -146.035 ;
        RECT 15.475 -147.725 15.805 -147.395 ;
        RECT 15.475 -149.085 15.805 -148.755 ;
        RECT 15.475 -150.445 15.805 -150.115 ;
        RECT 15.475 -151.805 15.805 -151.475 ;
        RECT 15.475 -153.165 15.805 -152.835 ;
        RECT 15.475 -154.525 15.805 -154.195 ;
        RECT 15.475 -155.885 15.805 -155.555 ;
        RECT 15.475 -157.245 15.805 -156.915 ;
        RECT 15.475 -158.605 15.805 -158.275 ;
        RECT 15.475 -159.965 15.805 -159.635 ;
        RECT 15.475 -161.325 15.805 -160.995 ;
        RECT 15.475 -162.685 15.805 -162.355 ;
        RECT 15.475 -164.045 15.805 -163.715 ;
        RECT 15.475 -165.405 15.805 -165.075 ;
        RECT 15.475 -166.765 15.805 -166.435 ;
        RECT 15.475 -168.125 15.805 -167.795 ;
        RECT 15.475 -169.485 15.805 -169.155 ;
        RECT 15.475 -170.845 15.805 -170.515 ;
        RECT 15.475 -172.205 15.805 -171.875 ;
        RECT 15.475 -173.565 15.805 -173.235 ;
        RECT 15.475 -174.925 15.805 -174.595 ;
        RECT 15.475 -176.285 15.805 -175.955 ;
        RECT 15.475 -177.645 15.805 -177.315 ;
        RECT 15.475 -183.29 15.805 -182.16 ;
        RECT 15.48 -183.405 15.8 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.835 244.04 17.165 245.17 ;
        RECT 16.835 239.875 17.165 240.205 ;
        RECT 16.835 238.515 17.165 238.845 ;
        RECT 16.835 237.155 17.165 237.485 ;
        RECT 16.84 237.155 17.16 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.835 -0.845 17.165 -0.515 ;
        RECT 16.835 -2.205 17.165 -1.875 ;
        RECT 16.835 -3.565 17.165 -3.235 ;
        RECT 16.84 -3.565 17.16 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.195 244.04 18.525 245.17 ;
        RECT 18.195 239.875 18.525 240.205 ;
        RECT 18.195 238.515 18.525 238.845 ;
        RECT 18.195 237.155 18.525 237.485 ;
        RECT 18.2 237.155 18.52 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.195 -0.845 18.525 -0.515 ;
        RECT 18.195 -2.205 18.525 -1.875 ;
        RECT 18.195 -3.565 18.525 -3.235 ;
        RECT 18.2 -3.565 18.52 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.555 244.04 19.885 245.17 ;
        RECT 19.555 239.875 19.885 240.205 ;
        RECT 19.555 238.515 19.885 238.845 ;
        RECT 19.555 237.155 19.885 237.485 ;
        RECT 19.56 237.155 19.88 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.555 -0.845 19.885 -0.515 ;
        RECT 19.555 -2.205 19.885 -1.875 ;
        RECT 19.555 -3.565 19.885 -3.235 ;
        RECT 19.56 -3.565 19.88 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.555 -91.965 19.885 -91.635 ;
        RECT 19.555 -93.325 19.885 -92.995 ;
        RECT 19.555 -94.685 19.885 -94.355 ;
        RECT 19.555 -96.045 19.885 -95.715 ;
        RECT 19.555 -97.405 19.885 -97.075 ;
        RECT 19.555 -98.765 19.885 -98.435 ;
        RECT 19.555 -100.125 19.885 -99.795 ;
        RECT 19.555 -101.485 19.885 -101.155 ;
        RECT 19.555 -102.845 19.885 -102.515 ;
        RECT 19.555 -104.205 19.885 -103.875 ;
        RECT 19.555 -105.565 19.885 -105.235 ;
        RECT 19.555 -106.925 19.885 -106.595 ;
        RECT 19.555 -108.285 19.885 -107.955 ;
        RECT 19.555 -109.645 19.885 -109.315 ;
        RECT 19.555 -111.005 19.885 -110.675 ;
        RECT 19.555 -112.365 19.885 -112.035 ;
        RECT 19.555 -113.725 19.885 -113.395 ;
        RECT 19.555 -115.085 19.885 -114.755 ;
        RECT 19.555 -116.445 19.885 -116.115 ;
        RECT 19.555 -117.805 19.885 -117.475 ;
        RECT 19.555 -119.165 19.885 -118.835 ;
        RECT 19.555 -120.525 19.885 -120.195 ;
        RECT 19.555 -121.885 19.885 -121.555 ;
        RECT 19.555 -123.245 19.885 -122.915 ;
        RECT 19.555 -124.605 19.885 -124.275 ;
        RECT 19.555 -125.965 19.885 -125.635 ;
        RECT 19.555 -127.325 19.885 -126.995 ;
        RECT 19.555 -128.685 19.885 -128.355 ;
        RECT 19.555 -130.045 19.885 -129.715 ;
        RECT 19.555 -131.405 19.885 -131.075 ;
        RECT 19.555 -132.765 19.885 -132.435 ;
        RECT 19.555 -134.125 19.885 -133.795 ;
        RECT 19.555 -135.485 19.885 -135.155 ;
        RECT 19.555 -136.845 19.885 -136.515 ;
        RECT 19.555 -138.205 19.885 -137.875 ;
        RECT 19.555 -139.565 19.885 -139.235 ;
        RECT 19.555 -140.925 19.885 -140.595 ;
        RECT 19.555 -142.285 19.885 -141.955 ;
        RECT 19.555 -143.645 19.885 -143.315 ;
        RECT 19.555 -145.005 19.885 -144.675 ;
        RECT 19.555 -146.365 19.885 -146.035 ;
        RECT 19.555 -147.725 19.885 -147.395 ;
        RECT 19.555 -149.085 19.885 -148.755 ;
        RECT 19.555 -150.445 19.885 -150.115 ;
        RECT 19.555 -151.805 19.885 -151.475 ;
        RECT 19.555 -153.165 19.885 -152.835 ;
        RECT 19.555 -154.525 19.885 -154.195 ;
        RECT 19.555 -155.885 19.885 -155.555 ;
        RECT 19.555 -157.245 19.885 -156.915 ;
        RECT 19.555 -158.605 19.885 -158.275 ;
        RECT 19.555 -159.965 19.885 -159.635 ;
        RECT 19.555 -161.325 19.885 -160.995 ;
        RECT 19.555 -162.685 19.885 -162.355 ;
        RECT 19.555 -164.045 19.885 -163.715 ;
        RECT 19.555 -165.405 19.885 -165.075 ;
        RECT 19.555 -166.765 19.885 -166.435 ;
        RECT 19.555 -168.125 19.885 -167.795 ;
        RECT 19.555 -169.485 19.885 -169.155 ;
        RECT 19.555 -170.845 19.885 -170.515 ;
        RECT 19.555 -172.205 19.885 -171.875 ;
        RECT 19.555 -173.565 19.885 -173.235 ;
        RECT 19.555 -174.925 19.885 -174.595 ;
        RECT 19.555 -176.285 19.885 -175.955 ;
        RECT 19.555 -177.645 19.885 -177.315 ;
        RECT 19.555 -183.29 19.885 -182.16 ;
        RECT 19.56 -183.405 19.88 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.915 244.04 21.245 245.17 ;
        RECT 20.915 239.875 21.245 240.205 ;
        RECT 20.915 238.515 21.245 238.845 ;
        RECT 20.915 237.155 21.245 237.485 ;
        RECT 20.92 237.155 21.24 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.915 -96.045 21.245 -95.715 ;
        RECT 20.915 -97.405 21.245 -97.075 ;
        RECT 20.915 -98.765 21.245 -98.435 ;
        RECT 20.915 -100.125 21.245 -99.795 ;
        RECT 20.915 -101.485 21.245 -101.155 ;
        RECT 20.915 -102.845 21.245 -102.515 ;
        RECT 20.915 -104.205 21.245 -103.875 ;
        RECT 20.915 -105.565 21.245 -105.235 ;
        RECT 20.915 -106.925 21.245 -106.595 ;
        RECT 20.915 -108.285 21.245 -107.955 ;
        RECT 20.915 -109.645 21.245 -109.315 ;
        RECT 20.915 -111.005 21.245 -110.675 ;
        RECT 20.915 -112.365 21.245 -112.035 ;
        RECT 20.915 -113.725 21.245 -113.395 ;
        RECT 20.915 -115.085 21.245 -114.755 ;
        RECT 20.915 -116.445 21.245 -116.115 ;
        RECT 20.915 -117.805 21.245 -117.475 ;
        RECT 20.915 -119.165 21.245 -118.835 ;
        RECT 20.915 -120.525 21.245 -120.195 ;
        RECT 20.915 -121.885 21.245 -121.555 ;
        RECT 20.915 -123.245 21.245 -122.915 ;
        RECT 20.915 -124.605 21.245 -124.275 ;
        RECT 20.915 -125.965 21.245 -125.635 ;
        RECT 20.915 -127.325 21.245 -126.995 ;
        RECT 20.915 -128.685 21.245 -128.355 ;
        RECT 20.915 -130.045 21.245 -129.715 ;
        RECT 20.915 -131.405 21.245 -131.075 ;
        RECT 20.915 -132.765 21.245 -132.435 ;
        RECT 20.915 -134.125 21.245 -133.795 ;
        RECT 20.915 -135.485 21.245 -135.155 ;
        RECT 20.915 -136.845 21.245 -136.515 ;
        RECT 20.915 -138.205 21.245 -137.875 ;
        RECT 20.915 -139.565 21.245 -139.235 ;
        RECT 20.915 -140.925 21.245 -140.595 ;
        RECT 20.915 -142.285 21.245 -141.955 ;
        RECT 20.915 -143.645 21.245 -143.315 ;
        RECT 20.915 -145.005 21.245 -144.675 ;
        RECT 20.915 -146.365 21.245 -146.035 ;
        RECT 20.915 -147.725 21.245 -147.395 ;
        RECT 20.915 -149.085 21.245 -148.755 ;
        RECT 20.915 -150.445 21.245 -150.115 ;
        RECT 20.915 -151.805 21.245 -151.475 ;
        RECT 20.915 -153.165 21.245 -152.835 ;
        RECT 20.915 -154.525 21.245 -154.195 ;
        RECT 20.915 -155.885 21.245 -155.555 ;
        RECT 20.915 -157.245 21.245 -156.915 ;
        RECT 20.915 -158.605 21.245 -158.275 ;
        RECT 20.915 -159.965 21.245 -159.635 ;
        RECT 20.915 -161.325 21.245 -160.995 ;
        RECT 20.915 -162.685 21.245 -162.355 ;
        RECT 20.915 -164.045 21.245 -163.715 ;
        RECT 20.915 -165.405 21.245 -165.075 ;
        RECT 20.915 -166.765 21.245 -166.435 ;
        RECT 20.915 -168.125 21.245 -167.795 ;
        RECT 20.915 -169.485 21.245 -169.155 ;
        RECT 20.915 -170.845 21.245 -170.515 ;
        RECT 20.915 -172.205 21.245 -171.875 ;
        RECT 20.915 -173.565 21.245 -173.235 ;
        RECT 20.915 -174.925 21.245 -174.595 ;
        RECT 20.915 -176.285 21.245 -175.955 ;
        RECT 20.915 -177.645 21.245 -177.315 ;
        RECT 20.915 -183.29 21.245 -182.16 ;
        RECT 20.92 -183.405 21.24 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.96 -94.075 21.29 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.275 244.04 22.605 245.17 ;
        RECT 22.275 239.875 22.605 240.205 ;
        RECT 22.275 238.515 22.605 238.845 ;
        RECT 22.275 237.155 22.605 237.485 ;
        RECT 22.28 237.155 22.6 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.635 244.04 23.965 245.17 ;
        RECT 23.635 239.875 23.965 240.205 ;
        RECT 23.635 238.515 23.965 238.845 ;
        RECT 23.635 237.155 23.965 237.485 ;
        RECT 23.64 237.155 23.96 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.635 -0.845 23.965 -0.515 ;
        RECT 23.635 -2.205 23.965 -1.875 ;
        RECT 23.635 -3.565 23.965 -3.235 ;
        RECT 23.64 -3.565 23.96 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.995 244.04 25.325 245.17 ;
        RECT 24.995 239.875 25.325 240.205 ;
        RECT 24.995 238.515 25.325 238.845 ;
        RECT 24.995 237.155 25.325 237.485 ;
        RECT 25 237.155 25.32 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.995 -0.845 25.325 -0.515 ;
        RECT 24.995 -2.205 25.325 -1.875 ;
        RECT 24.995 -3.565 25.325 -3.235 ;
        RECT 25 -3.565 25.32 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.995 -91.965 25.325 -91.635 ;
        RECT 24.995 -93.325 25.325 -92.995 ;
        RECT 24.995 -94.685 25.325 -94.355 ;
        RECT 24.995 -96.045 25.325 -95.715 ;
        RECT 24.995 -97.405 25.325 -97.075 ;
        RECT 24.995 -98.765 25.325 -98.435 ;
        RECT 24.995 -100.125 25.325 -99.795 ;
        RECT 24.995 -101.485 25.325 -101.155 ;
        RECT 24.995 -102.845 25.325 -102.515 ;
        RECT 24.995 -104.205 25.325 -103.875 ;
        RECT 24.995 -105.565 25.325 -105.235 ;
        RECT 24.995 -106.925 25.325 -106.595 ;
        RECT 24.995 -108.285 25.325 -107.955 ;
        RECT 24.995 -109.645 25.325 -109.315 ;
        RECT 24.995 -111.005 25.325 -110.675 ;
        RECT 24.995 -112.365 25.325 -112.035 ;
        RECT 24.995 -113.725 25.325 -113.395 ;
        RECT 24.995 -115.085 25.325 -114.755 ;
        RECT 24.995 -116.445 25.325 -116.115 ;
        RECT 24.995 -117.805 25.325 -117.475 ;
        RECT 24.995 -119.165 25.325 -118.835 ;
        RECT 24.995 -120.525 25.325 -120.195 ;
        RECT 24.995 -121.885 25.325 -121.555 ;
        RECT 24.995 -123.245 25.325 -122.915 ;
        RECT 24.995 -124.605 25.325 -124.275 ;
        RECT 24.995 -125.965 25.325 -125.635 ;
        RECT 24.995 -127.325 25.325 -126.995 ;
        RECT 24.995 -128.685 25.325 -128.355 ;
        RECT 24.995 -130.045 25.325 -129.715 ;
        RECT 24.995 -131.405 25.325 -131.075 ;
        RECT 24.995 -132.765 25.325 -132.435 ;
        RECT 24.995 -134.125 25.325 -133.795 ;
        RECT 24.995 -135.485 25.325 -135.155 ;
        RECT 24.995 -136.845 25.325 -136.515 ;
        RECT 24.995 -138.205 25.325 -137.875 ;
        RECT 24.995 -139.565 25.325 -139.235 ;
        RECT 24.995 -140.925 25.325 -140.595 ;
        RECT 24.995 -142.285 25.325 -141.955 ;
        RECT 24.995 -143.645 25.325 -143.315 ;
        RECT 24.995 -145.005 25.325 -144.675 ;
        RECT 24.995 -146.365 25.325 -146.035 ;
        RECT 24.995 -147.725 25.325 -147.395 ;
        RECT 24.995 -149.085 25.325 -148.755 ;
        RECT 24.995 -150.445 25.325 -150.115 ;
        RECT 24.995 -151.805 25.325 -151.475 ;
        RECT 24.995 -153.165 25.325 -152.835 ;
        RECT 24.995 -154.525 25.325 -154.195 ;
        RECT 24.995 -155.885 25.325 -155.555 ;
        RECT 24.995 -157.245 25.325 -156.915 ;
        RECT 24.995 -158.605 25.325 -158.275 ;
        RECT 24.995 -159.965 25.325 -159.635 ;
        RECT 24.995 -161.325 25.325 -160.995 ;
        RECT 24.995 -162.685 25.325 -162.355 ;
        RECT 24.995 -164.045 25.325 -163.715 ;
        RECT 24.995 -165.405 25.325 -165.075 ;
        RECT 24.995 -166.765 25.325 -166.435 ;
        RECT 24.995 -168.125 25.325 -167.795 ;
        RECT 24.995 -169.485 25.325 -169.155 ;
        RECT 24.995 -170.845 25.325 -170.515 ;
        RECT 24.995 -172.205 25.325 -171.875 ;
        RECT 24.995 -173.565 25.325 -173.235 ;
        RECT 24.995 -174.925 25.325 -174.595 ;
        RECT 24.995 -176.285 25.325 -175.955 ;
        RECT 24.995 -177.645 25.325 -177.315 ;
        RECT 24.995 -183.29 25.325 -182.16 ;
        RECT 25 -183.405 25.32 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.355 244.04 26.685 245.17 ;
        RECT 26.355 239.875 26.685 240.205 ;
        RECT 26.355 238.515 26.685 238.845 ;
        RECT 26.355 237.155 26.685 237.485 ;
        RECT 26.36 237.155 26.68 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.355 -0.845 26.685 -0.515 ;
        RECT 26.355 -2.205 26.685 -1.875 ;
        RECT 26.355 -3.565 26.685 -3.235 ;
        RECT 26.36 -3.565 26.68 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.355 -91.965 26.685 -91.635 ;
        RECT 26.355 -93.325 26.685 -92.995 ;
        RECT 26.355 -94.685 26.685 -94.355 ;
        RECT 26.355 -96.045 26.685 -95.715 ;
        RECT 26.355 -97.405 26.685 -97.075 ;
        RECT 26.355 -98.765 26.685 -98.435 ;
        RECT 26.355 -100.125 26.685 -99.795 ;
        RECT 26.355 -101.485 26.685 -101.155 ;
        RECT 26.355 -102.845 26.685 -102.515 ;
        RECT 26.355 -104.205 26.685 -103.875 ;
        RECT 26.355 -105.565 26.685 -105.235 ;
        RECT 26.355 -106.925 26.685 -106.595 ;
        RECT 26.355 -108.285 26.685 -107.955 ;
        RECT 26.355 -109.645 26.685 -109.315 ;
        RECT 26.355 -111.005 26.685 -110.675 ;
        RECT 26.355 -112.365 26.685 -112.035 ;
        RECT 26.355 -113.725 26.685 -113.395 ;
        RECT 26.355 -115.085 26.685 -114.755 ;
        RECT 26.355 -116.445 26.685 -116.115 ;
        RECT 26.355 -117.805 26.685 -117.475 ;
        RECT 26.355 -119.165 26.685 -118.835 ;
        RECT 26.355 -120.525 26.685 -120.195 ;
        RECT 26.355 -121.885 26.685 -121.555 ;
        RECT 26.355 -123.245 26.685 -122.915 ;
        RECT 26.355 -124.605 26.685 -124.275 ;
        RECT 26.355 -125.965 26.685 -125.635 ;
        RECT 26.355 -127.325 26.685 -126.995 ;
        RECT 26.355 -128.685 26.685 -128.355 ;
        RECT 26.355 -130.045 26.685 -129.715 ;
        RECT 26.355 -131.405 26.685 -131.075 ;
        RECT 26.355 -132.765 26.685 -132.435 ;
        RECT 26.355 -134.125 26.685 -133.795 ;
        RECT 26.355 -135.485 26.685 -135.155 ;
        RECT 26.355 -136.845 26.685 -136.515 ;
        RECT 26.355 -138.205 26.685 -137.875 ;
        RECT 26.355 -139.565 26.685 -139.235 ;
        RECT 26.355 -140.925 26.685 -140.595 ;
        RECT 26.355 -142.285 26.685 -141.955 ;
        RECT 26.355 -143.645 26.685 -143.315 ;
        RECT 26.355 -145.005 26.685 -144.675 ;
        RECT 26.355 -146.365 26.685 -146.035 ;
        RECT 26.355 -147.725 26.685 -147.395 ;
        RECT 26.355 -149.085 26.685 -148.755 ;
        RECT 26.355 -150.445 26.685 -150.115 ;
        RECT 26.355 -151.805 26.685 -151.475 ;
        RECT 26.355 -153.165 26.685 -152.835 ;
        RECT 26.355 -154.525 26.685 -154.195 ;
        RECT 26.355 -155.885 26.685 -155.555 ;
        RECT 26.355 -157.245 26.685 -156.915 ;
        RECT 26.355 -158.605 26.685 -158.275 ;
        RECT 26.355 -159.965 26.685 -159.635 ;
        RECT 26.355 -161.325 26.685 -160.995 ;
        RECT 26.355 -162.685 26.685 -162.355 ;
        RECT 26.355 -164.045 26.685 -163.715 ;
        RECT 26.355 -165.405 26.685 -165.075 ;
        RECT 26.355 -166.765 26.685 -166.435 ;
        RECT 26.355 -168.125 26.685 -167.795 ;
        RECT 26.355 -169.485 26.685 -169.155 ;
        RECT 26.355 -170.845 26.685 -170.515 ;
        RECT 26.355 -172.205 26.685 -171.875 ;
        RECT 26.355 -173.565 26.685 -173.235 ;
        RECT 26.355 -174.925 26.685 -174.595 ;
        RECT 26.355 -176.285 26.685 -175.955 ;
        RECT 26.355 -177.645 26.685 -177.315 ;
        RECT 26.355 -183.29 26.685 -182.16 ;
        RECT 26.36 -183.405 26.68 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.06 -94.075 27.39 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.715 244.04 28.045 245.17 ;
        RECT 27.715 239.875 28.045 240.205 ;
        RECT 27.715 238.515 28.045 238.845 ;
        RECT 27.715 237.155 28.045 237.485 ;
        RECT 27.72 237.155 28.04 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.715 -96.045 28.045 -95.715 ;
        RECT 27.715 -97.405 28.045 -97.075 ;
        RECT 27.715 -98.765 28.045 -98.435 ;
        RECT 27.715 -100.125 28.045 -99.795 ;
        RECT 27.715 -101.485 28.045 -101.155 ;
        RECT 27.715 -102.845 28.045 -102.515 ;
        RECT 27.715 -104.205 28.045 -103.875 ;
        RECT 27.715 -105.565 28.045 -105.235 ;
        RECT 27.715 -106.925 28.045 -106.595 ;
        RECT 27.715 -108.285 28.045 -107.955 ;
        RECT 27.715 -109.645 28.045 -109.315 ;
        RECT 27.715 -111.005 28.045 -110.675 ;
        RECT 27.715 -112.365 28.045 -112.035 ;
        RECT 27.715 -113.725 28.045 -113.395 ;
        RECT 27.715 -115.085 28.045 -114.755 ;
        RECT 27.715 -116.445 28.045 -116.115 ;
        RECT 27.715 -117.805 28.045 -117.475 ;
        RECT 27.715 -119.165 28.045 -118.835 ;
        RECT 27.715 -120.525 28.045 -120.195 ;
        RECT 27.715 -121.885 28.045 -121.555 ;
        RECT 27.715 -123.245 28.045 -122.915 ;
        RECT 27.715 -124.605 28.045 -124.275 ;
        RECT 27.715 -125.965 28.045 -125.635 ;
        RECT 27.715 -127.325 28.045 -126.995 ;
        RECT 27.715 -128.685 28.045 -128.355 ;
        RECT 27.715 -130.045 28.045 -129.715 ;
        RECT 27.715 -131.405 28.045 -131.075 ;
        RECT 27.715 -132.765 28.045 -132.435 ;
        RECT 27.715 -134.125 28.045 -133.795 ;
        RECT 27.715 -135.485 28.045 -135.155 ;
        RECT 27.715 -136.845 28.045 -136.515 ;
        RECT 27.715 -138.205 28.045 -137.875 ;
        RECT 27.715 -139.565 28.045 -139.235 ;
        RECT 27.715 -140.925 28.045 -140.595 ;
        RECT 27.715 -142.285 28.045 -141.955 ;
        RECT 27.715 -143.645 28.045 -143.315 ;
        RECT 27.715 -145.005 28.045 -144.675 ;
        RECT 27.715 -146.365 28.045 -146.035 ;
        RECT 27.715 -147.725 28.045 -147.395 ;
        RECT 27.715 -149.085 28.045 -148.755 ;
        RECT 27.715 -150.445 28.045 -150.115 ;
        RECT 27.715 -151.805 28.045 -151.475 ;
        RECT 27.715 -153.165 28.045 -152.835 ;
        RECT 27.715 -154.525 28.045 -154.195 ;
        RECT 27.715 -155.885 28.045 -155.555 ;
        RECT 27.715 -157.245 28.045 -156.915 ;
        RECT 27.715 -158.605 28.045 -158.275 ;
        RECT 27.715 -159.965 28.045 -159.635 ;
        RECT 27.715 -161.325 28.045 -160.995 ;
        RECT 27.715 -162.685 28.045 -162.355 ;
        RECT 27.715 -164.045 28.045 -163.715 ;
        RECT 27.715 -165.405 28.045 -165.075 ;
        RECT 27.715 -166.765 28.045 -166.435 ;
        RECT 27.715 -168.125 28.045 -167.795 ;
        RECT 27.715 -169.485 28.045 -169.155 ;
        RECT 27.715 -170.845 28.045 -170.515 ;
        RECT 27.715 -172.205 28.045 -171.875 ;
        RECT 27.715 -173.565 28.045 -173.235 ;
        RECT 27.715 -174.925 28.045 -174.595 ;
        RECT 27.715 -176.285 28.045 -175.955 ;
        RECT 27.715 -177.645 28.045 -177.315 ;
        RECT 27.715 -183.29 28.045 -182.16 ;
        RECT 27.72 -183.405 28.04 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.075 244.04 29.405 245.17 ;
        RECT 29.075 239.875 29.405 240.205 ;
        RECT 29.075 238.515 29.405 238.845 ;
        RECT 29.075 237.155 29.405 237.485 ;
        RECT 29.08 237.155 29.4 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.075 -0.845 29.405 -0.515 ;
        RECT 29.075 -2.205 29.405 -1.875 ;
        RECT 29.075 -3.565 29.405 -3.235 ;
        RECT 29.08 -3.565 29.4 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.435 244.04 30.765 245.17 ;
        RECT 30.435 239.875 30.765 240.205 ;
        RECT 30.435 238.515 30.765 238.845 ;
        RECT 30.435 237.155 30.765 237.485 ;
        RECT 30.44 237.155 30.76 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.435 -0.845 30.765 -0.515 ;
        RECT 30.435 -2.205 30.765 -1.875 ;
        RECT 30.435 -3.565 30.765 -3.235 ;
        RECT 30.44 -3.565 30.76 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.795 244.04 32.125 245.17 ;
        RECT 31.795 239.875 32.125 240.205 ;
        RECT 31.795 238.515 32.125 238.845 ;
        RECT 31.795 237.155 32.125 237.485 ;
        RECT 31.8 237.155 32.12 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.795 -0.845 32.125 -0.515 ;
        RECT 31.795 -2.205 32.125 -1.875 ;
        RECT 31.795 -3.565 32.125 -3.235 ;
        RECT 31.8 -3.565 32.12 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.795 -91.965 32.125 -91.635 ;
        RECT 31.795 -93.325 32.125 -92.995 ;
        RECT 31.795 -94.685 32.125 -94.355 ;
        RECT 31.795 -96.045 32.125 -95.715 ;
        RECT 31.795 -97.405 32.125 -97.075 ;
        RECT 31.795 -98.765 32.125 -98.435 ;
        RECT 31.795 -100.125 32.125 -99.795 ;
        RECT 31.795 -101.485 32.125 -101.155 ;
        RECT 31.795 -102.845 32.125 -102.515 ;
        RECT 31.795 -104.205 32.125 -103.875 ;
        RECT 31.795 -105.565 32.125 -105.235 ;
        RECT 31.795 -106.925 32.125 -106.595 ;
        RECT 31.795 -108.285 32.125 -107.955 ;
        RECT 31.795 -109.645 32.125 -109.315 ;
        RECT 31.795 -111.005 32.125 -110.675 ;
        RECT 31.795 -112.365 32.125 -112.035 ;
        RECT 31.795 -113.725 32.125 -113.395 ;
        RECT 31.795 -115.085 32.125 -114.755 ;
        RECT 31.795 -116.445 32.125 -116.115 ;
        RECT 31.795 -117.805 32.125 -117.475 ;
        RECT 31.795 -119.165 32.125 -118.835 ;
        RECT 31.795 -120.525 32.125 -120.195 ;
        RECT 31.795 -121.885 32.125 -121.555 ;
        RECT 31.795 -123.245 32.125 -122.915 ;
        RECT 31.795 -124.605 32.125 -124.275 ;
        RECT 31.795 -125.965 32.125 -125.635 ;
        RECT 31.795 -127.325 32.125 -126.995 ;
        RECT 31.795 -128.685 32.125 -128.355 ;
        RECT 31.795 -130.045 32.125 -129.715 ;
        RECT 31.795 -131.405 32.125 -131.075 ;
        RECT 31.795 -132.765 32.125 -132.435 ;
        RECT 31.795 -134.125 32.125 -133.795 ;
        RECT 31.795 -135.485 32.125 -135.155 ;
        RECT 31.795 -136.845 32.125 -136.515 ;
        RECT 31.795 -138.205 32.125 -137.875 ;
        RECT 31.795 -139.565 32.125 -139.235 ;
        RECT 31.795 -140.925 32.125 -140.595 ;
        RECT 31.795 -142.285 32.125 -141.955 ;
        RECT 31.795 -143.645 32.125 -143.315 ;
        RECT 31.795 -145.005 32.125 -144.675 ;
        RECT 31.795 -146.365 32.125 -146.035 ;
        RECT 31.795 -147.725 32.125 -147.395 ;
        RECT 31.795 -149.085 32.125 -148.755 ;
        RECT 31.795 -150.445 32.125 -150.115 ;
        RECT 31.795 -151.805 32.125 -151.475 ;
        RECT 31.795 -153.165 32.125 -152.835 ;
        RECT 31.795 -154.525 32.125 -154.195 ;
        RECT 31.795 -155.885 32.125 -155.555 ;
        RECT 31.795 -157.245 32.125 -156.915 ;
        RECT 31.795 -158.605 32.125 -158.275 ;
        RECT 31.795 -159.965 32.125 -159.635 ;
        RECT 31.795 -161.325 32.125 -160.995 ;
        RECT 31.795 -162.685 32.125 -162.355 ;
        RECT 31.795 -164.045 32.125 -163.715 ;
        RECT 31.795 -165.405 32.125 -165.075 ;
        RECT 31.795 -166.765 32.125 -166.435 ;
        RECT 31.795 -168.125 32.125 -167.795 ;
        RECT 31.795 -169.485 32.125 -169.155 ;
        RECT 31.795 -170.845 32.125 -170.515 ;
        RECT 31.795 -172.205 32.125 -171.875 ;
        RECT 31.795 -173.565 32.125 -173.235 ;
        RECT 31.795 -174.925 32.125 -174.595 ;
        RECT 31.795 -176.285 32.125 -175.955 ;
        RECT 31.795 -177.645 32.125 -177.315 ;
        RECT 31.795 -183.29 32.125 -182.16 ;
        RECT 31.8 -183.405 32.12 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.155 244.04 33.485 245.17 ;
        RECT 33.155 239.875 33.485 240.205 ;
        RECT 33.155 238.515 33.485 238.845 ;
        RECT 33.155 237.155 33.485 237.485 ;
        RECT 33.16 237.155 33.48 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.155 -96.045 33.485 -95.715 ;
        RECT 33.155 -97.405 33.485 -97.075 ;
        RECT 33.155 -98.765 33.485 -98.435 ;
        RECT 33.155 -100.125 33.485 -99.795 ;
        RECT 33.155 -101.485 33.485 -101.155 ;
        RECT 33.155 -102.845 33.485 -102.515 ;
        RECT 33.155 -104.205 33.485 -103.875 ;
        RECT 33.155 -105.565 33.485 -105.235 ;
        RECT 33.155 -106.925 33.485 -106.595 ;
        RECT 33.155 -108.285 33.485 -107.955 ;
        RECT 33.155 -109.645 33.485 -109.315 ;
        RECT 33.155 -111.005 33.485 -110.675 ;
        RECT 33.155 -112.365 33.485 -112.035 ;
        RECT 33.155 -113.725 33.485 -113.395 ;
        RECT 33.155 -115.085 33.485 -114.755 ;
        RECT 33.155 -116.445 33.485 -116.115 ;
        RECT 33.155 -117.805 33.485 -117.475 ;
        RECT 33.155 -119.165 33.485 -118.835 ;
        RECT 33.155 -120.525 33.485 -120.195 ;
        RECT 33.155 -121.885 33.485 -121.555 ;
        RECT 33.155 -123.245 33.485 -122.915 ;
        RECT 33.155 -124.605 33.485 -124.275 ;
        RECT 33.155 -125.965 33.485 -125.635 ;
        RECT 33.155 -127.325 33.485 -126.995 ;
        RECT 33.155 -128.685 33.485 -128.355 ;
        RECT 33.155 -130.045 33.485 -129.715 ;
        RECT 33.155 -131.405 33.485 -131.075 ;
        RECT 33.155 -132.765 33.485 -132.435 ;
        RECT 33.155 -134.125 33.485 -133.795 ;
        RECT 33.155 -135.485 33.485 -135.155 ;
        RECT 33.155 -136.845 33.485 -136.515 ;
        RECT 33.155 -138.205 33.485 -137.875 ;
        RECT 33.155 -139.565 33.485 -139.235 ;
        RECT 33.155 -140.925 33.485 -140.595 ;
        RECT 33.155 -142.285 33.485 -141.955 ;
        RECT 33.155 -143.645 33.485 -143.315 ;
        RECT 33.155 -145.005 33.485 -144.675 ;
        RECT 33.155 -146.365 33.485 -146.035 ;
        RECT 33.155 -147.725 33.485 -147.395 ;
        RECT 33.155 -149.085 33.485 -148.755 ;
        RECT 33.155 -150.445 33.485 -150.115 ;
        RECT 33.155 -151.805 33.485 -151.475 ;
        RECT 33.155 -153.165 33.485 -152.835 ;
        RECT 33.155 -154.525 33.485 -154.195 ;
        RECT 33.155 -155.885 33.485 -155.555 ;
        RECT 33.155 -157.245 33.485 -156.915 ;
        RECT 33.155 -158.605 33.485 -158.275 ;
        RECT 33.155 -159.965 33.485 -159.635 ;
        RECT 33.155 -161.325 33.485 -160.995 ;
        RECT 33.155 -162.685 33.485 -162.355 ;
        RECT 33.155 -164.045 33.485 -163.715 ;
        RECT 33.155 -165.405 33.485 -165.075 ;
        RECT 33.155 -166.765 33.485 -166.435 ;
        RECT 33.155 -168.125 33.485 -167.795 ;
        RECT 33.155 -169.485 33.485 -169.155 ;
        RECT 33.155 -170.845 33.485 -170.515 ;
        RECT 33.155 -172.205 33.485 -171.875 ;
        RECT 33.155 -173.565 33.485 -173.235 ;
        RECT 33.155 -174.925 33.485 -174.595 ;
        RECT 33.155 -176.285 33.485 -175.955 ;
        RECT 33.155 -177.645 33.485 -177.315 ;
        RECT 33.155 -183.29 33.485 -182.16 ;
        RECT 33.16 -183.405 33.48 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.16 -94.075 33.49 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.515 244.04 34.845 245.17 ;
        RECT 34.515 239.875 34.845 240.205 ;
        RECT 34.515 238.515 34.845 238.845 ;
        RECT 34.515 237.155 34.845 237.485 ;
        RECT 34.52 237.155 34.84 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.515 -0.845 34.845 -0.515 ;
        RECT 34.515 -2.205 34.845 -1.875 ;
        RECT 34.515 -3.565 34.845 -3.235 ;
        RECT 34.52 -3.565 34.84 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.875 244.04 36.205 245.17 ;
        RECT 35.875 239.875 36.205 240.205 ;
        RECT 35.875 238.515 36.205 238.845 ;
        RECT 35.875 237.155 36.205 237.485 ;
        RECT 35.88 237.155 36.2 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.875 -0.845 36.205 -0.515 ;
        RECT 35.875 -2.205 36.205 -1.875 ;
        RECT 35.875 -3.565 36.205 -3.235 ;
        RECT 35.88 -3.565 36.2 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.235 244.04 37.565 245.17 ;
        RECT 37.235 239.875 37.565 240.205 ;
        RECT 37.235 238.515 37.565 238.845 ;
        RECT 37.235 237.155 37.565 237.485 ;
        RECT 37.24 237.155 37.56 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.235 -0.845 37.565 -0.515 ;
        RECT 37.235 -2.205 37.565 -1.875 ;
        RECT 37.235 -3.565 37.565 -3.235 ;
        RECT 37.24 -3.565 37.56 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.235 -91.965 37.565 -91.635 ;
        RECT 37.235 -93.325 37.565 -92.995 ;
        RECT 37.235 -94.685 37.565 -94.355 ;
        RECT 37.235 -96.045 37.565 -95.715 ;
        RECT 37.235 -97.405 37.565 -97.075 ;
        RECT 37.235 -98.765 37.565 -98.435 ;
        RECT 37.235 -100.125 37.565 -99.795 ;
        RECT 37.235 -101.485 37.565 -101.155 ;
        RECT 37.235 -102.845 37.565 -102.515 ;
        RECT 37.235 -104.205 37.565 -103.875 ;
        RECT 37.235 -105.565 37.565 -105.235 ;
        RECT 37.235 -106.925 37.565 -106.595 ;
        RECT 37.235 -108.285 37.565 -107.955 ;
        RECT 37.235 -109.645 37.565 -109.315 ;
        RECT 37.235 -111.005 37.565 -110.675 ;
        RECT 37.235 -112.365 37.565 -112.035 ;
        RECT 37.235 -113.725 37.565 -113.395 ;
        RECT 37.235 -115.085 37.565 -114.755 ;
        RECT 37.235 -116.445 37.565 -116.115 ;
        RECT 37.235 -117.805 37.565 -117.475 ;
        RECT 37.235 -119.165 37.565 -118.835 ;
        RECT 37.235 -120.525 37.565 -120.195 ;
        RECT 37.235 -121.885 37.565 -121.555 ;
        RECT 37.235 -123.245 37.565 -122.915 ;
        RECT 37.235 -124.605 37.565 -124.275 ;
        RECT 37.235 -125.965 37.565 -125.635 ;
        RECT 37.235 -127.325 37.565 -126.995 ;
        RECT 37.235 -128.685 37.565 -128.355 ;
        RECT 37.235 -130.045 37.565 -129.715 ;
        RECT 37.235 -131.405 37.565 -131.075 ;
        RECT 37.235 -132.765 37.565 -132.435 ;
        RECT 37.235 -134.125 37.565 -133.795 ;
        RECT 37.235 -135.485 37.565 -135.155 ;
        RECT 37.235 -136.845 37.565 -136.515 ;
        RECT 37.235 -138.205 37.565 -137.875 ;
        RECT 37.235 -139.565 37.565 -139.235 ;
        RECT 37.235 -140.925 37.565 -140.595 ;
        RECT 37.235 -142.285 37.565 -141.955 ;
        RECT 37.235 -143.645 37.565 -143.315 ;
        RECT 37.235 -145.005 37.565 -144.675 ;
        RECT 37.235 -146.365 37.565 -146.035 ;
        RECT 37.235 -147.725 37.565 -147.395 ;
        RECT 37.235 -149.085 37.565 -148.755 ;
        RECT 37.235 -150.445 37.565 -150.115 ;
        RECT 37.235 -151.805 37.565 -151.475 ;
        RECT 37.235 -153.165 37.565 -152.835 ;
        RECT 37.235 -154.525 37.565 -154.195 ;
        RECT 37.235 -155.885 37.565 -155.555 ;
        RECT 37.235 -157.245 37.565 -156.915 ;
        RECT 37.235 -158.605 37.565 -158.275 ;
        RECT 37.235 -159.965 37.565 -159.635 ;
        RECT 37.235 -161.325 37.565 -160.995 ;
        RECT 37.235 -162.685 37.565 -162.355 ;
        RECT 37.235 -164.045 37.565 -163.715 ;
        RECT 37.235 -165.405 37.565 -165.075 ;
        RECT 37.235 -166.765 37.565 -166.435 ;
        RECT 37.235 -168.125 37.565 -167.795 ;
        RECT 37.235 -169.485 37.565 -169.155 ;
        RECT 37.235 -170.845 37.565 -170.515 ;
        RECT 37.235 -172.205 37.565 -171.875 ;
        RECT 37.235 -173.565 37.565 -173.235 ;
        RECT 37.235 -174.925 37.565 -174.595 ;
        RECT 37.235 -176.285 37.565 -175.955 ;
        RECT 37.235 -177.645 37.565 -177.315 ;
        RECT 37.235 -183.29 37.565 -182.16 ;
        RECT 37.24 -183.405 37.56 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.595 244.04 38.925 245.17 ;
        RECT 38.595 239.875 38.925 240.205 ;
        RECT 38.595 238.515 38.925 238.845 ;
        RECT 38.595 237.155 38.925 237.485 ;
        RECT 38.6 237.155 38.92 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.595 -96.045 38.925 -95.715 ;
        RECT 38.595 -97.405 38.925 -97.075 ;
        RECT 38.595 -98.765 38.925 -98.435 ;
        RECT 38.595 -100.125 38.925 -99.795 ;
        RECT 38.595 -101.485 38.925 -101.155 ;
        RECT 38.595 -102.845 38.925 -102.515 ;
        RECT 38.595 -104.205 38.925 -103.875 ;
        RECT 38.595 -105.565 38.925 -105.235 ;
        RECT 38.595 -106.925 38.925 -106.595 ;
        RECT 38.595 -108.285 38.925 -107.955 ;
        RECT 38.595 -109.645 38.925 -109.315 ;
        RECT 38.595 -111.005 38.925 -110.675 ;
        RECT 38.595 -112.365 38.925 -112.035 ;
        RECT 38.595 -113.725 38.925 -113.395 ;
        RECT 38.595 -115.085 38.925 -114.755 ;
        RECT 38.595 -116.445 38.925 -116.115 ;
        RECT 38.595 -117.805 38.925 -117.475 ;
        RECT 38.595 -119.165 38.925 -118.835 ;
        RECT 38.595 -120.525 38.925 -120.195 ;
        RECT 38.595 -121.885 38.925 -121.555 ;
        RECT 38.595 -123.245 38.925 -122.915 ;
        RECT 38.595 -124.605 38.925 -124.275 ;
        RECT 38.595 -125.965 38.925 -125.635 ;
        RECT 38.595 -127.325 38.925 -126.995 ;
        RECT 38.595 -128.685 38.925 -128.355 ;
        RECT 38.595 -130.045 38.925 -129.715 ;
        RECT 38.595 -131.405 38.925 -131.075 ;
        RECT 38.595 -132.765 38.925 -132.435 ;
        RECT 38.595 -134.125 38.925 -133.795 ;
        RECT 38.595 -135.485 38.925 -135.155 ;
        RECT 38.595 -136.845 38.925 -136.515 ;
        RECT 38.595 -138.205 38.925 -137.875 ;
        RECT 38.595 -139.565 38.925 -139.235 ;
        RECT 38.595 -140.925 38.925 -140.595 ;
        RECT 38.595 -142.285 38.925 -141.955 ;
        RECT 38.595 -143.645 38.925 -143.315 ;
        RECT 38.595 -145.005 38.925 -144.675 ;
        RECT 38.595 -146.365 38.925 -146.035 ;
        RECT 38.595 -147.725 38.925 -147.395 ;
        RECT 38.595 -149.085 38.925 -148.755 ;
        RECT 38.595 -150.445 38.925 -150.115 ;
        RECT 38.595 -151.805 38.925 -151.475 ;
        RECT 38.595 -153.165 38.925 -152.835 ;
        RECT 38.595 -154.525 38.925 -154.195 ;
        RECT 38.595 -155.885 38.925 -155.555 ;
        RECT 38.595 -157.245 38.925 -156.915 ;
        RECT 38.595 -158.605 38.925 -158.275 ;
        RECT 38.595 -159.965 38.925 -159.635 ;
        RECT 38.595 -161.325 38.925 -160.995 ;
        RECT 38.595 -162.685 38.925 -162.355 ;
        RECT 38.595 -164.045 38.925 -163.715 ;
        RECT 38.595 -165.405 38.925 -165.075 ;
        RECT 38.595 -166.765 38.925 -166.435 ;
        RECT 38.595 -168.125 38.925 -167.795 ;
        RECT 38.595 -169.485 38.925 -169.155 ;
        RECT 38.595 -170.845 38.925 -170.515 ;
        RECT 38.595 -172.205 38.925 -171.875 ;
        RECT 38.595 -173.565 38.925 -173.235 ;
        RECT 38.595 -174.925 38.925 -174.595 ;
        RECT 38.595 -176.285 38.925 -175.955 ;
        RECT 38.595 -177.645 38.925 -177.315 ;
        RECT 38.595 -183.29 38.925 -182.16 ;
        RECT 38.6 -183.405 38.92 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.26 -94.075 39.59 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.955 244.04 40.285 245.17 ;
        RECT 39.955 239.875 40.285 240.205 ;
        RECT 39.955 238.515 40.285 238.845 ;
        RECT 39.955 237.155 40.285 237.485 ;
        RECT 39.96 237.155 40.28 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.315 244.04 41.645 245.17 ;
        RECT 41.315 239.875 41.645 240.205 ;
        RECT 41.315 238.515 41.645 238.845 ;
        RECT 41.315 237.155 41.645 237.485 ;
        RECT 41.32 237.155 41.64 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.315 -0.845 41.645 -0.515 ;
        RECT 41.315 -2.205 41.645 -1.875 ;
        RECT 41.315 -3.565 41.645 -3.235 ;
        RECT 41.32 -3.565 41.64 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.675 244.04 43.005 245.17 ;
        RECT 42.675 239.875 43.005 240.205 ;
        RECT 42.675 238.515 43.005 238.845 ;
        RECT 42.675 237.155 43.005 237.485 ;
        RECT 42.68 237.155 43 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.675 -0.845 43.005 -0.515 ;
        RECT 42.675 -2.205 43.005 -1.875 ;
        RECT 42.675 -3.565 43.005 -3.235 ;
        RECT 42.68 -3.565 43 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.035 244.04 44.365 245.17 ;
        RECT 44.035 239.875 44.365 240.205 ;
        RECT 44.035 238.515 44.365 238.845 ;
        RECT 44.035 237.155 44.365 237.485 ;
        RECT 44.04 237.155 44.36 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.035 -3.565 44.365 -3.235 ;
        RECT 44.04 -3.565 44.36 -0.515 ;
        RECT 44.035 -0.845 44.365 -0.515 ;
        RECT 44.035 -2.205 44.365 -1.875 ;
    END
    PORT
      LAYER met3 ;
        RECT -2.205 244.04 -1.875 245.17 ;
        RECT -2.205 239.875 -1.875 240.205 ;
        RECT -2.205 238.515 -1.875 238.845 ;
        RECT -2.205 237.155 -1.875 237.485 ;
        RECT -2.205 235.17 -1.875 235.5 ;
        RECT -2.205 232.995 -1.875 233.325 ;
        RECT -2.205 231.415 -1.875 231.745 ;
        RECT -2.205 230.565 -1.875 230.895 ;
        RECT -2.205 228.255 -1.875 228.585 ;
        RECT -2.205 227.405 -1.875 227.735 ;
        RECT -2.205 225.095 -1.875 225.425 ;
        RECT -2.205 224.245 -1.875 224.575 ;
        RECT -2.205 221.935 -1.875 222.265 ;
        RECT -2.205 221.085 -1.875 221.415 ;
        RECT -2.205 218.775 -1.875 219.105 ;
        RECT -2.205 217.195 -1.875 217.525 ;
        RECT -2.205 216.345 -1.875 216.675 ;
        RECT -2.205 214.035 -1.875 214.365 ;
        RECT -2.205 213.185 -1.875 213.515 ;
        RECT -2.205 210.875 -1.875 211.205 ;
        RECT -2.205 210.025 -1.875 210.355 ;
        RECT -2.205 207.715 -1.875 208.045 ;
        RECT -2.205 206.865 -1.875 207.195 ;
        RECT -2.205 204.555 -1.875 204.885 ;
        RECT -2.205 202.975 -1.875 203.305 ;
        RECT -2.205 202.125 -1.875 202.455 ;
        RECT -2.205 199.815 -1.875 200.145 ;
        RECT -2.205 198.965 -1.875 199.295 ;
        RECT -2.205 196.655 -1.875 196.985 ;
        RECT -2.205 195.805 -1.875 196.135 ;
        RECT -2.205 193.495 -1.875 193.825 ;
        RECT -2.205 192.645 -1.875 192.975 ;
        RECT -2.205 190.335 -1.875 190.665 ;
        RECT -2.205 188.755 -1.875 189.085 ;
        RECT -2.205 187.905 -1.875 188.235 ;
        RECT -2.205 185.595 -1.875 185.925 ;
        RECT -2.205 184.745 -1.875 185.075 ;
        RECT -2.205 182.435 -1.875 182.765 ;
        RECT -2.205 181.585 -1.875 181.915 ;
        RECT -2.205 179.275 -1.875 179.605 ;
        RECT -2.205 178.425 -1.875 178.755 ;
        RECT -2.205 176.115 -1.875 176.445 ;
        RECT -2.205 174.535 -1.875 174.865 ;
        RECT -2.205 173.685 -1.875 174.015 ;
        RECT -2.205 171.375 -1.875 171.705 ;
        RECT -2.205 170.525 -1.875 170.855 ;
        RECT -2.205 168.215 -1.875 168.545 ;
        RECT -2.205 167.365 -1.875 167.695 ;
        RECT -2.205 165.055 -1.875 165.385 ;
        RECT -2.205 164.205 -1.875 164.535 ;
        RECT -2.205 161.895 -1.875 162.225 ;
        RECT -2.205 160.315 -1.875 160.645 ;
        RECT -2.205 159.465 -1.875 159.795 ;
        RECT -2.205 157.155 -1.875 157.485 ;
        RECT -2.205 156.305 -1.875 156.635 ;
        RECT -2.205 153.995 -1.875 154.325 ;
        RECT -2.205 153.145 -1.875 153.475 ;
        RECT -2.205 150.835 -1.875 151.165 ;
        RECT -2.205 149.985 -1.875 150.315 ;
        RECT -2.205 147.675 -1.875 148.005 ;
        RECT -2.205 146.095 -1.875 146.425 ;
        RECT -2.205 145.245 -1.875 145.575 ;
        RECT -2.205 142.935 -1.875 143.265 ;
        RECT -2.205 142.085 -1.875 142.415 ;
        RECT -2.205 139.775 -1.875 140.105 ;
        RECT -2.205 138.925 -1.875 139.255 ;
        RECT -2.205 136.615 -1.875 136.945 ;
        RECT -2.205 135.765 -1.875 136.095 ;
        RECT -2.205 133.455 -1.875 133.785 ;
        RECT -2.205 131.875 -1.875 132.205 ;
        RECT -2.205 131.025 -1.875 131.355 ;
        RECT -2.205 128.715 -1.875 129.045 ;
        RECT -2.205 127.865 -1.875 128.195 ;
        RECT -2.205 125.555 -1.875 125.885 ;
        RECT -2.205 124.705 -1.875 125.035 ;
        RECT -2.205 122.395 -1.875 122.725 ;
        RECT -2.205 121.545 -1.875 121.875 ;
        RECT -2.205 119.235 -1.875 119.565 ;
        RECT -2.205 117.655 -1.875 117.985 ;
        RECT -2.205 116.805 -1.875 117.135 ;
        RECT -2.205 114.495 -1.875 114.825 ;
        RECT -2.205 113.645 -1.875 113.975 ;
        RECT -2.205 111.335 -1.875 111.665 ;
        RECT -2.205 110.485 -1.875 110.815 ;
        RECT -2.205 108.175 -1.875 108.505 ;
        RECT -2.205 107.325 -1.875 107.655 ;
        RECT -2.205 105.015 -1.875 105.345 ;
        RECT -2.205 103.435 -1.875 103.765 ;
        RECT -2.205 102.585 -1.875 102.915 ;
        RECT -2.205 100.275 -1.875 100.605 ;
        RECT -2.205 99.425 -1.875 99.755 ;
        RECT -2.205 97.115 -1.875 97.445 ;
        RECT -2.205 96.265 -1.875 96.595 ;
        RECT -2.205 93.955 -1.875 94.285 ;
        RECT -2.205 93.105 -1.875 93.435 ;
        RECT -2.205 90.795 -1.875 91.125 ;
        RECT -2.205 89.215 -1.875 89.545 ;
        RECT -2.205 88.365 -1.875 88.695 ;
        RECT -2.205 86.055 -1.875 86.385 ;
        RECT -2.205 85.205 -1.875 85.535 ;
        RECT -2.205 82.895 -1.875 83.225 ;
        RECT -2.205 82.045 -1.875 82.375 ;
        RECT -2.205 79.735 -1.875 80.065 ;
        RECT -2.205 78.885 -1.875 79.215 ;
        RECT -2.205 76.575 -1.875 76.905 ;
        RECT -2.205 74.995 -1.875 75.325 ;
        RECT -2.205 74.145 -1.875 74.475 ;
        RECT -2.205 71.835 -1.875 72.165 ;
        RECT -2.205 70.985 -1.875 71.315 ;
        RECT -2.205 68.675 -1.875 69.005 ;
        RECT -2.205 67.825 -1.875 68.155 ;
        RECT -2.205 65.515 -1.875 65.845 ;
        RECT -2.205 64.665 -1.875 64.995 ;
        RECT -2.205 62.355 -1.875 62.685 ;
        RECT -2.205 60.775 -1.875 61.105 ;
        RECT -2.205 59.925 -1.875 60.255 ;
        RECT -2.205 57.615 -1.875 57.945 ;
        RECT -2.205 56.765 -1.875 57.095 ;
        RECT -2.205 54.455 -1.875 54.785 ;
        RECT -2.205 53.605 -1.875 53.935 ;
        RECT -2.205 51.295 -1.875 51.625 ;
        RECT -2.205 50.445 -1.875 50.775 ;
        RECT -2.205 48.135 -1.875 48.465 ;
        RECT -2.205 46.555 -1.875 46.885 ;
        RECT -2.205 45.705 -1.875 46.035 ;
        RECT -2.205 43.395 -1.875 43.725 ;
        RECT -2.205 42.545 -1.875 42.875 ;
        RECT -2.205 40.235 -1.875 40.565 ;
        RECT -2.205 39.385 -1.875 39.715 ;
        RECT -2.205 37.075 -1.875 37.405 ;
        RECT -2.205 36.225 -1.875 36.555 ;
        RECT -2.205 33.915 -1.875 34.245 ;
        RECT -2.205 32.335 -1.875 32.665 ;
        RECT -2.205 31.485 -1.875 31.815 ;
        RECT -2.205 29.175 -1.875 29.505 ;
        RECT -2.205 28.325 -1.875 28.655 ;
        RECT -2.205 26.015 -1.875 26.345 ;
        RECT -2.205 25.165 -1.875 25.495 ;
        RECT -2.205 22.855 -1.875 23.185 ;
        RECT -2.205 22.005 -1.875 22.335 ;
        RECT -2.205 19.695 -1.875 20.025 ;
        RECT -2.205 18.115 -1.875 18.445 ;
        RECT -2.205 17.265 -1.875 17.595 ;
        RECT -2.205 14.955 -1.875 15.285 ;
        RECT -2.205 14.105 -1.875 14.435 ;
        RECT -2.205 11.795 -1.875 12.125 ;
        RECT -2.205 10.945 -1.875 11.275 ;
        RECT -2.205 8.635 -1.875 8.965 ;
        RECT -2.205 7.785 -1.875 8.115 ;
        RECT -2.205 5.475 -1.875 5.805 ;
        RECT -2.205 3.895 -1.875 4.225 ;
        RECT -2.205 3.045 -1.875 3.375 ;
        RECT -2.205 0.87 -1.875 1.2 ;
        RECT -2.205 -0.845 -1.875 -0.515 ;
        RECT -2.205 -2.205 -1.875 -1.875 ;
        RECT -2.205 -3.565 -1.875 -3.235 ;
        RECT -2.205 -4.925 -1.875 -4.595 ;
        RECT -2.205 -6.285 -1.875 -5.955 ;
        RECT -2.205 -7.645 -1.875 -7.315 ;
        RECT -2.205 -9.005 -1.875 -8.675 ;
        RECT -2.205 -10.365 -1.875 -10.035 ;
        RECT -2.205 -11.725 -1.875 -11.395 ;
        RECT -2.205 -13.085 -1.875 -12.755 ;
        RECT -2.205 -14.445 -1.875 -14.115 ;
        RECT -2.205 -15.805 -1.875 -15.475 ;
        RECT -2.205 -17.165 -1.875 -16.835 ;
        RECT -2.205 -21.245 -1.875 -20.915 ;
        RECT -2.205 -22.605 -1.875 -22.275 ;
        RECT -2.205 -23.965 -1.875 -23.635 ;
        RECT -2.205 -25.325 -1.875 -24.995 ;
        RECT -2.205 -26.685 -1.875 -26.355 ;
        RECT -2.205 -28.045 -1.875 -27.715 ;
        RECT -2.205 -29.405 -1.875 -29.075 ;
        RECT -2.205 -30.765 -1.875 -30.435 ;
        RECT -2.205 -32.125 -1.875 -31.795 ;
        RECT -2.205 -33.485 -1.875 -33.155 ;
        RECT -2.205 -36.205 -1.875 -35.875 ;
        RECT -2.205 -37.565 -1.875 -37.235 ;
        RECT -2.205 -38.925 -1.875 -38.595 ;
        RECT -2.205 -40.285 -1.875 -39.955 ;
        RECT -2.205 -41.645 -1.875 -41.315 ;
        RECT -2.205 -43.005 -1.875 -42.675 ;
        RECT -2.205 -44.365 -1.875 -44.035 ;
        RECT -2.205 -45.725 -1.875 -45.395 ;
        RECT -2.205 -47.085 -1.875 -46.755 ;
        RECT -2.205 -48.445 -1.875 -48.115 ;
        RECT -2.205 -51.165 -1.875 -50.835 ;
        RECT -2.205 -52.525 -1.875 -52.195 ;
        RECT -2.205 -53.885 -1.875 -53.555 ;
        RECT -2.205 -55.245 -1.875 -54.915 ;
        RECT -2.205 -56.605 -1.875 -56.275 ;
        RECT -2.205 -57.965 -1.875 -57.635 ;
        RECT -2.205 -59.325 -1.875 -58.995 ;
        RECT -2.205 -60.685 -1.875 -60.355 ;
        RECT -2.205 -62.045 -1.875 -61.715 ;
        RECT -2.205 -63.405 -1.875 -63.075 ;
        RECT -2.205 -64.765 -1.875 -64.435 ;
        RECT -2.205 -66.125 -1.875 -65.795 ;
        RECT -2.205 -67.485 -1.875 -67.155 ;
        RECT -2.205 -68.845 -1.875 -68.515 ;
        RECT -2.205 -70.205 -1.875 -69.875 ;
        RECT -2.205 -71.565 -1.875 -71.235 ;
        RECT -2.205 -72.925 -1.875 -72.595 ;
        RECT -2.205 -74.285 -1.875 -73.955 ;
        RECT -2.205 -75.645 -1.875 -75.315 ;
        RECT -2.205 -77.005 -1.875 -76.675 ;
        RECT -2.205 -78.365 -1.875 -78.035 ;
        RECT -2.205 -79.725 -1.875 -79.395 ;
        RECT -2.205 -81.085 -1.875 -80.755 ;
        RECT -2.205 -82.445 -1.875 -82.115 ;
        RECT -2.205 -83.805 -1.875 -83.475 ;
        RECT -2.205 -85.165 -1.875 -84.835 ;
        RECT -2.205 -87.885 -1.875 -87.555 ;
        RECT -2.205 -89.245 -1.875 -88.915 ;
        RECT -2.205 -90.605 -1.875 -90.275 ;
        RECT -2.205 -91.965 -1.875 -91.635 ;
        RECT -2.205 -93.325 -1.875 -92.995 ;
        RECT -2.205 -94.685 -1.875 -94.355 ;
        RECT -2.205 -96.045 -1.875 -95.715 ;
        RECT -2.205 -97.405 -1.875 -97.075 ;
        RECT -2.205 -98.765 -1.875 -98.435 ;
        RECT -2.205 -100.125 -1.875 -99.795 ;
        RECT -2.205 -101.485 -1.875 -101.155 ;
        RECT -2.205 -102.845 -1.875 -102.515 ;
        RECT -2.205 -104.205 -1.875 -103.875 ;
        RECT -2.205 -105.565 -1.875 -105.235 ;
        RECT -2.205 -106.925 -1.875 -106.595 ;
        RECT -2.205 -108.285 -1.875 -107.955 ;
        RECT -2.205 -109.645 -1.875 -109.315 ;
        RECT -2.205 -111.005 -1.875 -110.675 ;
        RECT -2.205 -112.365 -1.875 -112.035 ;
        RECT -2.205 -113.725 -1.875 -113.395 ;
        RECT -2.205 -115.085 -1.875 -114.755 ;
        RECT -2.205 -116.445 -1.875 -116.115 ;
        RECT -2.205 -117.805 -1.875 -117.475 ;
        RECT -2.205 -119.165 -1.875 -118.835 ;
        RECT -2.205 -120.525 -1.875 -120.195 ;
        RECT -2.205 -121.885 -1.875 -121.555 ;
        RECT -2.205 -123.245 -1.875 -122.915 ;
        RECT -2.205 -124.605 -1.875 -124.275 ;
        RECT -2.205 -125.965 -1.875 -125.635 ;
        RECT -2.205 -127.325 -1.875 -126.995 ;
        RECT -2.205 -128.685 -1.875 -128.355 ;
        RECT -2.205 -130.045 -1.875 -129.715 ;
        RECT -2.205 -131.405 -1.875 -131.075 ;
        RECT -2.205 -132.765 -1.875 -132.435 ;
        RECT -2.205 -134.125 -1.875 -133.795 ;
        RECT -2.205 -135.485 -1.875 -135.155 ;
        RECT -2.205 -136.845 -1.875 -136.515 ;
        RECT -2.205 -138.205 -1.875 -137.875 ;
        RECT -2.205 -139.565 -1.875 -139.235 ;
        RECT -2.205 -140.925 -1.875 -140.595 ;
        RECT -2.205 -142.285 -1.875 -141.955 ;
        RECT -2.205 -143.645 -1.875 -143.315 ;
        RECT -2.205 -145.005 -1.875 -144.675 ;
        RECT -2.205 -146.365 -1.875 -146.035 ;
        RECT -2.205 -147.725 -1.875 -147.395 ;
        RECT -2.205 -149.085 -1.875 -148.755 ;
        RECT -2.205 -150.445 -1.875 -150.115 ;
        RECT -2.205 -151.805 -1.875 -151.475 ;
        RECT -2.205 -153.165 -1.875 -152.835 ;
        RECT -2.205 -154.525 -1.875 -154.195 ;
        RECT -2.205 -155.885 -1.875 -155.555 ;
        RECT -2.205 -157.245 -1.875 -156.915 ;
        RECT -2.205 -158.605 -1.875 -158.275 ;
        RECT -2.205 -159.965 -1.875 -159.635 ;
        RECT -2.205 -161.325 -1.875 -160.995 ;
        RECT -2.205 -162.685 -1.875 -162.355 ;
        RECT -2.205 -164.045 -1.875 -163.715 ;
        RECT -2.205 -165.405 -1.875 -165.075 ;
        RECT -2.205 -166.765 -1.875 -166.435 ;
        RECT -2.205 -168.125 -1.875 -167.795 ;
        RECT -2.205 -169.485 -1.875 -169.155 ;
        RECT -2.205 -170.845 -1.875 -170.515 ;
        RECT -2.205 -172.205 -1.875 -171.875 ;
        RECT -2.205 -173.565 -1.875 -173.235 ;
        RECT -2.205 -174.925 -1.875 -174.595 ;
        RECT -2.205 -176.285 -1.875 -175.955 ;
        RECT -2.205 -177.645 -1.875 -177.315 ;
        RECT -2.205 -183.29 -1.875 -182.16 ;
        RECT -2.2 -183.405 -1.88 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -0.845 244.04 -0.515 245.17 ;
        RECT -0.845 239.875 -0.515 240.205 ;
        RECT -0.845 238.515 -0.515 238.845 ;
        RECT -0.845 237.155 -0.515 237.485 ;
        RECT -0.845 235.17 -0.515 235.5 ;
        RECT -0.845 232.995 -0.515 233.325 ;
        RECT -0.845 231.415 -0.515 231.745 ;
        RECT -0.845 230.565 -0.515 230.895 ;
        RECT -0.845 228.255 -0.515 228.585 ;
        RECT -0.845 227.405 -0.515 227.735 ;
        RECT -0.845 225.095 -0.515 225.425 ;
        RECT -0.845 224.245 -0.515 224.575 ;
        RECT -0.845 221.935 -0.515 222.265 ;
        RECT -0.845 221.085 -0.515 221.415 ;
        RECT -0.845 218.775 -0.515 219.105 ;
        RECT -0.845 217.195 -0.515 217.525 ;
        RECT -0.845 216.345 -0.515 216.675 ;
        RECT -0.845 214.035 -0.515 214.365 ;
        RECT -0.845 213.185 -0.515 213.515 ;
        RECT -0.845 210.875 -0.515 211.205 ;
        RECT -0.845 210.025 -0.515 210.355 ;
        RECT -0.845 207.715 -0.515 208.045 ;
        RECT -0.845 206.865 -0.515 207.195 ;
        RECT -0.845 204.555 -0.515 204.885 ;
        RECT -0.845 202.975 -0.515 203.305 ;
        RECT -0.845 202.125 -0.515 202.455 ;
        RECT -0.845 199.815 -0.515 200.145 ;
        RECT -0.845 198.965 -0.515 199.295 ;
        RECT -0.845 196.655 -0.515 196.985 ;
        RECT -0.845 195.805 -0.515 196.135 ;
        RECT -0.845 193.495 -0.515 193.825 ;
        RECT -0.845 192.645 -0.515 192.975 ;
        RECT -0.845 190.335 -0.515 190.665 ;
        RECT -0.845 188.755 -0.515 189.085 ;
        RECT -0.845 187.905 -0.515 188.235 ;
        RECT -0.845 185.595 -0.515 185.925 ;
        RECT -0.845 184.745 -0.515 185.075 ;
        RECT -0.845 182.435 -0.515 182.765 ;
        RECT -0.845 181.585 -0.515 181.915 ;
        RECT -0.845 179.275 -0.515 179.605 ;
        RECT -0.845 178.425 -0.515 178.755 ;
        RECT -0.845 176.115 -0.515 176.445 ;
        RECT -0.845 174.535 -0.515 174.865 ;
        RECT -0.845 173.685 -0.515 174.015 ;
        RECT -0.845 171.375 -0.515 171.705 ;
        RECT -0.845 170.525 -0.515 170.855 ;
        RECT -0.845 168.215 -0.515 168.545 ;
        RECT -0.845 167.365 -0.515 167.695 ;
        RECT -0.845 165.055 -0.515 165.385 ;
        RECT -0.845 164.205 -0.515 164.535 ;
        RECT -0.845 161.895 -0.515 162.225 ;
        RECT -0.845 160.315 -0.515 160.645 ;
        RECT -0.845 159.465 -0.515 159.795 ;
        RECT -0.845 157.155 -0.515 157.485 ;
        RECT -0.845 156.305 -0.515 156.635 ;
        RECT -0.845 153.995 -0.515 154.325 ;
        RECT -0.845 153.145 -0.515 153.475 ;
        RECT -0.845 150.835 -0.515 151.165 ;
        RECT -0.845 149.985 -0.515 150.315 ;
        RECT -0.845 147.675 -0.515 148.005 ;
        RECT -0.845 146.095 -0.515 146.425 ;
        RECT -0.845 145.245 -0.515 145.575 ;
        RECT -0.845 142.935 -0.515 143.265 ;
        RECT -0.845 142.085 -0.515 142.415 ;
        RECT -0.845 139.775 -0.515 140.105 ;
        RECT -0.845 138.925 -0.515 139.255 ;
        RECT -0.845 136.615 -0.515 136.945 ;
        RECT -0.845 135.765 -0.515 136.095 ;
        RECT -0.845 133.455 -0.515 133.785 ;
        RECT -0.845 131.875 -0.515 132.205 ;
        RECT -0.845 131.025 -0.515 131.355 ;
        RECT -0.845 128.715 -0.515 129.045 ;
        RECT -0.845 127.865 -0.515 128.195 ;
        RECT -0.845 125.555 -0.515 125.885 ;
        RECT -0.845 124.705 -0.515 125.035 ;
        RECT -0.845 122.395 -0.515 122.725 ;
        RECT -0.845 121.545 -0.515 121.875 ;
        RECT -0.845 119.235 -0.515 119.565 ;
        RECT -0.845 117.655 -0.515 117.985 ;
        RECT -0.845 116.805 -0.515 117.135 ;
        RECT -0.845 114.495 -0.515 114.825 ;
        RECT -0.845 113.645 -0.515 113.975 ;
        RECT -0.845 111.335 -0.515 111.665 ;
        RECT -0.845 110.485 -0.515 110.815 ;
        RECT -0.845 108.175 -0.515 108.505 ;
        RECT -0.845 107.325 -0.515 107.655 ;
        RECT -0.845 105.015 -0.515 105.345 ;
        RECT -0.845 103.435 -0.515 103.765 ;
        RECT -0.845 102.585 -0.515 102.915 ;
        RECT -0.845 100.275 -0.515 100.605 ;
        RECT -0.845 99.425 -0.515 99.755 ;
        RECT -0.845 97.115 -0.515 97.445 ;
        RECT -0.845 96.265 -0.515 96.595 ;
        RECT -0.845 93.955 -0.515 94.285 ;
        RECT -0.845 93.105 -0.515 93.435 ;
        RECT -0.845 90.795 -0.515 91.125 ;
        RECT -0.845 89.215 -0.515 89.545 ;
        RECT -0.845 88.365 -0.515 88.695 ;
        RECT -0.845 86.055 -0.515 86.385 ;
        RECT -0.845 85.205 -0.515 85.535 ;
        RECT -0.845 82.895 -0.515 83.225 ;
        RECT -0.845 82.045 -0.515 82.375 ;
        RECT -0.845 79.735 -0.515 80.065 ;
        RECT -0.845 78.885 -0.515 79.215 ;
        RECT -0.845 76.575 -0.515 76.905 ;
        RECT -0.845 74.995 -0.515 75.325 ;
        RECT -0.845 74.145 -0.515 74.475 ;
        RECT -0.845 71.835 -0.515 72.165 ;
        RECT -0.845 70.985 -0.515 71.315 ;
        RECT -0.845 68.675 -0.515 69.005 ;
        RECT -0.845 67.825 -0.515 68.155 ;
        RECT -0.845 65.515 -0.515 65.845 ;
        RECT -0.845 64.665 -0.515 64.995 ;
        RECT -0.845 62.355 -0.515 62.685 ;
        RECT -0.845 60.775 -0.515 61.105 ;
        RECT -0.845 59.925 -0.515 60.255 ;
        RECT -0.845 57.615 -0.515 57.945 ;
        RECT -0.845 56.765 -0.515 57.095 ;
        RECT -0.845 54.455 -0.515 54.785 ;
        RECT -0.845 53.605 -0.515 53.935 ;
        RECT -0.845 51.295 -0.515 51.625 ;
        RECT -0.845 50.445 -0.515 50.775 ;
        RECT -0.845 48.135 -0.515 48.465 ;
        RECT -0.845 46.555 -0.515 46.885 ;
        RECT -0.845 45.705 -0.515 46.035 ;
        RECT -0.845 43.395 -0.515 43.725 ;
        RECT -0.845 42.545 -0.515 42.875 ;
        RECT -0.845 40.235 -0.515 40.565 ;
        RECT -0.845 39.385 -0.515 39.715 ;
        RECT -0.845 37.075 -0.515 37.405 ;
        RECT -0.845 36.225 -0.515 36.555 ;
        RECT -0.845 33.915 -0.515 34.245 ;
        RECT -0.845 32.335 -0.515 32.665 ;
        RECT -0.845 31.485 -0.515 31.815 ;
        RECT -0.845 29.175 -0.515 29.505 ;
        RECT -0.845 28.325 -0.515 28.655 ;
        RECT -0.845 26.015 -0.515 26.345 ;
        RECT -0.845 25.165 -0.515 25.495 ;
        RECT -0.845 22.855 -0.515 23.185 ;
        RECT -0.845 22.005 -0.515 22.335 ;
        RECT -0.845 19.695 -0.515 20.025 ;
        RECT -0.845 18.115 -0.515 18.445 ;
        RECT -0.845 17.265 -0.515 17.595 ;
        RECT -0.845 14.955 -0.515 15.285 ;
        RECT -0.845 14.105 -0.515 14.435 ;
        RECT -0.845 11.795 -0.515 12.125 ;
        RECT -0.845 10.945 -0.515 11.275 ;
        RECT -0.845 8.635 -0.515 8.965 ;
        RECT -0.845 7.785 -0.515 8.115 ;
        RECT -0.845 5.475 -0.515 5.805 ;
        RECT -0.845 3.895 -0.515 4.225 ;
        RECT -0.845 3.045 -0.515 3.375 ;
        RECT -0.845 0.87 -0.515 1.2 ;
        RECT -0.845 -0.845 -0.515 -0.515 ;
        RECT -0.845 -2.205 -0.515 -1.875 ;
        RECT -0.845 -3.565 -0.515 -3.235 ;
        RECT -0.845 -4.925 -0.515 -4.595 ;
        RECT -0.845 -6.285 -0.515 -5.955 ;
        RECT -0.845 -7.645 -0.515 -7.315 ;
        RECT -0.845 -9.005 -0.515 -8.675 ;
        RECT -0.845 -10.365 -0.515 -10.035 ;
        RECT -0.845 -13.085 -0.515 -12.755 ;
        RECT -0.845 -14.445 -0.515 -14.115 ;
        RECT -0.845 -15.805 -0.515 -15.475 ;
        RECT -0.845 -17.165 -0.515 -16.835 ;
        RECT -0.845 -21.245 -0.515 -20.915 ;
        RECT -0.845 -22.605 -0.515 -22.275 ;
        RECT -0.845 -23.965 -0.515 -23.635 ;
        RECT -0.845 -25.325 -0.515 -24.995 ;
        RECT -0.845 -26.685 -0.515 -26.355 ;
        RECT -0.845 -28.045 -0.515 -27.715 ;
        RECT -0.845 -29.405 -0.515 -29.075 ;
        RECT -0.845 -30.765 -0.515 -30.435 ;
        RECT -0.845 -32.125 -0.515 -31.795 ;
        RECT -0.845 -33.485 -0.515 -33.155 ;
        RECT -0.845 -36.205 -0.515 -35.875 ;
        RECT -0.845 -37.565 -0.515 -37.235 ;
        RECT -0.845 -38.925 -0.515 -38.595 ;
        RECT -0.845 -40.285 -0.515 -39.955 ;
        RECT -0.845 -41.645 -0.515 -41.315 ;
        RECT -0.845 -43.005 -0.515 -42.675 ;
        RECT -0.845 -44.365 -0.515 -44.035 ;
        RECT -0.845 -45.725 -0.515 -45.395 ;
        RECT -0.845 -47.085 -0.515 -46.755 ;
        RECT -0.845 -48.445 -0.515 -48.115 ;
        RECT -0.845 -51.165 -0.515 -50.835 ;
        RECT -0.845 -52.525 -0.515 -52.195 ;
        RECT -0.845 -53.885 -0.515 -53.555 ;
        RECT -0.845 -55.245 -0.515 -54.915 ;
        RECT -0.845 -56.605 -0.515 -56.275 ;
        RECT -0.845 -57.965 -0.515 -57.635 ;
        RECT -0.845 -59.325 -0.515 -58.995 ;
        RECT -0.845 -60.685 -0.515 -60.355 ;
        RECT -0.845 -62.045 -0.515 -61.715 ;
        RECT -0.845 -63.405 -0.515 -63.075 ;
        RECT -0.845 -64.765 -0.515 -64.435 ;
        RECT -0.845 -66.125 -0.515 -65.795 ;
        RECT -0.845 -67.485 -0.515 -67.155 ;
        RECT -0.845 -68.845 -0.515 -68.515 ;
        RECT -0.845 -70.205 -0.515 -69.875 ;
        RECT -0.845 -71.565 -0.515 -71.235 ;
        RECT -0.845 -72.925 -0.515 -72.595 ;
        RECT -0.845 -74.285 -0.515 -73.955 ;
        RECT -0.845 -75.645 -0.515 -75.315 ;
        RECT -0.845 -77.005 -0.515 -76.675 ;
        RECT -0.845 -78.365 -0.515 -78.035 ;
        RECT -0.845 -79.725 -0.515 -79.395 ;
        RECT -0.845 -81.085 -0.515 -80.755 ;
        RECT -0.845 -82.445 -0.515 -82.115 ;
        RECT -0.845 -83.805 -0.515 -83.475 ;
        RECT -0.845 -85.165 -0.515 -84.835 ;
        RECT -0.845 -87.885 -0.515 -87.555 ;
        RECT -0.845 -89.245 -0.515 -88.915 ;
        RECT -0.845 -90.605 -0.515 -90.275 ;
        RECT -0.845 -91.965 -0.515 -91.635 ;
        RECT -0.845 -93.325 -0.515 -92.995 ;
        RECT -0.845 -94.685 -0.515 -94.355 ;
        RECT -0.845 -96.045 -0.515 -95.715 ;
        RECT -0.845 -97.405 -0.515 -97.075 ;
        RECT -0.845 -98.765 -0.515 -98.435 ;
        RECT -0.845 -100.125 -0.515 -99.795 ;
        RECT -0.845 -101.485 -0.515 -101.155 ;
        RECT -0.845 -102.845 -0.515 -102.515 ;
        RECT -0.845 -104.205 -0.515 -103.875 ;
        RECT -0.845 -105.565 -0.515 -105.235 ;
        RECT -0.845 -106.925 -0.515 -106.595 ;
        RECT -0.845 -108.285 -0.515 -107.955 ;
        RECT -0.845 -109.645 -0.515 -109.315 ;
        RECT -0.845 -111.005 -0.515 -110.675 ;
        RECT -0.845 -112.365 -0.515 -112.035 ;
        RECT -0.845 -113.725 -0.515 -113.395 ;
        RECT -0.845 -115.085 -0.515 -114.755 ;
        RECT -0.845 -116.445 -0.515 -116.115 ;
        RECT -0.845 -117.805 -0.515 -117.475 ;
        RECT -0.845 -119.165 -0.515 -118.835 ;
        RECT -0.845 -120.525 -0.515 -120.195 ;
        RECT -0.845 -121.885 -0.515 -121.555 ;
        RECT -0.845 -123.245 -0.515 -122.915 ;
        RECT -0.845 -124.605 -0.515 -124.275 ;
        RECT -0.845 -125.965 -0.515 -125.635 ;
        RECT -0.845 -127.325 -0.515 -126.995 ;
        RECT -0.845 -128.685 -0.515 -128.355 ;
        RECT -0.845 -130.045 -0.515 -129.715 ;
        RECT -0.845 -131.405 -0.515 -131.075 ;
        RECT -0.845 -132.765 -0.515 -132.435 ;
        RECT -0.845 -134.125 -0.515 -133.795 ;
        RECT -0.845 -135.485 -0.515 -135.155 ;
        RECT -0.845 -136.845 -0.515 -136.515 ;
        RECT -0.845 -138.205 -0.515 -137.875 ;
        RECT -0.845 -139.565 -0.515 -139.235 ;
        RECT -0.845 -140.925 -0.515 -140.595 ;
        RECT -0.845 -142.285 -0.515 -141.955 ;
        RECT -0.845 -143.645 -0.515 -143.315 ;
        RECT -0.845 -145.005 -0.515 -144.675 ;
        RECT -0.845 -146.365 -0.515 -146.035 ;
        RECT -0.845 -147.725 -0.515 -147.395 ;
        RECT -0.845 -149.085 -0.515 -148.755 ;
        RECT -0.845 -150.445 -0.515 -150.115 ;
        RECT -0.845 -151.805 -0.515 -151.475 ;
        RECT -0.845 -153.165 -0.515 -152.835 ;
        RECT -0.845 -154.525 -0.515 -154.195 ;
        RECT -0.845 -155.885 -0.515 -155.555 ;
        RECT -0.845 -157.245 -0.515 -156.915 ;
        RECT -0.845 -158.605 -0.515 -158.275 ;
        RECT -0.845 -159.965 -0.515 -159.635 ;
        RECT -0.845 -161.325 -0.515 -160.995 ;
        RECT -0.845 -162.685 -0.515 -162.355 ;
        RECT -0.845 -164.045 -0.515 -163.715 ;
        RECT -0.845 -165.405 -0.515 -165.075 ;
        RECT -0.845 -166.765 -0.515 -166.435 ;
        RECT -0.845 -168.125 -0.515 -167.795 ;
        RECT -0.845 -169.485 -0.515 -169.155 ;
        RECT -0.845 -170.845 -0.515 -170.515 ;
        RECT -0.845 -172.205 -0.515 -171.875 ;
        RECT -0.845 -173.565 -0.515 -173.235 ;
        RECT -0.845 -174.925 -0.515 -174.595 ;
        RECT -0.845 -176.285 -0.515 -175.955 ;
        RECT -0.845 -177.645 -0.515 -177.315 ;
        RECT -0.845 -183.29 -0.515 -182.16 ;
        RECT -0.84 -183.405 -0.52 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.515 244.04 0.845 245.17 ;
        RECT 0.515 239.875 0.845 240.205 ;
        RECT 0.515 238.515 0.845 238.845 ;
        RECT 0.515 237.155 0.845 237.485 ;
        RECT 0.52 237.155 0.84 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.515 -0.845 0.845 -0.515 ;
        RECT 0.515 -2.205 0.845 -1.875 ;
        RECT 0.515 -3.565 0.845 -3.235 ;
        RECT 0.52 -3.565 0.84 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.515 -91.965 0.845 -91.635 ;
        RECT 0.515 -93.325 0.845 -92.995 ;
        RECT 0.515 -94.685 0.845 -94.355 ;
        RECT 0.515 -96.045 0.845 -95.715 ;
        RECT 0.515 -97.405 0.845 -97.075 ;
        RECT 0.515 -98.765 0.845 -98.435 ;
        RECT 0.515 -100.125 0.845 -99.795 ;
        RECT 0.515 -101.485 0.845 -101.155 ;
        RECT 0.515 -102.845 0.845 -102.515 ;
        RECT 0.515 -104.205 0.845 -103.875 ;
        RECT 0.515 -105.565 0.845 -105.235 ;
        RECT 0.515 -106.925 0.845 -106.595 ;
        RECT 0.515 -108.285 0.845 -107.955 ;
        RECT 0.515 -109.645 0.845 -109.315 ;
        RECT 0.515 -111.005 0.845 -110.675 ;
        RECT 0.515 -112.365 0.845 -112.035 ;
        RECT 0.515 -113.725 0.845 -113.395 ;
        RECT 0.515 -115.085 0.845 -114.755 ;
        RECT 0.515 -116.445 0.845 -116.115 ;
        RECT 0.515 -117.805 0.845 -117.475 ;
        RECT 0.515 -119.165 0.845 -118.835 ;
        RECT 0.515 -120.525 0.845 -120.195 ;
        RECT 0.515 -121.885 0.845 -121.555 ;
        RECT 0.515 -123.245 0.845 -122.915 ;
        RECT 0.515 -124.605 0.845 -124.275 ;
        RECT 0.515 -125.965 0.845 -125.635 ;
        RECT 0.515 -127.325 0.845 -126.995 ;
        RECT 0.515 -128.685 0.845 -128.355 ;
        RECT 0.515 -130.045 0.845 -129.715 ;
        RECT 0.515 -131.405 0.845 -131.075 ;
        RECT 0.515 -132.765 0.845 -132.435 ;
        RECT 0.515 -134.125 0.845 -133.795 ;
        RECT 0.515 -135.485 0.845 -135.155 ;
        RECT 0.515 -136.845 0.845 -136.515 ;
        RECT 0.515 -138.205 0.845 -137.875 ;
        RECT 0.515 -139.565 0.845 -139.235 ;
        RECT 0.515 -140.925 0.845 -140.595 ;
        RECT 0.515 -142.285 0.845 -141.955 ;
        RECT 0.515 -143.645 0.845 -143.315 ;
        RECT 0.515 -145.005 0.845 -144.675 ;
        RECT 0.515 -146.365 0.845 -146.035 ;
        RECT 0.515 -147.725 0.845 -147.395 ;
        RECT 0.515 -149.085 0.845 -148.755 ;
        RECT 0.515 -150.445 0.845 -150.115 ;
        RECT 0.515 -151.805 0.845 -151.475 ;
        RECT 0.515 -153.165 0.845 -152.835 ;
        RECT 0.515 -154.525 0.845 -154.195 ;
        RECT 0.515 -155.885 0.845 -155.555 ;
        RECT 0.515 -157.245 0.845 -156.915 ;
        RECT 0.515 -158.605 0.845 -158.275 ;
        RECT 0.515 -159.965 0.845 -159.635 ;
        RECT 0.515 -161.325 0.845 -160.995 ;
        RECT 0.515 -162.685 0.845 -162.355 ;
        RECT 0.515 -164.045 0.845 -163.715 ;
        RECT 0.515 -165.405 0.845 -165.075 ;
        RECT 0.515 -166.765 0.845 -166.435 ;
        RECT 0.515 -168.125 0.845 -167.795 ;
        RECT 0.515 -169.485 0.845 -169.155 ;
        RECT 0.515 -170.845 0.845 -170.515 ;
        RECT 0.515 -172.205 0.845 -171.875 ;
        RECT 0.515 -173.565 0.845 -173.235 ;
        RECT 0.515 -174.925 0.845 -174.595 ;
        RECT 0.515 -176.285 0.845 -175.955 ;
        RECT 0.515 -177.645 0.845 -177.315 ;
        RECT 0.515 -183.29 0.845 -182.16 ;
        RECT 0.52 -183.405 0.84 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.875 244.04 2.205 245.17 ;
        RECT 1.875 239.875 2.205 240.205 ;
        RECT 1.875 238.515 2.205 238.845 ;
        RECT 1.875 237.155 2.205 237.485 ;
        RECT 1.88 237.155 2.2 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.875 -0.845 2.205 -0.515 ;
        RECT 1.875 -2.205 2.205 -1.875 ;
        RECT 1.875 -3.565 2.205 -3.235 ;
        RECT 1.88 -3.565 2.2 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.875 -91.965 2.205 -91.635 ;
        RECT 1.875 -93.325 2.205 -92.995 ;
        RECT 1.875 -94.685 2.205 -94.355 ;
        RECT 1.875 -96.045 2.205 -95.715 ;
        RECT 1.875 -97.405 2.205 -97.075 ;
        RECT 1.875 -98.765 2.205 -98.435 ;
        RECT 1.875 -100.125 2.205 -99.795 ;
        RECT 1.875 -101.485 2.205 -101.155 ;
        RECT 1.875 -102.845 2.205 -102.515 ;
        RECT 1.875 -104.205 2.205 -103.875 ;
        RECT 1.875 -105.565 2.205 -105.235 ;
        RECT 1.875 -106.925 2.205 -106.595 ;
        RECT 1.875 -108.285 2.205 -107.955 ;
        RECT 1.875 -109.645 2.205 -109.315 ;
        RECT 1.875 -111.005 2.205 -110.675 ;
        RECT 1.875 -112.365 2.205 -112.035 ;
        RECT 1.875 -113.725 2.205 -113.395 ;
        RECT 1.875 -115.085 2.205 -114.755 ;
        RECT 1.875 -116.445 2.205 -116.115 ;
        RECT 1.875 -117.805 2.205 -117.475 ;
        RECT 1.875 -119.165 2.205 -118.835 ;
        RECT 1.875 -120.525 2.205 -120.195 ;
        RECT 1.875 -121.885 2.205 -121.555 ;
        RECT 1.875 -123.245 2.205 -122.915 ;
        RECT 1.875 -124.605 2.205 -124.275 ;
        RECT 1.875 -125.965 2.205 -125.635 ;
        RECT 1.875 -127.325 2.205 -126.995 ;
        RECT 1.875 -128.685 2.205 -128.355 ;
        RECT 1.875 -130.045 2.205 -129.715 ;
        RECT 1.875 -131.405 2.205 -131.075 ;
        RECT 1.875 -132.765 2.205 -132.435 ;
        RECT 1.875 -134.125 2.205 -133.795 ;
        RECT 1.875 -135.485 2.205 -135.155 ;
        RECT 1.875 -136.845 2.205 -136.515 ;
        RECT 1.875 -138.205 2.205 -137.875 ;
        RECT 1.875 -139.565 2.205 -139.235 ;
        RECT 1.875 -140.925 2.205 -140.595 ;
        RECT 1.875 -142.285 2.205 -141.955 ;
        RECT 1.875 -143.645 2.205 -143.315 ;
        RECT 1.875 -145.005 2.205 -144.675 ;
        RECT 1.875 -146.365 2.205 -146.035 ;
        RECT 1.875 -147.725 2.205 -147.395 ;
        RECT 1.875 -149.085 2.205 -148.755 ;
        RECT 1.875 -150.445 2.205 -150.115 ;
        RECT 1.875 -151.805 2.205 -151.475 ;
        RECT 1.875 -153.165 2.205 -152.835 ;
        RECT 1.875 -154.525 2.205 -154.195 ;
        RECT 1.875 -155.885 2.205 -155.555 ;
        RECT 1.875 -157.245 2.205 -156.915 ;
        RECT 1.875 -158.605 2.205 -158.275 ;
        RECT 1.875 -159.965 2.205 -159.635 ;
        RECT 1.875 -161.325 2.205 -160.995 ;
        RECT 1.875 -162.685 2.205 -162.355 ;
        RECT 1.875 -164.045 2.205 -163.715 ;
        RECT 1.875 -165.405 2.205 -165.075 ;
        RECT 1.875 -166.765 2.205 -166.435 ;
        RECT 1.875 -168.125 2.205 -167.795 ;
        RECT 1.875 -169.485 2.205 -169.155 ;
        RECT 1.875 -170.845 2.205 -170.515 ;
        RECT 1.875 -172.205 2.205 -171.875 ;
        RECT 1.875 -173.565 2.205 -173.235 ;
        RECT 1.875 -174.925 2.205 -174.595 ;
        RECT 1.875 -176.285 2.205 -175.955 ;
        RECT 1.875 -177.645 2.205 -177.315 ;
        RECT 1.875 -183.29 2.205 -182.16 ;
        RECT 1.88 -183.405 2.2 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.66 -94.075 2.99 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.235 244.04 3.565 245.17 ;
        RECT 3.235 239.875 3.565 240.205 ;
        RECT 3.235 238.515 3.565 238.845 ;
        RECT 3.235 237.155 3.565 237.485 ;
        RECT 3.24 237.155 3.56 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.235 -96.045 3.565 -95.715 ;
        RECT 3.235 -97.405 3.565 -97.075 ;
        RECT 3.235 -98.765 3.565 -98.435 ;
        RECT 3.235 -100.125 3.565 -99.795 ;
        RECT 3.235 -101.485 3.565 -101.155 ;
        RECT 3.235 -102.845 3.565 -102.515 ;
        RECT 3.235 -104.205 3.565 -103.875 ;
        RECT 3.235 -105.565 3.565 -105.235 ;
        RECT 3.235 -106.925 3.565 -106.595 ;
        RECT 3.235 -108.285 3.565 -107.955 ;
        RECT 3.235 -109.645 3.565 -109.315 ;
        RECT 3.235 -111.005 3.565 -110.675 ;
        RECT 3.235 -112.365 3.565 -112.035 ;
        RECT 3.235 -113.725 3.565 -113.395 ;
        RECT 3.235 -115.085 3.565 -114.755 ;
        RECT 3.235 -116.445 3.565 -116.115 ;
        RECT 3.235 -117.805 3.565 -117.475 ;
        RECT 3.235 -119.165 3.565 -118.835 ;
        RECT 3.235 -120.525 3.565 -120.195 ;
        RECT 3.235 -121.885 3.565 -121.555 ;
        RECT 3.235 -123.245 3.565 -122.915 ;
        RECT 3.235 -124.605 3.565 -124.275 ;
        RECT 3.235 -125.965 3.565 -125.635 ;
        RECT 3.235 -127.325 3.565 -126.995 ;
        RECT 3.235 -128.685 3.565 -128.355 ;
        RECT 3.235 -130.045 3.565 -129.715 ;
        RECT 3.235 -131.405 3.565 -131.075 ;
        RECT 3.235 -132.765 3.565 -132.435 ;
        RECT 3.235 -134.125 3.565 -133.795 ;
        RECT 3.235 -135.485 3.565 -135.155 ;
        RECT 3.235 -136.845 3.565 -136.515 ;
        RECT 3.235 -138.205 3.565 -137.875 ;
        RECT 3.235 -139.565 3.565 -139.235 ;
        RECT 3.235 -140.925 3.565 -140.595 ;
        RECT 3.235 -142.285 3.565 -141.955 ;
        RECT 3.235 -143.645 3.565 -143.315 ;
        RECT 3.235 -145.005 3.565 -144.675 ;
        RECT 3.235 -146.365 3.565 -146.035 ;
        RECT 3.235 -147.725 3.565 -147.395 ;
        RECT 3.235 -149.085 3.565 -148.755 ;
        RECT 3.235 -150.445 3.565 -150.115 ;
        RECT 3.235 -151.805 3.565 -151.475 ;
        RECT 3.235 -153.165 3.565 -152.835 ;
        RECT 3.235 -154.525 3.565 -154.195 ;
        RECT 3.235 -155.885 3.565 -155.555 ;
        RECT 3.235 -157.245 3.565 -156.915 ;
        RECT 3.235 -158.605 3.565 -158.275 ;
        RECT 3.235 -159.965 3.565 -159.635 ;
        RECT 3.235 -161.325 3.565 -160.995 ;
        RECT 3.235 -162.685 3.565 -162.355 ;
        RECT 3.235 -164.045 3.565 -163.715 ;
        RECT 3.235 -165.405 3.565 -165.075 ;
        RECT 3.235 -166.765 3.565 -166.435 ;
        RECT 3.235 -168.125 3.565 -167.795 ;
        RECT 3.235 -169.485 3.565 -169.155 ;
        RECT 3.235 -170.845 3.565 -170.515 ;
        RECT 3.235 -172.205 3.565 -171.875 ;
        RECT 3.235 -173.565 3.565 -173.235 ;
        RECT 3.235 -174.925 3.565 -174.595 ;
        RECT 3.235 -176.285 3.565 -175.955 ;
        RECT 3.235 -177.645 3.565 -177.315 ;
        RECT 3.235 -183.29 3.565 -182.16 ;
        RECT 3.24 -183.405 3.56 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.595 244.04 4.925 245.17 ;
        RECT 4.595 239.875 4.925 240.205 ;
        RECT 4.595 238.515 4.925 238.845 ;
        RECT 4.595 237.155 4.925 237.485 ;
        RECT 4.6 237.155 4.92 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.595 -0.845 4.925 -0.515 ;
        RECT 4.595 -2.205 4.925 -1.875 ;
        RECT 4.595 -3.565 4.925 -3.235 ;
        RECT 4.6 -3.565 4.92 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.955 244.04 6.285 245.17 ;
        RECT 5.955 239.875 6.285 240.205 ;
        RECT 5.955 238.515 6.285 238.845 ;
        RECT 5.955 237.155 6.285 237.485 ;
        RECT 5.96 237.155 6.28 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.955 -0.845 6.285 -0.515 ;
        RECT 5.955 -2.205 6.285 -1.875 ;
        RECT 5.955 -3.565 6.285 -3.235 ;
        RECT 5.96 -3.565 6.28 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.315 244.04 7.645 245.17 ;
        RECT 7.315 239.875 7.645 240.205 ;
        RECT 7.315 238.515 7.645 238.845 ;
        RECT 7.315 237.155 7.645 237.485 ;
        RECT 7.32 237.155 7.64 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.315 -0.845 7.645 -0.515 ;
        RECT 7.315 -2.205 7.645 -1.875 ;
        RECT 7.315 -3.565 7.645 -3.235 ;
        RECT 7.32 -3.565 7.64 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.315 -91.965 7.645 -91.635 ;
        RECT 7.315 -93.325 7.645 -92.995 ;
        RECT 7.315 -94.685 7.645 -94.355 ;
        RECT 7.315 -96.045 7.645 -95.715 ;
        RECT 7.315 -97.405 7.645 -97.075 ;
        RECT 7.315 -98.765 7.645 -98.435 ;
        RECT 7.315 -100.125 7.645 -99.795 ;
        RECT 7.315 -101.485 7.645 -101.155 ;
        RECT 7.315 -102.845 7.645 -102.515 ;
        RECT 7.315 -104.205 7.645 -103.875 ;
        RECT 7.315 -105.565 7.645 -105.235 ;
        RECT 7.315 -106.925 7.645 -106.595 ;
        RECT 7.315 -108.285 7.645 -107.955 ;
        RECT 7.315 -109.645 7.645 -109.315 ;
        RECT 7.315 -111.005 7.645 -110.675 ;
        RECT 7.315 -112.365 7.645 -112.035 ;
        RECT 7.315 -113.725 7.645 -113.395 ;
        RECT 7.315 -115.085 7.645 -114.755 ;
        RECT 7.315 -116.445 7.645 -116.115 ;
        RECT 7.315 -117.805 7.645 -117.475 ;
        RECT 7.315 -119.165 7.645 -118.835 ;
        RECT 7.315 -120.525 7.645 -120.195 ;
        RECT 7.315 -121.885 7.645 -121.555 ;
        RECT 7.315 -123.245 7.645 -122.915 ;
        RECT 7.315 -124.605 7.645 -124.275 ;
        RECT 7.315 -125.965 7.645 -125.635 ;
        RECT 7.315 -127.325 7.645 -126.995 ;
        RECT 7.315 -128.685 7.645 -128.355 ;
        RECT 7.315 -130.045 7.645 -129.715 ;
        RECT 7.315 -131.405 7.645 -131.075 ;
        RECT 7.315 -132.765 7.645 -132.435 ;
        RECT 7.315 -134.125 7.645 -133.795 ;
        RECT 7.315 -135.485 7.645 -135.155 ;
        RECT 7.315 -136.845 7.645 -136.515 ;
        RECT 7.315 -138.205 7.645 -137.875 ;
        RECT 7.315 -139.565 7.645 -139.235 ;
        RECT 7.315 -140.925 7.645 -140.595 ;
        RECT 7.315 -142.285 7.645 -141.955 ;
        RECT 7.315 -143.645 7.645 -143.315 ;
        RECT 7.315 -145.005 7.645 -144.675 ;
        RECT 7.315 -146.365 7.645 -146.035 ;
        RECT 7.315 -147.725 7.645 -147.395 ;
        RECT 7.315 -149.085 7.645 -148.755 ;
        RECT 7.315 -150.445 7.645 -150.115 ;
        RECT 7.315 -151.805 7.645 -151.475 ;
        RECT 7.315 -153.165 7.645 -152.835 ;
        RECT 7.315 -154.525 7.645 -154.195 ;
        RECT 7.315 -155.885 7.645 -155.555 ;
        RECT 7.315 -157.245 7.645 -156.915 ;
        RECT 7.315 -158.605 7.645 -158.275 ;
        RECT 7.315 -159.965 7.645 -159.635 ;
        RECT 7.315 -161.325 7.645 -160.995 ;
        RECT 7.315 -162.685 7.645 -162.355 ;
        RECT 7.315 -164.045 7.645 -163.715 ;
        RECT 7.315 -165.405 7.645 -165.075 ;
        RECT 7.315 -166.765 7.645 -166.435 ;
        RECT 7.315 -168.125 7.645 -167.795 ;
        RECT 7.315 -169.485 7.645 -169.155 ;
        RECT 7.315 -170.845 7.645 -170.515 ;
        RECT 7.315 -172.205 7.645 -171.875 ;
        RECT 7.315 -173.565 7.645 -173.235 ;
        RECT 7.315 -174.925 7.645 -174.595 ;
        RECT 7.315 -176.285 7.645 -175.955 ;
        RECT 7.315 -177.645 7.645 -177.315 ;
        RECT 7.315 -183.29 7.645 -182.16 ;
        RECT 7.32 -183.405 7.64 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.675 244.04 9.005 245.17 ;
        RECT 8.675 239.875 9.005 240.205 ;
        RECT 8.675 238.515 9.005 238.845 ;
        RECT 8.675 237.155 9.005 237.485 ;
        RECT 8.68 237.155 9 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.675 -119.165 9.005 -118.835 ;
        RECT 8.675 -120.525 9.005 -120.195 ;
        RECT 8.675 -121.885 9.005 -121.555 ;
        RECT 8.675 -123.245 9.005 -122.915 ;
        RECT 8.675 -124.605 9.005 -124.275 ;
        RECT 8.675 -125.965 9.005 -125.635 ;
        RECT 8.675 -127.325 9.005 -126.995 ;
        RECT 8.675 -128.685 9.005 -128.355 ;
        RECT 8.675 -130.045 9.005 -129.715 ;
        RECT 8.675 -131.405 9.005 -131.075 ;
        RECT 8.675 -132.765 9.005 -132.435 ;
        RECT 8.675 -134.125 9.005 -133.795 ;
        RECT 8.675 -135.485 9.005 -135.155 ;
        RECT 8.675 -136.845 9.005 -136.515 ;
        RECT 8.675 -138.205 9.005 -137.875 ;
        RECT 8.675 -139.565 9.005 -139.235 ;
        RECT 8.675 -140.925 9.005 -140.595 ;
        RECT 8.675 -142.285 9.005 -141.955 ;
        RECT 8.675 -143.645 9.005 -143.315 ;
        RECT 8.675 -145.005 9.005 -144.675 ;
        RECT 8.675 -146.365 9.005 -146.035 ;
        RECT 8.675 -147.725 9.005 -147.395 ;
        RECT 8.675 -149.085 9.005 -148.755 ;
        RECT 8.675 -150.445 9.005 -150.115 ;
        RECT 8.675 -151.805 9.005 -151.475 ;
        RECT 8.675 -153.165 9.005 -152.835 ;
        RECT 8.675 -154.525 9.005 -154.195 ;
        RECT 8.675 -155.885 9.005 -155.555 ;
        RECT 8.675 -157.245 9.005 -156.915 ;
        RECT 8.675 -158.605 9.005 -158.275 ;
        RECT 8.675 -159.965 9.005 -159.635 ;
        RECT 8.675 -161.325 9.005 -160.995 ;
        RECT 8.675 -162.685 9.005 -162.355 ;
        RECT 8.675 -164.045 9.005 -163.715 ;
        RECT 8.675 -165.405 9.005 -165.075 ;
        RECT 8.675 -166.765 9.005 -166.435 ;
        RECT 8.675 -168.125 9.005 -167.795 ;
        RECT 8.675 -169.485 9.005 -169.155 ;
        RECT 8.675 -170.845 9.005 -170.515 ;
        RECT 8.675 -172.205 9.005 -171.875 ;
        RECT 8.675 -173.565 9.005 -173.235 ;
        RECT 8.675 -174.925 9.005 -174.595 ;
        RECT 8.675 -176.285 9.005 -175.955 ;
        RECT 8.675 -177.645 9.005 -177.315 ;
        RECT 8.675 -183.29 9.005 -182.16 ;
        RECT 8.68 -183.405 9 -95.04 ;
        RECT 8.675 -96.045 9.005 -95.715 ;
        RECT 8.675 -97.405 9.005 -97.075 ;
        RECT 8.675 -98.765 9.005 -98.435 ;
        RECT 8.675 -100.125 9.005 -99.795 ;
        RECT 8.675 -101.485 9.005 -101.155 ;
        RECT 8.675 -102.845 9.005 -102.515 ;
        RECT 8.675 -104.205 9.005 -103.875 ;
        RECT 8.675 -105.565 9.005 -105.235 ;
        RECT 8.675 -106.925 9.005 -106.595 ;
        RECT 8.675 -108.285 9.005 -107.955 ;
        RECT 8.675 -109.645 9.005 -109.315 ;
        RECT 8.675 -111.005 9.005 -110.675 ;
        RECT 8.675 -112.365 9.005 -112.035 ;
        RECT 8.675 -113.725 9.005 -113.395 ;
        RECT 8.675 -115.085 9.005 -114.755 ;
        RECT 8.675 -116.445 9.005 -116.115 ;
        RECT 8.675 -117.805 9.005 -117.475 ;
    END
    PORT
      LAYER met3 ;
        RECT -10.365 -174.925 -10.035 -174.595 ;
        RECT -10.365 -177.645 -10.035 -177.315 ;
        RECT -10.365 -183.29 -10.035 -182.16 ;
        RECT -10.36 -183.405 -10.04 -173.24 ;
    END
    PORT
      LAYER met3 ;
        RECT -9.005 244.04 -8.675 245.17 ;
        RECT -9.005 239.875 -8.675 240.205 ;
        RECT -9.005 238.515 -8.675 238.845 ;
        RECT -9.005 237.155 -8.675 237.485 ;
        RECT -9.005 235.795 -8.675 236.125 ;
        RECT -9.005 234.435 -8.675 234.765 ;
        RECT -9.005 233.075 -8.675 233.405 ;
        RECT -9.005 231.715 -8.675 232.045 ;
        RECT -9.005 227.635 -8.675 227.965 ;
        RECT -9.005 224.915 -8.675 225.245 ;
        RECT -9.005 218.115 -8.675 218.445 ;
        RECT -9.005 216.755 -8.675 217.085 ;
        RECT -9.005 207.235 -8.675 207.565 ;
        RECT -9.005 204.515 -8.675 204.845 ;
        RECT -9.005 203.155 -8.675 203.485 ;
        RECT -9.005 199.075 -8.675 199.405 ;
        RECT -9.005 196.355 -8.675 196.685 ;
        RECT -9.005 189.555 -8.675 189.885 ;
        RECT -9.005 188.195 -8.675 188.525 ;
        RECT -9.005 185.475 -8.675 185.805 ;
        RECT -9.005 178.675 -8.675 179.005 ;
        RECT -9.005 175.955 -8.675 176.285 ;
        RECT -9.005 174.595 -8.675 174.925 ;
        RECT -9.005 167.795 -8.675 168.125 ;
        RECT -9.005 160.995 -8.675 161.325 ;
        RECT -9.005 159.635 -8.675 159.965 ;
        RECT -9.005 156.915 -8.675 157.245 ;
        RECT -9.005 150.115 -8.675 150.445 ;
        RECT -9.005 147.395 -8.675 147.725 ;
        RECT -9.005 146.035 -8.675 146.365 ;
        RECT -9.005 139.235 -8.675 139.565 ;
        RECT -9.005 136.515 -8.675 136.845 ;
        RECT -9.005 132.435 -8.675 132.765 ;
        RECT -9.005 131.075 -8.675 131.405 ;
        RECT -9.005 128.355 -8.675 128.685 ;
        RECT -9.005 118.835 -8.675 119.165 ;
        RECT -9.005 117.475 -8.675 117.805 ;
        RECT -9.005 110.675 -8.675 111.005 ;
        RECT -9.005 107.955 -8.675 108.285 ;
        RECT -9.005 103.875 -8.675 104.205 ;
        RECT -9.005 99.795 -8.675 100.125 ;
        RECT -9.005 97.075 -8.675 97.405 ;
        RECT -9.005 90.275 -8.675 90.605 ;
        RECT -9.005 88.915 -8.675 89.245 ;
        RECT -9.005 82.115 -8.675 82.445 ;
        RECT -9.005 79.395 -8.675 79.725 ;
        RECT -9.005 75.315 -8.675 75.645 ;
        RECT -9.005 71.235 -8.675 71.565 ;
        RECT -9.005 68.515 -8.675 68.845 ;
        RECT -9.005 61.715 -8.675 62.045 ;
        RECT -9.005 60.355 -8.675 60.685 ;
        RECT -9.005 50.835 -8.675 51.165 ;
        RECT -9.005 46.755 -8.675 47.085 ;
        RECT -9.005 42.675 -8.675 43.005 ;
        RECT -9.005 39.955 -8.675 40.285 ;
        RECT -9.005 33.155 -8.675 33.485 ;
        RECT -9.005 31.795 -8.675 32.125 ;
        RECT -9.005 29.075 -8.675 29.405 ;
        RECT -9.005 22.275 -8.675 22.605 ;
        RECT -9.005 19.555 -8.675 19.885 ;
        RECT -9.005 18.195 -8.675 18.525 ;
        RECT -9.005 11.395 -8.675 11.725 ;
        RECT -9.005 4.595 -8.675 4.925 ;
        RECT -9.005 3.235 -8.675 3.565 ;
        RECT -9.005 1.875 -8.675 2.205 ;
        RECT -9.005 0.515 -8.675 0.845 ;
        RECT -9.005 -0.845 -8.675 -0.515 ;
        RECT -9.005 -2.205 -8.675 -1.875 ;
        RECT -9.005 -3.565 -8.675 -3.235 ;
        RECT -9.005 -4.925 -8.675 -4.595 ;
        RECT -9.005 -6.285 -8.675 -5.955 ;
        RECT -9.005 -7.645 -8.675 -7.315 ;
        RECT -9.005 -9.005 -8.675 -8.675 ;
        RECT -9.005 -10.365 -8.675 -10.035 ;
        RECT -9.005 -11.725 -8.675 -11.395 ;
        RECT -9.005 -13.085 -8.675 -12.755 ;
        RECT -9.005 -14.445 -8.675 -14.115 ;
        RECT -9.005 -15.805 -8.675 -15.475 ;
        RECT -9.005 -17.165 -8.675 -16.835 ;
        RECT -9 -19.2 -8.68 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -9.005 -109.645 -8.675 -109.315 ;
        RECT -9.005 -111.005 -8.675 -110.675 ;
        RECT -9.005 -112.365 -8.675 -112.035 ;
        RECT -9.005 -113.725 -8.675 -113.395 ;
        RECT -9.005 -115.085 -8.675 -114.755 ;
        RECT -9.005 -116.445 -8.675 -116.115 ;
        RECT -9.005 -117.805 -8.675 -117.475 ;
        RECT -9.005 -119.165 -8.675 -118.835 ;
        RECT -9.005 -121.885 -8.675 -121.555 ;
        RECT -9.005 -123.245 -8.675 -122.915 ;
        RECT -9.005 -124.605 -8.675 -124.275 ;
        RECT -9.005 -125.965 -8.675 -125.635 ;
        RECT -9.005 -127.325 -8.675 -126.995 ;
        RECT -9.005 -128.685 -8.675 -128.355 ;
        RECT -9.005 -130.045 -8.675 -129.715 ;
        RECT -9.005 -131.405 -8.675 -131.075 ;
        RECT -9.005 -132.765 -8.675 -132.435 ;
        RECT -9.005 -134.125 -8.675 -133.795 ;
        RECT -9.005 -135.485 -8.675 -135.155 ;
        RECT -9.005 -136.845 -8.675 -136.515 ;
        RECT -9.005 -138.205 -8.675 -137.875 ;
        RECT -9.005 -139.565 -8.675 -139.235 ;
        RECT -9.005 -140.925 -8.675 -140.595 ;
        RECT -9.005 -142.285 -8.675 -141.955 ;
        RECT -9.005 -143.645 -8.675 -143.315 ;
        RECT -9.005 -145.005 -8.675 -144.675 ;
        RECT -9.005 -146.365 -8.675 -146.035 ;
        RECT -9.005 -147.725 -8.675 -147.395 ;
        RECT -9.005 -149.085 -8.675 -148.755 ;
        RECT -9.005 -150.445 -8.675 -150.115 ;
        RECT -9.005 -151.805 -8.675 -151.475 ;
        RECT -9.005 -153.165 -8.675 -152.835 ;
        RECT -9.005 -154.525 -8.675 -154.195 ;
        RECT -9.005 -155.885 -8.675 -155.555 ;
        RECT -9.005 -157.245 -8.675 -156.915 ;
        RECT -9.005 -158.605 -8.675 -158.275 ;
        RECT -9.005 -159.965 -8.675 -159.635 ;
        RECT -9.005 -161.325 -8.675 -160.995 ;
        RECT -9.005 -162.685 -8.675 -162.355 ;
        RECT -9.005 -164.045 -8.675 -163.715 ;
        RECT -9.005 -165.405 -8.675 -165.075 ;
        RECT -9.005 -166.765 -8.675 -166.435 ;
        RECT -9.005 -168.125 -8.675 -167.795 ;
        RECT -9.005 -169.485 -8.675 -169.155 ;
        RECT -9.005 -170.845 -8.675 -170.515 ;
        RECT -9.005 -172.205 -8.675 -171.875 ;
        RECT -9.005 -173.565 -8.675 -173.235 ;
        RECT -9.005 -174.925 -8.675 -174.595 ;
        RECT -9.005 -176.285 -8.675 -175.955 ;
        RECT -9.005 -177.645 -8.675 -177.315 ;
        RECT -9.005 -183.29 -8.675 -182.16 ;
        RECT -9 -183.405 -8.68 -109.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -7.645 244.04 -7.315 245.17 ;
        RECT -7.645 239.875 -7.315 240.205 ;
        RECT -7.645 238.515 -7.315 238.845 ;
        RECT -7.645 237.155 -7.315 237.485 ;
        RECT -7.645 235.795 -7.315 236.125 ;
        RECT -7.645 234.435 -7.315 234.765 ;
        RECT -7.645 233.075 -7.315 233.405 ;
        RECT -7.645 231.715 -7.315 232.045 ;
        RECT -7.645 227.635 -7.315 227.965 ;
        RECT -7.645 224.915 -7.315 225.245 ;
        RECT -7.645 218.115 -7.315 218.445 ;
        RECT -7.645 216.755 -7.315 217.085 ;
        RECT -7.645 207.235 -7.315 207.565 ;
        RECT -7.645 204.515 -7.315 204.845 ;
        RECT -7.645 203.155 -7.315 203.485 ;
        RECT -7.645 199.075 -7.315 199.405 ;
        RECT -7.645 196.355 -7.315 196.685 ;
        RECT -7.645 189.555 -7.315 189.885 ;
        RECT -7.645 188.195 -7.315 188.525 ;
        RECT -7.645 185.475 -7.315 185.805 ;
        RECT -7.645 178.675 -7.315 179.005 ;
        RECT -7.645 175.955 -7.315 176.285 ;
        RECT -7.645 174.595 -7.315 174.925 ;
        RECT -7.645 167.795 -7.315 168.125 ;
        RECT -7.645 160.995 -7.315 161.325 ;
        RECT -7.645 159.635 -7.315 159.965 ;
        RECT -7.645 156.915 -7.315 157.245 ;
        RECT -7.645 150.115 -7.315 150.445 ;
        RECT -7.645 147.395 -7.315 147.725 ;
        RECT -7.645 146.035 -7.315 146.365 ;
        RECT -7.645 139.235 -7.315 139.565 ;
        RECT -7.645 136.515 -7.315 136.845 ;
        RECT -7.645 132.435 -7.315 132.765 ;
        RECT -7.645 131.075 -7.315 131.405 ;
        RECT -7.645 128.355 -7.315 128.685 ;
        RECT -7.645 118.835 -7.315 119.165 ;
        RECT -7.645 117.475 -7.315 117.805 ;
        RECT -7.645 110.675 -7.315 111.005 ;
        RECT -7.645 107.955 -7.315 108.285 ;
        RECT -7.645 103.875 -7.315 104.205 ;
        RECT -7.645 99.795 -7.315 100.125 ;
        RECT -7.645 97.075 -7.315 97.405 ;
        RECT -7.645 90.275 -7.315 90.605 ;
        RECT -7.645 88.915 -7.315 89.245 ;
        RECT -7.645 82.115 -7.315 82.445 ;
        RECT -7.645 79.395 -7.315 79.725 ;
        RECT -7.645 75.315 -7.315 75.645 ;
        RECT -7.645 71.235 -7.315 71.565 ;
        RECT -7.645 68.515 -7.315 68.845 ;
        RECT -7.645 61.715 -7.315 62.045 ;
        RECT -7.645 60.355 -7.315 60.685 ;
        RECT -7.645 50.835 -7.315 51.165 ;
        RECT -7.645 46.755 -7.315 47.085 ;
        RECT -7.645 42.675 -7.315 43.005 ;
        RECT -7.645 39.955 -7.315 40.285 ;
        RECT -7.645 33.155 -7.315 33.485 ;
        RECT -7.645 31.795 -7.315 32.125 ;
        RECT -7.645 29.075 -7.315 29.405 ;
        RECT -7.645 22.275 -7.315 22.605 ;
        RECT -7.645 19.555 -7.315 19.885 ;
        RECT -7.645 18.195 -7.315 18.525 ;
        RECT -7.645 11.395 -7.315 11.725 ;
        RECT -7.645 4.595 -7.315 4.925 ;
        RECT -7.645 3.235 -7.315 3.565 ;
        RECT -7.645 1.875 -7.315 2.205 ;
        RECT -7.645 0.515 -7.315 0.845 ;
        RECT -7.645 -0.845 -7.315 -0.515 ;
        RECT -7.645 -2.205 -7.315 -1.875 ;
        RECT -7.645 -3.565 -7.315 -3.235 ;
        RECT -7.645 -4.925 -7.315 -4.595 ;
        RECT -7.645 -6.285 -7.315 -5.955 ;
        RECT -7.645 -7.645 -7.315 -7.315 ;
        RECT -7.645 -9.005 -7.315 -8.675 ;
        RECT -7.645 -10.365 -7.315 -10.035 ;
        RECT -7.645 -11.725 -7.315 -11.395 ;
        RECT -7.645 -13.085 -7.315 -12.755 ;
        RECT -7.645 -14.445 -7.315 -14.115 ;
        RECT -7.645 -15.805 -7.315 -15.475 ;
        RECT -7.645 -17.165 -7.315 -16.835 ;
        RECT -7.645 -21.245 -7.315 -20.915 ;
        RECT -7.645 -22.605 -7.315 -22.275 ;
        RECT -7.645 -23.965 -7.315 -23.635 ;
        RECT -7.645 -25.325 -7.315 -24.995 ;
        RECT -7.645 -26.685 -7.315 -26.355 ;
        RECT -7.645 -28.045 -7.315 -27.715 ;
        RECT -7.645 -29.405 -7.315 -29.075 ;
        RECT -7.645 -30.765 -7.315 -30.435 ;
        RECT -7.645 -32.125 -7.315 -31.795 ;
        RECT -7.645 -33.485 -7.315 -33.155 ;
        RECT -7.645 -36.205 -7.315 -35.875 ;
        RECT -7.645 -37.565 -7.315 -37.235 ;
        RECT -7.645 -38.925 -7.315 -38.595 ;
        RECT -7.645 -40.285 -7.315 -39.955 ;
        RECT -7.645 -41.645 -7.315 -41.315 ;
        RECT -7.645 -43.005 -7.315 -42.675 ;
        RECT -7.645 -44.365 -7.315 -44.035 ;
        RECT -7.645 -45.725 -7.315 -45.395 ;
        RECT -7.645 -47.085 -7.315 -46.755 ;
        RECT -7.645 -48.445 -7.315 -48.115 ;
        RECT -7.645 -51.165 -7.315 -50.835 ;
        RECT -7.645 -52.525 -7.315 -52.195 ;
        RECT -7.645 -53.885 -7.315 -53.555 ;
        RECT -7.645 -55.245 -7.315 -54.915 ;
        RECT -7.645 -56.605 -7.315 -56.275 ;
        RECT -7.645 -57.965 -7.315 -57.635 ;
        RECT -7.645 -59.325 -7.315 -58.995 ;
        RECT -7.645 -60.685 -7.315 -60.355 ;
        RECT -7.645 -62.045 -7.315 -61.715 ;
        RECT -7.645 -63.405 -7.315 -63.075 ;
        RECT -7.645 -64.765 -7.315 -64.435 ;
        RECT -7.645 -66.125 -7.315 -65.795 ;
        RECT -7.645 -67.485 -7.315 -67.155 ;
        RECT -7.645 -68.845 -7.315 -68.515 ;
        RECT -7.645 -70.205 -7.315 -69.875 ;
        RECT -7.645 -71.565 -7.315 -71.235 ;
        RECT -7.645 -72.925 -7.315 -72.595 ;
        RECT -7.645 -74.285 -7.315 -73.955 ;
        RECT -7.645 -75.645 -7.315 -75.315 ;
        RECT -7.645 -77.005 -7.315 -76.675 ;
        RECT -7.645 -78.365 -7.315 -78.035 ;
        RECT -7.645 -79.725 -7.315 -79.395 ;
        RECT -7.645 -81.085 -7.315 -80.755 ;
        RECT -7.645 -82.445 -7.315 -82.115 ;
        RECT -7.645 -83.805 -7.315 -83.475 ;
        RECT -7.645 -85.165 -7.315 -84.835 ;
        RECT -7.645 -87.885 -7.315 -87.555 ;
        RECT -7.645 -89.245 -7.315 -88.915 ;
        RECT -7.645 -90.605 -7.315 -90.275 ;
        RECT -7.645 -91.965 -7.315 -91.635 ;
        RECT -7.645 -93.325 -7.315 -92.995 ;
        RECT -7.645 -94.685 -7.315 -94.355 ;
        RECT -7.645 -96.045 -7.315 -95.715 ;
        RECT -7.645 -97.405 -7.315 -97.075 ;
        RECT -7.645 -98.765 -7.315 -98.435 ;
        RECT -7.645 -100.125 -7.315 -99.795 ;
        RECT -7.645 -101.485 -7.315 -101.155 ;
        RECT -7.645 -102.845 -7.315 -102.515 ;
        RECT -7.645 -104.205 -7.315 -103.875 ;
        RECT -7.645 -105.565 -7.315 -105.235 ;
        RECT -7.645 -106.925 -7.315 -106.595 ;
        RECT -7.645 -108.285 -7.315 -107.955 ;
        RECT -7.645 -109.645 -7.315 -109.315 ;
        RECT -7.645 -111.005 -7.315 -110.675 ;
        RECT -7.645 -112.365 -7.315 -112.035 ;
        RECT -7.645 -113.725 -7.315 -113.395 ;
        RECT -7.645 -115.085 -7.315 -114.755 ;
        RECT -7.645 -116.445 -7.315 -116.115 ;
        RECT -7.645 -117.805 -7.315 -117.475 ;
        RECT -7.645 -119.165 -7.315 -118.835 ;
        RECT -7.645 -120.525 -7.315 -120.195 ;
        RECT -7.645 -121.885 -7.315 -121.555 ;
        RECT -7.645 -123.245 -7.315 -122.915 ;
        RECT -7.645 -124.605 -7.315 -124.275 ;
        RECT -7.645 -125.965 -7.315 -125.635 ;
        RECT -7.645 -127.325 -7.315 -126.995 ;
        RECT -7.645 -128.685 -7.315 -128.355 ;
        RECT -7.645 -130.045 -7.315 -129.715 ;
        RECT -7.645 -131.405 -7.315 -131.075 ;
        RECT -7.645 -132.765 -7.315 -132.435 ;
        RECT -7.645 -134.125 -7.315 -133.795 ;
        RECT -7.645 -135.485 -7.315 -135.155 ;
        RECT -7.645 -136.845 -7.315 -136.515 ;
        RECT -7.645 -138.205 -7.315 -137.875 ;
        RECT -7.645 -139.565 -7.315 -139.235 ;
        RECT -7.645 -140.925 -7.315 -140.595 ;
        RECT -7.645 -142.285 -7.315 -141.955 ;
        RECT -7.645 -143.645 -7.315 -143.315 ;
        RECT -7.645 -145.005 -7.315 -144.675 ;
        RECT -7.645 -146.365 -7.315 -146.035 ;
        RECT -7.645 -147.725 -7.315 -147.395 ;
        RECT -7.645 -149.085 -7.315 -148.755 ;
        RECT -7.645 -150.445 -7.315 -150.115 ;
        RECT -7.645 -151.805 -7.315 -151.475 ;
        RECT -7.645 -153.165 -7.315 -152.835 ;
        RECT -7.645 -154.525 -7.315 -154.195 ;
        RECT -7.645 -155.885 -7.315 -155.555 ;
        RECT -7.645 -157.245 -7.315 -156.915 ;
        RECT -7.645 -158.605 -7.315 -158.275 ;
        RECT -7.645 -159.965 -7.315 -159.635 ;
        RECT -7.645 -161.325 -7.315 -160.995 ;
        RECT -7.645 -162.685 -7.315 -162.355 ;
        RECT -7.645 -164.045 -7.315 -163.715 ;
        RECT -7.645 -165.405 -7.315 -165.075 ;
        RECT -7.645 -166.765 -7.315 -166.435 ;
        RECT -7.645 -168.125 -7.315 -167.795 ;
        RECT -7.645 -169.485 -7.315 -169.155 ;
        RECT -7.645 -170.845 -7.315 -170.515 ;
        RECT -7.645 -172.205 -7.315 -171.875 ;
        RECT -7.645 -173.565 -7.315 -173.235 ;
        RECT -7.645 -174.925 -7.315 -174.595 ;
        RECT -7.645 -176.285 -7.315 -175.955 ;
        RECT -7.645 -177.645 -7.315 -177.315 ;
        RECT -7.645 -183.29 -7.315 -182.16 ;
        RECT -7.64 -183.405 -7.32 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -6.285 244.04 -5.955 245.17 ;
        RECT -6.285 239.875 -5.955 240.205 ;
        RECT -6.285 238.515 -5.955 238.845 ;
        RECT -6.285 237.155 -5.955 237.485 ;
        RECT -6.285 -0.845 -5.955 -0.515 ;
        RECT -6.285 -2.205 -5.955 -1.875 ;
        RECT -6.285 -3.565 -5.955 -3.235 ;
        RECT -6.285 -4.925 -5.955 -4.595 ;
        RECT -6.285 -6.285 -5.955 -5.955 ;
        RECT -6.285 -7.645 -5.955 -7.315 ;
        RECT -6.285 -9.005 -5.955 -8.675 ;
        RECT -6.285 -10.365 -5.955 -10.035 ;
        RECT -6.285 -11.725 -5.955 -11.395 ;
        RECT -6.285 -13.085 -5.955 -12.755 ;
        RECT -6.285 -14.445 -5.955 -14.115 ;
        RECT -6.285 -15.805 -5.955 -15.475 ;
        RECT -6.285 -17.165 -5.955 -16.835 ;
        RECT -6.285 -21.245 -5.955 -20.915 ;
        RECT -6.285 -22.605 -5.955 -22.275 ;
        RECT -6.285 -23.965 -5.955 -23.635 ;
        RECT -6.285 -25.325 -5.955 -24.995 ;
        RECT -6.285 -26.685 -5.955 -26.355 ;
        RECT -6.285 -28.045 -5.955 -27.715 ;
        RECT -6.285 -29.405 -5.955 -29.075 ;
        RECT -6.285 -30.765 -5.955 -30.435 ;
        RECT -6.285 -32.125 -5.955 -31.795 ;
        RECT -6.285 -33.485 -5.955 -33.155 ;
        RECT -6.285 -36.205 -5.955 -35.875 ;
        RECT -6.285 -37.565 -5.955 -37.235 ;
        RECT -6.285 -38.925 -5.955 -38.595 ;
        RECT -6.285 -40.285 -5.955 -39.955 ;
        RECT -6.285 -41.645 -5.955 -41.315 ;
        RECT -6.285 -43.005 -5.955 -42.675 ;
        RECT -6.285 -44.365 -5.955 -44.035 ;
        RECT -6.285 -45.725 -5.955 -45.395 ;
        RECT -6.285 -47.085 -5.955 -46.755 ;
        RECT -6.285 -48.445 -5.955 -48.115 ;
        RECT -6.285 -51.165 -5.955 -50.835 ;
        RECT -6.285 -52.525 -5.955 -52.195 ;
        RECT -6.285 -53.885 -5.955 -53.555 ;
        RECT -6.285 -55.245 -5.955 -54.915 ;
        RECT -6.285 -56.605 -5.955 -56.275 ;
        RECT -6.285 -57.965 -5.955 -57.635 ;
        RECT -6.285 -59.325 -5.955 -58.995 ;
        RECT -6.285 -60.685 -5.955 -60.355 ;
        RECT -6.285 -62.045 -5.955 -61.715 ;
        RECT -6.285 -63.405 -5.955 -63.075 ;
        RECT -6.285 -64.765 -5.955 -64.435 ;
        RECT -6.285 -66.125 -5.955 -65.795 ;
        RECT -6.285 -67.485 -5.955 -67.155 ;
        RECT -6.285 -68.845 -5.955 -68.515 ;
        RECT -6.285 -70.205 -5.955 -69.875 ;
        RECT -6.285 -71.565 -5.955 -71.235 ;
        RECT -6.285 -72.925 -5.955 -72.595 ;
        RECT -6.285 -74.285 -5.955 -73.955 ;
        RECT -6.285 -75.645 -5.955 -75.315 ;
        RECT -6.285 -77.005 -5.955 -76.675 ;
        RECT -6.285 -78.365 -5.955 -78.035 ;
        RECT -6.285 -79.725 -5.955 -79.395 ;
        RECT -6.285 -81.085 -5.955 -80.755 ;
        RECT -6.285 -82.445 -5.955 -82.115 ;
        RECT -6.285 -83.805 -5.955 -83.475 ;
        RECT -6.285 -85.165 -5.955 -84.835 ;
        RECT -6.285 -87.885 -5.955 -87.555 ;
        RECT -6.285 -89.245 -5.955 -88.915 ;
        RECT -6.285 -90.605 -5.955 -90.275 ;
        RECT -6.285 -91.965 -5.955 -91.635 ;
        RECT -6.285 -93.325 -5.955 -92.995 ;
        RECT -6.285 -94.685 -5.955 -94.355 ;
        RECT -6.285 -96.045 -5.955 -95.715 ;
        RECT -6.285 -97.405 -5.955 -97.075 ;
        RECT -6.285 -98.765 -5.955 -98.435 ;
        RECT -6.285 -100.125 -5.955 -99.795 ;
        RECT -6.285 -101.485 -5.955 -101.155 ;
        RECT -6.285 -102.845 -5.955 -102.515 ;
        RECT -6.285 -104.205 -5.955 -103.875 ;
        RECT -6.285 -105.565 -5.955 -105.235 ;
        RECT -6.285 -106.925 -5.955 -106.595 ;
        RECT -6.285 -108.285 -5.955 -107.955 ;
        RECT -6.285 -109.645 -5.955 -109.315 ;
        RECT -6.285 -111.005 -5.955 -110.675 ;
        RECT -6.285 -112.365 -5.955 -112.035 ;
        RECT -6.285 -113.725 -5.955 -113.395 ;
        RECT -6.285 -115.085 -5.955 -114.755 ;
        RECT -6.285 -116.445 -5.955 -116.115 ;
        RECT -6.285 -117.805 -5.955 -117.475 ;
        RECT -6.285 -119.165 -5.955 -118.835 ;
        RECT -6.285 -120.525 -5.955 -120.195 ;
        RECT -6.285 -121.885 -5.955 -121.555 ;
        RECT -6.285 -123.245 -5.955 -122.915 ;
        RECT -6.285 -124.605 -5.955 -124.275 ;
        RECT -6.285 -125.965 -5.955 -125.635 ;
        RECT -6.285 -127.325 -5.955 -126.995 ;
        RECT -6.285 -128.685 -5.955 -128.355 ;
        RECT -6.285 -130.045 -5.955 -129.715 ;
        RECT -6.285 -131.405 -5.955 -131.075 ;
        RECT -6.285 -132.765 -5.955 -132.435 ;
        RECT -6.285 -134.125 -5.955 -133.795 ;
        RECT -6.285 -135.485 -5.955 -135.155 ;
        RECT -6.285 -136.845 -5.955 -136.515 ;
        RECT -6.285 -138.205 -5.955 -137.875 ;
        RECT -6.285 -139.565 -5.955 -139.235 ;
        RECT -6.285 -140.925 -5.955 -140.595 ;
        RECT -6.285 -142.285 -5.955 -141.955 ;
        RECT -6.285 -143.645 -5.955 -143.315 ;
        RECT -6.285 -145.005 -5.955 -144.675 ;
        RECT -6.285 -146.365 -5.955 -146.035 ;
        RECT -6.285 -147.725 -5.955 -147.395 ;
        RECT -6.285 -149.085 -5.955 -148.755 ;
        RECT -6.285 -150.445 -5.955 -150.115 ;
        RECT -6.285 -151.805 -5.955 -151.475 ;
        RECT -6.285 -153.165 -5.955 -152.835 ;
        RECT -6.285 -154.525 -5.955 -154.195 ;
        RECT -6.285 -155.885 -5.955 -155.555 ;
        RECT -6.285 -157.245 -5.955 -156.915 ;
        RECT -6.285 -158.605 -5.955 -158.275 ;
        RECT -6.285 -159.965 -5.955 -159.635 ;
        RECT -6.285 -161.325 -5.955 -160.995 ;
        RECT -6.285 -162.685 -5.955 -162.355 ;
        RECT -6.285 -164.045 -5.955 -163.715 ;
        RECT -6.285 -165.405 -5.955 -165.075 ;
        RECT -6.285 -166.765 -5.955 -166.435 ;
        RECT -6.285 -168.125 -5.955 -167.795 ;
        RECT -6.285 -169.485 -5.955 -169.155 ;
        RECT -6.285 -170.845 -5.955 -170.515 ;
        RECT -6.285 -172.205 -5.955 -171.875 ;
        RECT -6.285 -173.565 -5.955 -173.235 ;
        RECT -6.285 -174.925 -5.955 -174.595 ;
        RECT -6.285 -176.285 -5.955 -175.955 ;
        RECT -6.285 -177.645 -5.955 -177.315 ;
        RECT -6.285 -183.29 -5.955 -182.16 ;
        RECT -6.28 -183.405 -5.96 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -4.925 244.04 -4.595 245.17 ;
        RECT -4.925 239.875 -4.595 240.205 ;
        RECT -4.925 238.515 -4.595 238.845 ;
        RECT -4.925 237.155 -4.595 237.485 ;
        RECT -4.925 235.17 -4.595 235.5 ;
        RECT -4.925 232.995 -4.595 233.325 ;
        RECT -4.925 231.415 -4.595 231.745 ;
        RECT -4.925 230.565 -4.595 230.895 ;
        RECT -4.925 228.255 -4.595 228.585 ;
        RECT -4.925 227.405 -4.595 227.735 ;
        RECT -4.925 225.095 -4.595 225.425 ;
        RECT -4.925 224.245 -4.595 224.575 ;
        RECT -4.925 221.935 -4.595 222.265 ;
        RECT -4.925 221.085 -4.595 221.415 ;
        RECT -4.925 218.775 -4.595 219.105 ;
        RECT -4.925 217.195 -4.595 217.525 ;
        RECT -4.925 216.345 -4.595 216.675 ;
        RECT -4.925 214.035 -4.595 214.365 ;
        RECT -4.925 213.185 -4.595 213.515 ;
        RECT -4.925 210.875 -4.595 211.205 ;
        RECT -4.925 210.025 -4.595 210.355 ;
        RECT -4.925 207.715 -4.595 208.045 ;
        RECT -4.925 206.865 -4.595 207.195 ;
        RECT -4.925 204.555 -4.595 204.885 ;
        RECT -4.925 202.975 -4.595 203.305 ;
        RECT -4.925 202.125 -4.595 202.455 ;
        RECT -4.925 199.815 -4.595 200.145 ;
        RECT -4.925 198.965 -4.595 199.295 ;
        RECT -4.925 196.655 -4.595 196.985 ;
        RECT -4.925 195.805 -4.595 196.135 ;
        RECT -4.925 193.495 -4.595 193.825 ;
        RECT -4.925 192.645 -4.595 192.975 ;
        RECT -4.925 190.335 -4.595 190.665 ;
        RECT -4.925 188.755 -4.595 189.085 ;
        RECT -4.925 187.905 -4.595 188.235 ;
        RECT -4.925 185.595 -4.595 185.925 ;
        RECT -4.925 184.745 -4.595 185.075 ;
        RECT -4.925 182.435 -4.595 182.765 ;
        RECT -4.925 181.585 -4.595 181.915 ;
        RECT -4.925 179.275 -4.595 179.605 ;
        RECT -4.925 178.425 -4.595 178.755 ;
        RECT -4.925 176.115 -4.595 176.445 ;
        RECT -4.925 174.535 -4.595 174.865 ;
        RECT -4.925 173.685 -4.595 174.015 ;
        RECT -4.925 171.375 -4.595 171.705 ;
        RECT -4.925 170.525 -4.595 170.855 ;
        RECT -4.925 168.215 -4.595 168.545 ;
        RECT -4.925 167.365 -4.595 167.695 ;
        RECT -4.925 165.055 -4.595 165.385 ;
        RECT -4.925 164.205 -4.595 164.535 ;
        RECT -4.925 161.895 -4.595 162.225 ;
        RECT -4.925 160.315 -4.595 160.645 ;
        RECT -4.925 159.465 -4.595 159.795 ;
        RECT -4.925 157.155 -4.595 157.485 ;
        RECT -4.925 156.305 -4.595 156.635 ;
        RECT -4.925 153.995 -4.595 154.325 ;
        RECT -4.925 153.145 -4.595 153.475 ;
        RECT -4.925 150.835 -4.595 151.165 ;
        RECT -4.925 149.985 -4.595 150.315 ;
        RECT -4.925 147.675 -4.595 148.005 ;
        RECT -4.925 146.095 -4.595 146.425 ;
        RECT -4.925 145.245 -4.595 145.575 ;
        RECT -4.925 142.935 -4.595 143.265 ;
        RECT -4.925 142.085 -4.595 142.415 ;
        RECT -4.925 139.775 -4.595 140.105 ;
        RECT -4.925 138.925 -4.595 139.255 ;
        RECT -4.925 136.615 -4.595 136.945 ;
        RECT -4.925 135.765 -4.595 136.095 ;
        RECT -4.925 133.455 -4.595 133.785 ;
        RECT -4.925 131.875 -4.595 132.205 ;
        RECT -4.925 131.025 -4.595 131.355 ;
        RECT -4.925 128.715 -4.595 129.045 ;
        RECT -4.925 127.865 -4.595 128.195 ;
        RECT -4.925 125.555 -4.595 125.885 ;
        RECT -4.925 124.705 -4.595 125.035 ;
        RECT -4.925 122.395 -4.595 122.725 ;
        RECT -4.925 121.545 -4.595 121.875 ;
        RECT -4.925 119.235 -4.595 119.565 ;
        RECT -4.925 117.655 -4.595 117.985 ;
        RECT -4.925 116.805 -4.595 117.135 ;
        RECT -4.925 114.495 -4.595 114.825 ;
        RECT -4.925 113.645 -4.595 113.975 ;
        RECT -4.925 111.335 -4.595 111.665 ;
        RECT -4.925 110.485 -4.595 110.815 ;
        RECT -4.925 108.175 -4.595 108.505 ;
        RECT -4.925 107.325 -4.595 107.655 ;
        RECT -4.925 105.015 -4.595 105.345 ;
        RECT -4.925 103.435 -4.595 103.765 ;
        RECT -4.925 102.585 -4.595 102.915 ;
        RECT -4.925 100.275 -4.595 100.605 ;
        RECT -4.925 99.425 -4.595 99.755 ;
        RECT -4.925 97.115 -4.595 97.445 ;
        RECT -4.925 96.265 -4.595 96.595 ;
        RECT -4.925 93.955 -4.595 94.285 ;
        RECT -4.925 93.105 -4.595 93.435 ;
        RECT -4.925 90.795 -4.595 91.125 ;
        RECT -4.925 89.215 -4.595 89.545 ;
        RECT -4.925 88.365 -4.595 88.695 ;
        RECT -4.925 86.055 -4.595 86.385 ;
        RECT -4.925 85.205 -4.595 85.535 ;
        RECT -4.925 82.895 -4.595 83.225 ;
        RECT -4.925 82.045 -4.595 82.375 ;
        RECT -4.925 79.735 -4.595 80.065 ;
        RECT -4.925 78.885 -4.595 79.215 ;
        RECT -4.925 76.575 -4.595 76.905 ;
        RECT -4.925 74.995 -4.595 75.325 ;
        RECT -4.925 74.145 -4.595 74.475 ;
        RECT -4.925 71.835 -4.595 72.165 ;
        RECT -4.925 70.985 -4.595 71.315 ;
        RECT -4.925 68.675 -4.595 69.005 ;
        RECT -4.925 67.825 -4.595 68.155 ;
        RECT -4.925 65.515 -4.595 65.845 ;
        RECT -4.925 64.665 -4.595 64.995 ;
        RECT -4.925 62.355 -4.595 62.685 ;
        RECT -4.925 60.775 -4.595 61.105 ;
        RECT -4.925 59.925 -4.595 60.255 ;
        RECT -4.925 57.615 -4.595 57.945 ;
        RECT -4.925 56.765 -4.595 57.095 ;
        RECT -4.925 54.455 -4.595 54.785 ;
        RECT -4.925 53.605 -4.595 53.935 ;
        RECT -4.925 51.295 -4.595 51.625 ;
        RECT -4.925 50.445 -4.595 50.775 ;
        RECT -4.925 48.135 -4.595 48.465 ;
        RECT -4.925 46.555 -4.595 46.885 ;
        RECT -4.925 45.705 -4.595 46.035 ;
        RECT -4.925 43.395 -4.595 43.725 ;
        RECT -4.925 42.545 -4.595 42.875 ;
        RECT -4.925 40.235 -4.595 40.565 ;
        RECT -4.925 39.385 -4.595 39.715 ;
        RECT -4.925 37.075 -4.595 37.405 ;
        RECT -4.925 36.225 -4.595 36.555 ;
        RECT -4.925 33.915 -4.595 34.245 ;
        RECT -4.925 32.335 -4.595 32.665 ;
        RECT -4.925 31.485 -4.595 31.815 ;
        RECT -4.925 29.175 -4.595 29.505 ;
        RECT -4.925 28.325 -4.595 28.655 ;
        RECT -4.925 26.015 -4.595 26.345 ;
        RECT -4.925 25.165 -4.595 25.495 ;
        RECT -4.925 22.855 -4.595 23.185 ;
        RECT -4.925 22.005 -4.595 22.335 ;
        RECT -4.925 19.695 -4.595 20.025 ;
        RECT -4.925 18.115 -4.595 18.445 ;
        RECT -4.925 17.265 -4.595 17.595 ;
        RECT -4.925 14.955 -4.595 15.285 ;
        RECT -4.925 14.105 -4.595 14.435 ;
        RECT -4.925 11.795 -4.595 12.125 ;
        RECT -4.925 10.945 -4.595 11.275 ;
        RECT -4.925 8.635 -4.595 8.965 ;
        RECT -4.925 7.785 -4.595 8.115 ;
        RECT -4.925 5.475 -4.595 5.805 ;
        RECT -4.925 3.895 -4.595 4.225 ;
        RECT -4.925 3.045 -4.595 3.375 ;
        RECT -4.925 0.87 -4.595 1.2 ;
        RECT -4.925 -0.845 -4.595 -0.515 ;
        RECT -4.925 -2.205 -4.595 -1.875 ;
        RECT -4.925 -3.565 -4.595 -3.235 ;
        RECT -4.925 -4.925 -4.595 -4.595 ;
        RECT -4.925 -6.285 -4.595 -5.955 ;
        RECT -4.925 -7.645 -4.595 -7.315 ;
        RECT -4.925 -9.005 -4.595 -8.675 ;
        RECT -4.925 -10.365 -4.595 -10.035 ;
        RECT -4.925 -11.725 -4.595 -11.395 ;
        RECT -4.925 -13.085 -4.595 -12.755 ;
        RECT -4.925 -14.445 -4.595 -14.115 ;
        RECT -4.925 -15.805 -4.595 -15.475 ;
        RECT -4.925 -17.165 -4.595 -16.835 ;
        RECT -4.925 -21.245 -4.595 -20.915 ;
        RECT -4.925 -22.605 -4.595 -22.275 ;
        RECT -4.925 -23.965 -4.595 -23.635 ;
        RECT -4.925 -25.325 -4.595 -24.995 ;
        RECT -4.925 -26.685 -4.595 -26.355 ;
        RECT -4.925 -28.045 -4.595 -27.715 ;
        RECT -4.925 -29.405 -4.595 -29.075 ;
        RECT -4.925 -30.765 -4.595 -30.435 ;
        RECT -4.925 -32.125 -4.595 -31.795 ;
        RECT -4.925 -33.485 -4.595 -33.155 ;
        RECT -4.925 -36.205 -4.595 -35.875 ;
        RECT -4.925 -37.565 -4.595 -37.235 ;
        RECT -4.925 -38.925 -4.595 -38.595 ;
        RECT -4.925 -40.285 -4.595 -39.955 ;
        RECT -4.925 -41.645 -4.595 -41.315 ;
        RECT -4.925 -43.005 -4.595 -42.675 ;
        RECT -4.925 -44.365 -4.595 -44.035 ;
        RECT -4.925 -45.725 -4.595 -45.395 ;
        RECT -4.925 -47.085 -4.595 -46.755 ;
        RECT -4.925 -48.445 -4.595 -48.115 ;
        RECT -4.925 -51.165 -4.595 -50.835 ;
        RECT -4.925 -52.525 -4.595 -52.195 ;
        RECT -4.925 -53.885 -4.595 -53.555 ;
        RECT -4.925 -55.245 -4.595 -54.915 ;
        RECT -4.925 -56.605 -4.595 -56.275 ;
        RECT -4.925 -57.965 -4.595 -57.635 ;
        RECT -4.925 -59.325 -4.595 -58.995 ;
        RECT -4.925 -60.685 -4.595 -60.355 ;
        RECT -4.925 -62.045 -4.595 -61.715 ;
        RECT -4.925 -63.405 -4.595 -63.075 ;
        RECT -4.925 -64.765 -4.595 -64.435 ;
        RECT -4.925 -66.125 -4.595 -65.795 ;
        RECT -4.925 -67.485 -4.595 -67.155 ;
        RECT -4.925 -68.845 -4.595 -68.515 ;
        RECT -4.925 -70.205 -4.595 -69.875 ;
        RECT -4.925 -71.565 -4.595 -71.235 ;
        RECT -4.925 -72.925 -4.595 -72.595 ;
        RECT -4.925 -74.285 -4.595 -73.955 ;
        RECT -4.925 -75.645 -4.595 -75.315 ;
        RECT -4.925 -77.005 -4.595 -76.675 ;
        RECT -4.925 -78.365 -4.595 -78.035 ;
        RECT -4.925 -79.725 -4.595 -79.395 ;
        RECT -4.925 -81.085 -4.595 -80.755 ;
        RECT -4.925 -82.445 -4.595 -82.115 ;
        RECT -4.925 -83.805 -4.595 -83.475 ;
        RECT -4.925 -85.165 -4.595 -84.835 ;
        RECT -4.925 -87.885 -4.595 -87.555 ;
        RECT -4.925 -89.245 -4.595 -88.915 ;
        RECT -4.925 -90.605 -4.595 -90.275 ;
        RECT -4.925 -91.965 -4.595 -91.635 ;
        RECT -4.925 -93.325 -4.595 -92.995 ;
        RECT -4.925 -94.685 -4.595 -94.355 ;
        RECT -4.925 -96.045 -4.595 -95.715 ;
        RECT -4.925 -97.405 -4.595 -97.075 ;
        RECT -4.925 -98.765 -4.595 -98.435 ;
        RECT -4.925 -100.125 -4.595 -99.795 ;
        RECT -4.925 -101.485 -4.595 -101.155 ;
        RECT -4.925 -102.845 -4.595 -102.515 ;
        RECT -4.925 -104.205 -4.595 -103.875 ;
        RECT -4.925 -105.565 -4.595 -105.235 ;
        RECT -4.925 -106.925 -4.595 -106.595 ;
        RECT -4.925 -108.285 -4.595 -107.955 ;
        RECT -4.925 -109.645 -4.595 -109.315 ;
        RECT -4.925 -111.005 -4.595 -110.675 ;
        RECT -4.925 -112.365 -4.595 -112.035 ;
        RECT -4.925 -113.725 -4.595 -113.395 ;
        RECT -4.925 -115.085 -4.595 -114.755 ;
        RECT -4.925 -116.445 -4.595 -116.115 ;
        RECT -4.925 -117.805 -4.595 -117.475 ;
        RECT -4.925 -119.165 -4.595 -118.835 ;
        RECT -4.925 -120.525 -4.595 -120.195 ;
        RECT -4.925 -121.885 -4.595 -121.555 ;
        RECT -4.925 -123.245 -4.595 -122.915 ;
        RECT -4.925 -124.605 -4.595 -124.275 ;
        RECT -4.925 -125.965 -4.595 -125.635 ;
        RECT -4.925 -127.325 -4.595 -126.995 ;
        RECT -4.925 -128.685 -4.595 -128.355 ;
        RECT -4.925 -130.045 -4.595 -129.715 ;
        RECT -4.925 -131.405 -4.595 -131.075 ;
        RECT -4.925 -132.765 -4.595 -132.435 ;
        RECT -4.925 -134.125 -4.595 -133.795 ;
        RECT -4.925 -135.485 -4.595 -135.155 ;
        RECT -4.925 -136.845 -4.595 -136.515 ;
        RECT -4.925 -138.205 -4.595 -137.875 ;
        RECT -4.925 -139.565 -4.595 -139.235 ;
        RECT -4.925 -140.925 -4.595 -140.595 ;
        RECT -4.925 -142.285 -4.595 -141.955 ;
        RECT -4.925 -143.645 -4.595 -143.315 ;
        RECT -4.925 -145.005 -4.595 -144.675 ;
        RECT -4.925 -146.365 -4.595 -146.035 ;
        RECT -4.925 -147.725 -4.595 -147.395 ;
        RECT -4.925 -149.085 -4.595 -148.755 ;
        RECT -4.925 -150.445 -4.595 -150.115 ;
        RECT -4.925 -151.805 -4.595 -151.475 ;
        RECT -4.925 -153.165 -4.595 -152.835 ;
        RECT -4.925 -154.525 -4.595 -154.195 ;
        RECT -4.925 -155.885 -4.595 -155.555 ;
        RECT -4.925 -157.245 -4.595 -156.915 ;
        RECT -4.925 -158.605 -4.595 -158.275 ;
        RECT -4.925 -159.965 -4.595 -159.635 ;
        RECT -4.925 -161.325 -4.595 -160.995 ;
        RECT -4.925 -162.685 -4.595 -162.355 ;
        RECT -4.925 -164.045 -4.595 -163.715 ;
        RECT -4.925 -165.405 -4.595 -165.075 ;
        RECT -4.925 -166.765 -4.595 -166.435 ;
        RECT -4.925 -168.125 -4.595 -167.795 ;
        RECT -4.925 -169.485 -4.595 -169.155 ;
        RECT -4.925 -170.845 -4.595 -170.515 ;
        RECT -4.925 -172.205 -4.595 -171.875 ;
        RECT -4.925 -173.565 -4.595 -173.235 ;
        RECT -4.925 -174.925 -4.595 -174.595 ;
        RECT -4.925 -176.285 -4.595 -175.955 ;
        RECT -4.925 -177.645 -4.595 -177.315 ;
        RECT -4.925 -183.29 -4.595 -182.16 ;
        RECT -4.92 -183.405 -4.6 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -3.565 121.545 -3.235 121.875 ;
        RECT -3.565 119.235 -3.235 119.565 ;
        RECT -3.565 117.655 -3.235 117.985 ;
        RECT -3.565 116.805 -3.235 117.135 ;
        RECT -3.565 114.495 -3.235 114.825 ;
        RECT -3.565 113.645 -3.235 113.975 ;
        RECT -3.565 111.335 -3.235 111.665 ;
        RECT -3.565 110.485 -3.235 110.815 ;
        RECT -3.565 108.175 -3.235 108.505 ;
        RECT -3.565 107.325 -3.235 107.655 ;
        RECT -3.565 105.015 -3.235 105.345 ;
        RECT -3.565 103.435 -3.235 103.765 ;
        RECT -3.565 102.585 -3.235 102.915 ;
        RECT -3.565 100.275 -3.235 100.605 ;
        RECT -3.565 99.425 -3.235 99.755 ;
        RECT -3.565 97.115 -3.235 97.445 ;
        RECT -3.565 96.265 -3.235 96.595 ;
        RECT -3.565 93.955 -3.235 94.285 ;
        RECT -3.565 93.105 -3.235 93.435 ;
        RECT -3.565 90.795 -3.235 91.125 ;
        RECT -3.565 89.215 -3.235 89.545 ;
        RECT -3.565 88.365 -3.235 88.695 ;
        RECT -3.565 86.055 -3.235 86.385 ;
        RECT -3.565 85.205 -3.235 85.535 ;
        RECT -3.565 82.895 -3.235 83.225 ;
        RECT -3.565 82.045 -3.235 82.375 ;
        RECT -3.565 79.735 -3.235 80.065 ;
        RECT -3.565 78.885 -3.235 79.215 ;
        RECT -3.565 76.575 -3.235 76.905 ;
        RECT -3.565 74.995 -3.235 75.325 ;
        RECT -3.565 74.145 -3.235 74.475 ;
        RECT -3.565 71.835 -3.235 72.165 ;
        RECT -3.565 70.985 -3.235 71.315 ;
        RECT -3.565 68.675 -3.235 69.005 ;
        RECT -3.565 67.825 -3.235 68.155 ;
        RECT -3.565 65.515 -3.235 65.845 ;
        RECT -3.565 64.665 -3.235 64.995 ;
        RECT -3.565 62.355 -3.235 62.685 ;
        RECT -3.565 60.775 -3.235 61.105 ;
        RECT -3.565 59.925 -3.235 60.255 ;
        RECT -3.565 57.615 -3.235 57.945 ;
        RECT -3.565 56.765 -3.235 57.095 ;
        RECT -3.565 54.455 -3.235 54.785 ;
        RECT -3.565 53.605 -3.235 53.935 ;
        RECT -3.565 51.295 -3.235 51.625 ;
        RECT -3.565 50.445 -3.235 50.775 ;
        RECT -3.565 48.135 -3.235 48.465 ;
        RECT -3.565 46.555 -3.235 46.885 ;
        RECT -3.565 45.705 -3.235 46.035 ;
        RECT -3.565 43.395 -3.235 43.725 ;
        RECT -3.565 42.545 -3.235 42.875 ;
        RECT -3.565 40.235 -3.235 40.565 ;
        RECT -3.565 39.385 -3.235 39.715 ;
        RECT -3.565 37.075 -3.235 37.405 ;
        RECT -3.565 36.225 -3.235 36.555 ;
        RECT -3.565 33.915 -3.235 34.245 ;
        RECT -3.565 32.335 -3.235 32.665 ;
        RECT -3.565 31.485 -3.235 31.815 ;
        RECT -3.565 29.175 -3.235 29.505 ;
        RECT -3.565 28.325 -3.235 28.655 ;
        RECT -3.565 26.015 -3.235 26.345 ;
        RECT -3.565 25.165 -3.235 25.495 ;
        RECT -3.565 22.855 -3.235 23.185 ;
        RECT -3.565 22.005 -3.235 22.335 ;
        RECT -3.565 19.695 -3.235 20.025 ;
        RECT -3.565 18.115 -3.235 18.445 ;
        RECT -3.565 17.265 -3.235 17.595 ;
        RECT -3.565 14.955 -3.235 15.285 ;
        RECT -3.565 14.105 -3.235 14.435 ;
        RECT -3.565 11.795 -3.235 12.125 ;
        RECT -3.565 10.945 -3.235 11.275 ;
        RECT -3.565 8.635 -3.235 8.965 ;
        RECT -3.565 7.785 -3.235 8.115 ;
        RECT -3.565 5.475 -3.235 5.805 ;
        RECT -3.565 3.895 -3.235 4.225 ;
        RECT -3.565 3.045 -3.235 3.375 ;
        RECT -3.565 0.87 -3.235 1.2 ;
        RECT -3.565 -0.845 -3.235 -0.515 ;
        RECT -3.565 -2.205 -3.235 -1.875 ;
        RECT -3.565 -3.565 -3.235 -3.235 ;
        RECT -3.565 -4.925 -3.235 -4.595 ;
        RECT -3.565 -6.285 -3.235 -5.955 ;
        RECT -3.565 -7.645 -3.235 -7.315 ;
        RECT -3.565 -9.005 -3.235 -8.675 ;
        RECT -3.565 -10.365 -3.235 -10.035 ;
        RECT -3.565 -11.725 -3.235 -11.395 ;
        RECT -3.565 -13.085 -3.235 -12.755 ;
        RECT -3.565 -14.445 -3.235 -14.115 ;
        RECT -3.565 -15.805 -3.235 -15.475 ;
        RECT -3.565 -17.165 -3.235 -16.835 ;
        RECT -3.565 -21.245 -3.235 -20.915 ;
        RECT -3.565 -22.605 -3.235 -22.275 ;
        RECT -3.565 -23.965 -3.235 -23.635 ;
        RECT -3.565 -25.325 -3.235 -24.995 ;
        RECT -3.565 -26.685 -3.235 -26.355 ;
        RECT -3.565 -28.045 -3.235 -27.715 ;
        RECT -3.565 -29.405 -3.235 -29.075 ;
        RECT -3.565 -30.765 -3.235 -30.435 ;
        RECT -3.565 -32.125 -3.235 -31.795 ;
        RECT -3.565 -33.485 -3.235 -33.155 ;
        RECT -3.565 -36.205 -3.235 -35.875 ;
        RECT -3.565 -37.565 -3.235 -37.235 ;
        RECT -3.565 -38.925 -3.235 -38.595 ;
        RECT -3.565 -40.285 -3.235 -39.955 ;
        RECT -3.565 -41.645 -3.235 -41.315 ;
        RECT -3.565 -43.005 -3.235 -42.675 ;
        RECT -3.565 -44.365 -3.235 -44.035 ;
        RECT -3.565 -45.725 -3.235 -45.395 ;
        RECT -3.565 -47.085 -3.235 -46.755 ;
        RECT -3.565 -48.445 -3.235 -48.115 ;
        RECT -3.565 -51.165 -3.235 -50.835 ;
        RECT -3.565 -52.525 -3.235 -52.195 ;
        RECT -3.565 -53.885 -3.235 -53.555 ;
        RECT -3.565 -55.245 -3.235 -54.915 ;
        RECT -3.565 -56.605 -3.235 -56.275 ;
        RECT -3.565 -57.965 -3.235 -57.635 ;
        RECT -3.565 -59.325 -3.235 -58.995 ;
        RECT -3.565 -60.685 -3.235 -60.355 ;
        RECT -3.565 -62.045 -3.235 -61.715 ;
        RECT -3.565 -63.405 -3.235 -63.075 ;
        RECT -3.565 -64.765 -3.235 -64.435 ;
        RECT -3.565 -66.125 -3.235 -65.795 ;
        RECT -3.565 -67.485 -3.235 -67.155 ;
        RECT -3.565 -68.845 -3.235 -68.515 ;
        RECT -3.565 -70.205 -3.235 -69.875 ;
        RECT -3.565 -71.565 -3.235 -71.235 ;
        RECT -3.565 -72.925 -3.235 -72.595 ;
        RECT -3.565 -74.285 -3.235 -73.955 ;
        RECT -3.565 -75.645 -3.235 -75.315 ;
        RECT -3.565 -77.005 -3.235 -76.675 ;
        RECT -3.565 -78.365 -3.235 -78.035 ;
        RECT -3.565 -79.725 -3.235 -79.395 ;
        RECT -3.565 -81.085 -3.235 -80.755 ;
        RECT -3.565 -82.445 -3.235 -82.115 ;
        RECT -3.565 -83.805 -3.235 -83.475 ;
        RECT -3.565 -85.165 -3.235 -84.835 ;
        RECT -3.565 -87.885 -3.235 -87.555 ;
        RECT -3.565 -89.245 -3.235 -88.915 ;
        RECT -3.565 -90.605 -3.235 -90.275 ;
        RECT -3.565 -91.965 -3.235 -91.635 ;
        RECT -3.565 -93.325 -3.235 -92.995 ;
        RECT -3.565 -94.685 -3.235 -94.355 ;
        RECT -3.565 -96.045 -3.235 -95.715 ;
        RECT -3.565 -97.405 -3.235 -97.075 ;
        RECT -3.565 -98.765 -3.235 -98.435 ;
        RECT -3.565 -100.125 -3.235 -99.795 ;
        RECT -3.565 -101.485 -3.235 -101.155 ;
        RECT -3.565 -102.845 -3.235 -102.515 ;
        RECT -3.565 -104.205 -3.235 -103.875 ;
        RECT -3.565 -105.565 -3.235 -105.235 ;
        RECT -3.565 -106.925 -3.235 -106.595 ;
        RECT -3.565 -108.285 -3.235 -107.955 ;
        RECT -3.565 -109.645 -3.235 -109.315 ;
        RECT -3.565 -111.005 -3.235 -110.675 ;
        RECT -3.565 -112.365 -3.235 -112.035 ;
        RECT -3.565 -113.725 -3.235 -113.395 ;
        RECT -3.565 -115.085 -3.235 -114.755 ;
        RECT -3.565 -116.445 -3.235 -116.115 ;
        RECT -3.565 -117.805 -3.235 -117.475 ;
        RECT -3.565 -119.165 -3.235 -118.835 ;
        RECT -3.565 -120.525 -3.235 -120.195 ;
        RECT -3.565 -121.885 -3.235 -121.555 ;
        RECT -3.565 -123.245 -3.235 -122.915 ;
        RECT -3.565 -124.605 -3.235 -124.275 ;
        RECT -3.565 -125.965 -3.235 -125.635 ;
        RECT -3.565 -127.325 -3.235 -126.995 ;
        RECT -3.565 -128.685 -3.235 -128.355 ;
        RECT -3.565 -130.045 -3.235 -129.715 ;
        RECT -3.565 -131.405 -3.235 -131.075 ;
        RECT -3.565 -132.765 -3.235 -132.435 ;
        RECT -3.565 -134.125 -3.235 -133.795 ;
        RECT -3.565 -135.485 -3.235 -135.155 ;
        RECT -3.565 -136.845 -3.235 -136.515 ;
        RECT -3.565 -138.205 -3.235 -137.875 ;
        RECT -3.565 -139.565 -3.235 -139.235 ;
        RECT -3.565 -140.925 -3.235 -140.595 ;
        RECT -3.565 -142.285 -3.235 -141.955 ;
        RECT -3.565 -143.645 -3.235 -143.315 ;
        RECT -3.565 -145.005 -3.235 -144.675 ;
        RECT -3.565 -146.365 -3.235 -146.035 ;
        RECT -3.565 -147.725 -3.235 -147.395 ;
        RECT -3.565 -149.085 -3.235 -148.755 ;
        RECT -3.565 -150.445 -3.235 -150.115 ;
        RECT -3.565 -151.805 -3.235 -151.475 ;
        RECT -3.565 -153.165 -3.235 -152.835 ;
        RECT -3.565 -154.525 -3.235 -154.195 ;
        RECT -3.565 -155.885 -3.235 -155.555 ;
        RECT -3.565 -157.245 -3.235 -156.915 ;
        RECT -3.565 -158.605 -3.235 -158.275 ;
        RECT -3.565 -159.965 -3.235 -159.635 ;
        RECT -3.565 -161.325 -3.235 -160.995 ;
        RECT -3.565 -162.685 -3.235 -162.355 ;
        RECT -3.565 -164.045 -3.235 -163.715 ;
        RECT -3.565 -165.405 -3.235 -165.075 ;
        RECT -3.565 -166.765 -3.235 -166.435 ;
        RECT -3.565 -168.125 -3.235 -167.795 ;
        RECT -3.565 -169.485 -3.235 -169.155 ;
        RECT -3.565 -170.845 -3.235 -170.515 ;
        RECT -3.565 -172.205 -3.235 -171.875 ;
        RECT -3.565 -173.565 -3.235 -173.235 ;
        RECT -3.565 -174.925 -3.235 -174.595 ;
        RECT -3.565 -176.285 -3.235 -175.955 ;
        RECT -3.565 -177.645 -3.235 -177.315 ;
        RECT -3.565 -183.29 -3.235 -182.16 ;
        RECT -3.56 -183.405 -3.24 245.285 ;
        RECT -3.565 244.04 -3.235 245.17 ;
        RECT -3.565 239.875 -3.235 240.205 ;
        RECT -3.565 238.515 -3.235 238.845 ;
        RECT -3.565 237.155 -3.235 237.485 ;
        RECT -3.565 235.17 -3.235 235.5 ;
        RECT -3.565 232.995 -3.235 233.325 ;
        RECT -3.565 231.415 -3.235 231.745 ;
        RECT -3.565 230.565 -3.235 230.895 ;
        RECT -3.565 228.255 -3.235 228.585 ;
        RECT -3.565 227.405 -3.235 227.735 ;
        RECT -3.565 225.095 -3.235 225.425 ;
        RECT -3.565 224.245 -3.235 224.575 ;
        RECT -3.565 221.935 -3.235 222.265 ;
        RECT -3.565 221.085 -3.235 221.415 ;
        RECT -3.565 218.775 -3.235 219.105 ;
        RECT -3.565 217.195 -3.235 217.525 ;
        RECT -3.565 216.345 -3.235 216.675 ;
        RECT -3.565 214.035 -3.235 214.365 ;
        RECT -3.565 213.185 -3.235 213.515 ;
        RECT -3.565 210.875 -3.235 211.205 ;
        RECT -3.565 210.025 -3.235 210.355 ;
        RECT -3.565 207.715 -3.235 208.045 ;
        RECT -3.565 206.865 -3.235 207.195 ;
        RECT -3.565 204.555 -3.235 204.885 ;
        RECT -3.565 202.975 -3.235 203.305 ;
        RECT -3.565 202.125 -3.235 202.455 ;
        RECT -3.565 199.815 -3.235 200.145 ;
        RECT -3.565 198.965 -3.235 199.295 ;
        RECT -3.565 196.655 -3.235 196.985 ;
        RECT -3.565 195.805 -3.235 196.135 ;
        RECT -3.565 193.495 -3.235 193.825 ;
        RECT -3.565 192.645 -3.235 192.975 ;
        RECT -3.565 190.335 -3.235 190.665 ;
        RECT -3.565 188.755 -3.235 189.085 ;
        RECT -3.565 187.905 -3.235 188.235 ;
        RECT -3.565 185.595 -3.235 185.925 ;
        RECT -3.565 184.745 -3.235 185.075 ;
        RECT -3.565 182.435 -3.235 182.765 ;
        RECT -3.565 181.585 -3.235 181.915 ;
        RECT -3.565 179.275 -3.235 179.605 ;
        RECT -3.565 178.425 -3.235 178.755 ;
        RECT -3.565 176.115 -3.235 176.445 ;
        RECT -3.565 174.535 -3.235 174.865 ;
        RECT -3.565 173.685 -3.235 174.015 ;
        RECT -3.565 171.375 -3.235 171.705 ;
        RECT -3.565 170.525 -3.235 170.855 ;
        RECT -3.565 168.215 -3.235 168.545 ;
        RECT -3.565 167.365 -3.235 167.695 ;
        RECT -3.565 165.055 -3.235 165.385 ;
        RECT -3.565 164.205 -3.235 164.535 ;
        RECT -3.565 161.895 -3.235 162.225 ;
        RECT -3.565 160.315 -3.235 160.645 ;
        RECT -3.565 159.465 -3.235 159.795 ;
        RECT -3.565 157.155 -3.235 157.485 ;
        RECT -3.565 156.305 -3.235 156.635 ;
        RECT -3.565 153.995 -3.235 154.325 ;
        RECT -3.565 153.145 -3.235 153.475 ;
        RECT -3.565 150.835 -3.235 151.165 ;
        RECT -3.565 149.985 -3.235 150.315 ;
        RECT -3.565 147.675 -3.235 148.005 ;
        RECT -3.565 146.095 -3.235 146.425 ;
        RECT -3.565 145.245 -3.235 145.575 ;
        RECT -3.565 142.935 -3.235 143.265 ;
        RECT -3.565 142.085 -3.235 142.415 ;
        RECT -3.565 139.775 -3.235 140.105 ;
        RECT -3.565 138.925 -3.235 139.255 ;
        RECT -3.565 136.615 -3.235 136.945 ;
        RECT -3.565 135.765 -3.235 136.095 ;
        RECT -3.565 133.455 -3.235 133.785 ;
        RECT -3.565 131.875 -3.235 132.205 ;
        RECT -3.565 131.025 -3.235 131.355 ;
        RECT -3.565 128.715 -3.235 129.045 ;
        RECT -3.565 127.865 -3.235 128.195 ;
        RECT -3.565 125.555 -3.235 125.885 ;
        RECT -3.565 124.705 -3.235 125.035 ;
        RECT -3.565 122.395 -3.235 122.725 ;
    END
    PORT
      LAYER met3 ;
        RECT -15.805 -102.91 -15.475 -102.58 ;
        RECT -15.805 -104.205 -15.475 -103.875 ;
        RECT -15.805 -105.565 -15.475 -105.235 ;
        RECT -15.805 -108.285 -15.475 -107.955 ;
        RECT -15.8 -110.32 -15.48 -101.84 ;
    END
    PORT
      LAYER met3 ;
        RECT -15.805 -115.085 -15.475 -114.755 ;
        RECT -15.805 -116.445 -15.475 -116.115 ;
        RECT -15.805 -124.605 -15.475 -124.275 ;
        RECT -15.805 -125.965 -15.475 -125.635 ;
        RECT -15.805 -136.845 -15.475 -136.515 ;
        RECT -15.805 -140.925 -15.475 -140.595 ;
        RECT -15.805 -151.805 -15.475 -151.475 ;
        RECT -15.805 -157.245 -15.475 -156.915 ;
        RECT -15.805 -158.605 -15.475 -158.275 ;
        RECT -15.805 -159.965 -15.475 -159.635 ;
        RECT -15.805 -161.325 -15.475 -160.995 ;
        RECT -15.805 -162.685 -15.475 -162.355 ;
        RECT -15.805 -164.045 -15.475 -163.715 ;
        RECT -15.805 -165.405 -15.475 -165.075 ;
        RECT -15.805 -166.765 -15.475 -166.435 ;
        RECT -15.805 -168.655 -15.475 -168.325 ;
        RECT -15.805 -169.485 -15.475 -169.155 ;
        RECT -15.805 -170.845 -15.475 -170.515 ;
        RECT -15.805 -172.205 -15.475 -171.875 ;
        RECT -15.805 -173.565 -15.475 -173.235 ;
        RECT -15.805 -174.925 -15.475 -174.595 ;
        RECT -15.805 -177.645 -15.475 -177.315 ;
        RECT -15.805 -183.29 -15.475 -182.16 ;
        RECT -15.8 -183.405 -15.48 -114.08 ;
    END
    PORT
      LAYER met3 ;
        RECT -14.445 244.04 -14.115 245.17 ;
        RECT -14.445 239.875 -14.115 240.205 ;
        RECT -14.445 238.515 -14.115 238.845 ;
        RECT -14.445 237.155 -14.115 237.485 ;
        RECT -14.445 235.795 -14.115 236.125 ;
        RECT -14.445 234.435 -14.115 234.765 ;
        RECT -14.445 233.075 -14.115 233.405 ;
        RECT -14.445 231.715 -14.115 232.045 ;
        RECT -14.445 230.355 -14.115 230.685 ;
        RECT -14.445 228.995 -14.115 229.325 ;
        RECT -14.445 227.635 -14.115 227.965 ;
        RECT -14.445 226.275 -14.115 226.605 ;
        RECT -14.445 224.915 -14.115 225.245 ;
        RECT -14.445 223.555 -14.115 223.885 ;
        RECT -14.445 222.195 -14.115 222.525 ;
        RECT -14.445 220.835 -14.115 221.165 ;
        RECT -14.445 219.475 -14.115 219.805 ;
        RECT -14.445 218.115 -14.115 218.445 ;
        RECT -14.445 216.755 -14.115 217.085 ;
        RECT -14.445 215.395 -14.115 215.725 ;
        RECT -14.445 214.035 -14.115 214.365 ;
        RECT -14.445 212.675 -14.115 213.005 ;
        RECT -14.445 211.315 -14.115 211.645 ;
        RECT -14.445 209.955 -14.115 210.285 ;
        RECT -14.445 208.595 -14.115 208.925 ;
        RECT -14.445 207.235 -14.115 207.565 ;
        RECT -14.445 205.875 -14.115 206.205 ;
        RECT -14.445 204.515 -14.115 204.845 ;
        RECT -14.445 203.155 -14.115 203.485 ;
        RECT -14.445 201.795 -14.115 202.125 ;
        RECT -14.445 200.435 -14.115 200.765 ;
        RECT -14.445 199.075 -14.115 199.405 ;
        RECT -14.445 197.715 -14.115 198.045 ;
        RECT -14.445 196.355 -14.115 196.685 ;
        RECT -14.445 194.995 -14.115 195.325 ;
        RECT -14.445 193.635 -14.115 193.965 ;
        RECT -14.445 192.275 -14.115 192.605 ;
        RECT -14.445 190.915 -14.115 191.245 ;
        RECT -14.445 189.555 -14.115 189.885 ;
        RECT -14.445 188.195 -14.115 188.525 ;
        RECT -14.445 186.835 -14.115 187.165 ;
        RECT -14.445 185.475 -14.115 185.805 ;
        RECT -14.445 184.115 -14.115 184.445 ;
        RECT -14.445 182.755 -14.115 183.085 ;
        RECT -14.445 181.395 -14.115 181.725 ;
        RECT -14.445 180.035 -14.115 180.365 ;
        RECT -14.445 178.675 -14.115 179.005 ;
        RECT -14.445 177.315 -14.115 177.645 ;
        RECT -14.445 175.955 -14.115 176.285 ;
        RECT -14.445 174.595 -14.115 174.925 ;
        RECT -14.445 173.235 -14.115 173.565 ;
        RECT -14.445 171.875 -14.115 172.205 ;
        RECT -14.445 170.515 -14.115 170.845 ;
        RECT -14.445 169.155 -14.115 169.485 ;
        RECT -14.445 167.795 -14.115 168.125 ;
        RECT -14.445 166.435 -14.115 166.765 ;
        RECT -14.445 165.075 -14.115 165.405 ;
        RECT -14.445 163.715 -14.115 164.045 ;
        RECT -14.445 162.355 -14.115 162.685 ;
        RECT -14.445 160.995 -14.115 161.325 ;
        RECT -14.445 159.635 -14.115 159.965 ;
        RECT -14.445 158.275 -14.115 158.605 ;
        RECT -14.445 156.915 -14.115 157.245 ;
        RECT -14.445 155.555 -14.115 155.885 ;
        RECT -14.445 154.195 -14.115 154.525 ;
        RECT -14.445 152.835 -14.115 153.165 ;
        RECT -14.445 151.475 -14.115 151.805 ;
        RECT -14.445 150.115 -14.115 150.445 ;
        RECT -14.445 148.755 -14.115 149.085 ;
        RECT -14.445 147.395 -14.115 147.725 ;
        RECT -14.445 146.035 -14.115 146.365 ;
        RECT -14.445 144.675 -14.115 145.005 ;
        RECT -14.445 143.315 -14.115 143.645 ;
        RECT -14.445 141.955 -14.115 142.285 ;
        RECT -14.445 140.595 -14.115 140.925 ;
        RECT -14.445 139.235 -14.115 139.565 ;
        RECT -14.445 137.875 -14.115 138.205 ;
        RECT -14.445 136.515 -14.115 136.845 ;
        RECT -14.445 135.155 -14.115 135.485 ;
        RECT -14.445 133.795 -14.115 134.125 ;
        RECT -14.445 132.435 -14.115 132.765 ;
        RECT -14.445 131.075 -14.115 131.405 ;
        RECT -14.445 129.715 -14.115 130.045 ;
        RECT -14.445 128.355 -14.115 128.685 ;
        RECT -14.445 126.995 -14.115 127.325 ;
        RECT -14.445 125.635 -14.115 125.965 ;
        RECT -14.445 124.275 -14.115 124.605 ;
        RECT -14.445 122.915 -14.115 123.245 ;
        RECT -14.445 121.555 -14.115 121.885 ;
        RECT -14.445 120.195 -14.115 120.525 ;
        RECT -14.445 118.835 -14.115 119.165 ;
        RECT -14.445 117.475 -14.115 117.805 ;
        RECT -14.445 116.115 -14.115 116.445 ;
        RECT -14.445 114.755 -14.115 115.085 ;
        RECT -14.445 113.395 -14.115 113.725 ;
        RECT -14.445 112.035 -14.115 112.365 ;
        RECT -14.445 110.675 -14.115 111.005 ;
        RECT -14.445 109.315 -14.115 109.645 ;
        RECT -14.445 107.955 -14.115 108.285 ;
        RECT -14.445 106.595 -14.115 106.925 ;
        RECT -14.445 105.235 -14.115 105.565 ;
        RECT -14.445 103.875 -14.115 104.205 ;
        RECT -14.445 102.515 -14.115 102.845 ;
        RECT -14.445 101.155 -14.115 101.485 ;
        RECT -14.445 99.795 -14.115 100.125 ;
        RECT -14.445 98.435 -14.115 98.765 ;
        RECT -14.445 97.075 -14.115 97.405 ;
        RECT -14.445 95.715 -14.115 96.045 ;
        RECT -14.445 94.355 -14.115 94.685 ;
        RECT -14.445 92.995 -14.115 93.325 ;
        RECT -14.445 91.635 -14.115 91.965 ;
        RECT -14.445 90.275 -14.115 90.605 ;
        RECT -14.445 88.915 -14.115 89.245 ;
        RECT -14.445 87.555 -14.115 87.885 ;
        RECT -14.445 86.195 -14.115 86.525 ;
        RECT -14.445 84.835 -14.115 85.165 ;
        RECT -14.445 83.475 -14.115 83.805 ;
        RECT -14.445 82.115 -14.115 82.445 ;
        RECT -14.445 80.755 -14.115 81.085 ;
        RECT -14.445 79.395 -14.115 79.725 ;
        RECT -14.445 78.035 -14.115 78.365 ;
        RECT -14.445 76.675 -14.115 77.005 ;
        RECT -14.445 75.315 -14.115 75.645 ;
        RECT -14.445 73.955 -14.115 74.285 ;
        RECT -14.445 72.595 -14.115 72.925 ;
        RECT -14.445 71.235 -14.115 71.565 ;
        RECT -14.445 69.875 -14.115 70.205 ;
        RECT -14.445 68.515 -14.115 68.845 ;
        RECT -14.445 67.155 -14.115 67.485 ;
        RECT -14.445 65.795 -14.115 66.125 ;
        RECT -14.445 64.435 -14.115 64.765 ;
        RECT -14.445 63.075 -14.115 63.405 ;
        RECT -14.445 61.715 -14.115 62.045 ;
        RECT -14.445 60.355 -14.115 60.685 ;
        RECT -14.445 58.995 -14.115 59.325 ;
        RECT -14.445 57.635 -14.115 57.965 ;
        RECT -14.445 56.275 -14.115 56.605 ;
        RECT -14.445 54.915 -14.115 55.245 ;
        RECT -14.445 53.555 -14.115 53.885 ;
        RECT -14.445 52.195 -14.115 52.525 ;
        RECT -14.445 50.835 -14.115 51.165 ;
        RECT -14.445 49.475 -14.115 49.805 ;
        RECT -14.445 48.115 -14.115 48.445 ;
        RECT -14.445 46.755 -14.115 47.085 ;
        RECT -14.445 45.395 -14.115 45.725 ;
        RECT -14.445 44.035 -14.115 44.365 ;
        RECT -14.445 42.675 -14.115 43.005 ;
        RECT -14.445 41.315 -14.115 41.645 ;
        RECT -14.445 39.955 -14.115 40.285 ;
        RECT -14.445 38.595 -14.115 38.925 ;
        RECT -14.445 37.235 -14.115 37.565 ;
        RECT -14.445 35.875 -14.115 36.205 ;
        RECT -14.445 34.515 -14.115 34.845 ;
        RECT -14.445 33.155 -14.115 33.485 ;
        RECT -14.445 31.795 -14.115 32.125 ;
        RECT -14.445 30.435 -14.115 30.765 ;
        RECT -14.445 29.075 -14.115 29.405 ;
        RECT -14.445 27.715 -14.115 28.045 ;
        RECT -14.445 26.355 -14.115 26.685 ;
        RECT -14.445 24.995 -14.115 25.325 ;
        RECT -14.445 23.635 -14.115 23.965 ;
        RECT -14.445 22.275 -14.115 22.605 ;
        RECT -14.445 20.915 -14.115 21.245 ;
        RECT -14.445 19.555 -14.115 19.885 ;
        RECT -14.445 18.195 -14.115 18.525 ;
        RECT -14.445 16.835 -14.115 17.165 ;
        RECT -14.445 15.475 -14.115 15.805 ;
        RECT -14.445 14.115 -14.115 14.445 ;
        RECT -14.445 12.755 -14.115 13.085 ;
        RECT -14.445 11.395 -14.115 11.725 ;
        RECT -14.445 10.035 -14.115 10.365 ;
        RECT -14.445 8.675 -14.115 9.005 ;
        RECT -14.445 7.315 -14.115 7.645 ;
        RECT -14.445 5.955 -14.115 6.285 ;
        RECT -14.445 4.595 -14.115 4.925 ;
        RECT -14.445 3.235 -14.115 3.565 ;
        RECT -14.445 1.875 -14.115 2.205 ;
        RECT -14.445 0.515 -14.115 0.845 ;
        RECT -14.445 -0.845 -14.115 -0.515 ;
        RECT -14.445 -2.205 -14.115 -1.875 ;
        RECT -14.445 -3.565 -14.115 -3.235 ;
        RECT -14.445 -4.925 -14.115 -4.595 ;
        RECT -14.445 -7.645 -14.115 -7.315 ;
        RECT -14.445 -9.005 -14.115 -8.675 ;
        RECT -14.445 -10.73 -14.115 -10.4 ;
        RECT -14.445 -11.725 -14.115 -11.395 ;
        RECT -14.445 -13.085 -14.115 -12.755 ;
        RECT -14.445 -15.805 -14.115 -15.475 ;
        RECT -14.445 -16.77 -14.115 -16.44 ;
        RECT -14.445 -18.525 -14.115 -18.195 ;
        RECT -14.445 -21.245 -14.115 -20.915 ;
        RECT -14.445 -26.685 -14.115 -26.355 ;
        RECT -14.445 -28.045 -14.115 -27.715 ;
        RECT -14.445 -29.405 -14.115 -29.075 ;
        RECT -14.445 -30.765 -14.115 -30.435 ;
        RECT -14.445 -32.125 -14.115 -31.795 ;
        RECT -14.445 -33.71 -14.115 -33.38 ;
        RECT -14.445 -34.845 -14.115 -34.515 ;
        RECT -14.445 -36.205 -14.115 -35.875 ;
        RECT -14.445 -38.925 -14.115 -38.595 ;
        RECT -14.445 -39.75 -14.115 -39.42 ;
        RECT -14.445 -41.645 -14.115 -41.315 ;
        RECT -14.445 -44.365 -14.115 -44.035 ;
        RECT -14.445 -51.165 -14.115 -50.835 ;
        RECT -14.445 -52.525 -14.115 -52.195 ;
        RECT -14.445 -53.885 -14.115 -53.555 ;
        RECT -14.445 -55.245 -14.115 -54.915 ;
        RECT -14.445 -56.605 -14.115 -56.275 ;
        RECT -14.445 -57.965 -14.115 -57.635 ;
        RECT -14.445 -59.325 -14.115 -58.995 ;
        RECT -14.445 -60.685 -14.115 -60.355 ;
        RECT -14.445 -62.045 -14.115 -61.715 ;
        RECT -14.445 -63.405 -14.115 -63.075 ;
        RECT -14.445 -64.765 -14.115 -64.435 ;
        RECT -14.445 -66.125 -14.115 -65.795 ;
        RECT -14.445 -67.485 -14.115 -67.155 ;
        RECT -14.445 -68.845 -14.115 -68.515 ;
        RECT -14.445 -70.205 -14.115 -69.875 ;
        RECT -14.445 -71.565 -14.115 -71.235 ;
        RECT -14.445 -73.19 -14.115 -72.86 ;
        RECT -14.445 -74.285 -14.115 -73.955 ;
        RECT -14.445 -75.645 -14.115 -75.315 ;
        RECT -14.445 -78.365 -14.115 -78.035 ;
        RECT -14.445 -79.725 -14.115 -79.395 ;
        RECT -14.445 -80.73 -14.115 -80.4 ;
        RECT -14.445 -82.445 -14.115 -82.115 ;
        RECT -14.445 -83.805 -14.115 -83.475 ;
        RECT -14.445 -86.525 -14.115 -86.195 ;
        RECT -14.445 -89.245 -14.115 -88.915 ;
        RECT -14.445 -90.605 -14.115 -90.275 ;
        RECT -14.445 -91.965 -14.115 -91.635 ;
        RECT -14.445 -93.325 -14.115 -92.995 ;
        RECT -14.445 -94.685 -14.115 -94.355 ;
        RECT -14.445 -95.37 -14.115 -95.04 ;
        RECT -14.445 -97.405 -14.115 -97.075 ;
        RECT -14.445 -100.125 -14.115 -99.795 ;
        RECT -14.445 -101.485 -14.115 -101.155 ;
        RECT -14.445 -102.91 -14.115 -102.58 ;
        RECT -14.445 -104.205 -14.115 -103.875 ;
        RECT -14.445 -105.565 -14.115 -105.235 ;
        RECT -14.445 -108.285 -14.115 -107.955 ;
        RECT -14.44 -108.96 -14.12 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -14.445 -113.725 -14.115 -113.395 ;
        RECT -14.445 -115.085 -14.115 -114.755 ;
        RECT -14.445 -116.445 -14.115 -116.115 ;
        RECT -14.445 -119.165 -14.115 -118.835 ;
        RECT -14.445 -124.605 -14.115 -124.275 ;
        RECT -14.445 -132.765 -14.115 -132.435 ;
        RECT -14.445 -134.125 -14.115 -133.795 ;
        RECT -14.445 -136.845 -14.115 -136.515 ;
        RECT -14.445 -140.925 -14.115 -140.595 ;
        RECT -14.445 -142.285 -14.115 -141.955 ;
        RECT -14.445 -146.365 -14.115 -146.035 ;
        RECT -14.445 -147.725 -14.115 -147.395 ;
        RECT -14.445 -151.805 -14.115 -151.475 ;
        RECT -14.445 -154.525 -14.115 -154.195 ;
        RECT -14.445 -157.245 -14.115 -156.915 ;
        RECT -14.445 -158.605 -14.115 -158.275 ;
        RECT -14.445 -159.965 -14.115 -159.635 ;
        RECT -14.445 -161.325 -14.115 -160.995 ;
        RECT -14.445 -162.685 -14.115 -162.355 ;
        RECT -14.445 -164.045 -14.115 -163.715 ;
        RECT -14.445 -165.405 -14.115 -165.075 ;
        RECT -14.445 -166.765 -14.115 -166.435 ;
        RECT -14.445 -168.655 -14.115 -168.325 ;
        RECT -14.445 -169.485 -14.115 -169.155 ;
        RECT -14.445 -170.845 -14.115 -170.515 ;
        RECT -14.445 -173.565 -14.115 -173.235 ;
        RECT -14.445 -174.925 -14.115 -174.595 ;
        RECT -14.445 -177.645 -14.115 -177.315 ;
        RECT -14.445 -183.29 -14.115 -182.16 ;
        RECT -14.44 -183.405 -14.12 -112.72 ;
    END
    PORT
      LAYER met3 ;
        RECT -13.085 244.04 -12.755 245.17 ;
        RECT -13.085 239.875 -12.755 240.205 ;
        RECT -13.085 238.515 -12.755 238.845 ;
        RECT -13.085 237.155 -12.755 237.485 ;
        RECT -13.085 235.795 -12.755 236.125 ;
        RECT -13.085 234.435 -12.755 234.765 ;
        RECT -13.085 233.075 -12.755 233.405 ;
        RECT -13.085 231.715 -12.755 232.045 ;
        RECT -13.085 230.355 -12.755 230.685 ;
        RECT -13.085 228.995 -12.755 229.325 ;
        RECT -13.085 227.635 -12.755 227.965 ;
        RECT -13.085 226.275 -12.755 226.605 ;
        RECT -13.085 224.915 -12.755 225.245 ;
        RECT -13.085 223.555 -12.755 223.885 ;
        RECT -13.085 222.195 -12.755 222.525 ;
        RECT -13.085 220.835 -12.755 221.165 ;
        RECT -13.085 219.475 -12.755 219.805 ;
        RECT -13.085 218.115 -12.755 218.445 ;
        RECT -13.085 216.755 -12.755 217.085 ;
        RECT -13.085 215.395 -12.755 215.725 ;
        RECT -13.085 214.035 -12.755 214.365 ;
        RECT -13.085 212.675 -12.755 213.005 ;
        RECT -13.085 211.315 -12.755 211.645 ;
        RECT -13.085 209.955 -12.755 210.285 ;
        RECT -13.085 208.595 -12.755 208.925 ;
        RECT -13.085 207.235 -12.755 207.565 ;
        RECT -13.085 205.875 -12.755 206.205 ;
        RECT -13.085 204.515 -12.755 204.845 ;
        RECT -13.085 203.155 -12.755 203.485 ;
        RECT -13.085 201.795 -12.755 202.125 ;
        RECT -13.085 200.435 -12.755 200.765 ;
        RECT -13.085 199.075 -12.755 199.405 ;
        RECT -13.085 197.715 -12.755 198.045 ;
        RECT -13.085 196.355 -12.755 196.685 ;
        RECT -13.085 194.995 -12.755 195.325 ;
        RECT -13.085 193.635 -12.755 193.965 ;
        RECT -13.085 192.275 -12.755 192.605 ;
        RECT -13.085 190.915 -12.755 191.245 ;
        RECT -13.085 189.555 -12.755 189.885 ;
        RECT -13.085 188.195 -12.755 188.525 ;
        RECT -13.085 186.835 -12.755 187.165 ;
        RECT -13.085 185.475 -12.755 185.805 ;
        RECT -13.085 184.115 -12.755 184.445 ;
        RECT -13.085 182.755 -12.755 183.085 ;
        RECT -13.085 181.395 -12.755 181.725 ;
        RECT -13.085 180.035 -12.755 180.365 ;
        RECT -13.085 178.675 -12.755 179.005 ;
        RECT -13.085 177.315 -12.755 177.645 ;
        RECT -13.085 175.955 -12.755 176.285 ;
        RECT -13.085 174.595 -12.755 174.925 ;
        RECT -13.085 173.235 -12.755 173.565 ;
        RECT -13.085 171.875 -12.755 172.205 ;
        RECT -13.085 170.515 -12.755 170.845 ;
        RECT -13.085 169.155 -12.755 169.485 ;
        RECT -13.085 167.795 -12.755 168.125 ;
        RECT -13.085 166.435 -12.755 166.765 ;
        RECT -13.085 165.075 -12.755 165.405 ;
        RECT -13.085 163.715 -12.755 164.045 ;
        RECT -13.085 162.355 -12.755 162.685 ;
        RECT -13.085 160.995 -12.755 161.325 ;
        RECT -13.085 159.635 -12.755 159.965 ;
        RECT -13.085 158.275 -12.755 158.605 ;
        RECT -13.085 156.915 -12.755 157.245 ;
        RECT -13.085 155.555 -12.755 155.885 ;
        RECT -13.085 154.195 -12.755 154.525 ;
        RECT -13.085 152.835 -12.755 153.165 ;
        RECT -13.085 151.475 -12.755 151.805 ;
        RECT -13.085 150.115 -12.755 150.445 ;
        RECT -13.085 148.755 -12.755 149.085 ;
        RECT -13.085 147.395 -12.755 147.725 ;
        RECT -13.085 146.035 -12.755 146.365 ;
        RECT -13.085 144.675 -12.755 145.005 ;
        RECT -13.085 143.315 -12.755 143.645 ;
        RECT -13.085 141.955 -12.755 142.285 ;
        RECT -13.085 140.595 -12.755 140.925 ;
        RECT -13.085 139.235 -12.755 139.565 ;
        RECT -13.085 137.875 -12.755 138.205 ;
        RECT -13.085 136.515 -12.755 136.845 ;
        RECT -13.085 135.155 -12.755 135.485 ;
        RECT -13.085 133.795 -12.755 134.125 ;
        RECT -13.085 132.435 -12.755 132.765 ;
        RECT -13.085 131.075 -12.755 131.405 ;
        RECT -13.085 129.715 -12.755 130.045 ;
        RECT -13.085 128.355 -12.755 128.685 ;
        RECT -13.085 126.995 -12.755 127.325 ;
        RECT -13.085 125.635 -12.755 125.965 ;
        RECT -13.085 124.275 -12.755 124.605 ;
        RECT -13.085 122.915 -12.755 123.245 ;
        RECT -13.085 121.555 -12.755 121.885 ;
        RECT -13.085 120.195 -12.755 120.525 ;
        RECT -13.085 118.835 -12.755 119.165 ;
        RECT -13.085 117.475 -12.755 117.805 ;
        RECT -13.085 116.115 -12.755 116.445 ;
        RECT -13.085 114.755 -12.755 115.085 ;
        RECT -13.085 113.395 -12.755 113.725 ;
        RECT -13.085 112.035 -12.755 112.365 ;
        RECT -13.085 110.675 -12.755 111.005 ;
        RECT -13.085 109.315 -12.755 109.645 ;
        RECT -13.085 107.955 -12.755 108.285 ;
        RECT -13.085 106.595 -12.755 106.925 ;
        RECT -13.085 105.235 -12.755 105.565 ;
        RECT -13.085 103.875 -12.755 104.205 ;
        RECT -13.085 102.515 -12.755 102.845 ;
        RECT -13.085 101.155 -12.755 101.485 ;
        RECT -13.085 99.795 -12.755 100.125 ;
        RECT -13.085 98.435 -12.755 98.765 ;
        RECT -13.085 97.075 -12.755 97.405 ;
        RECT -13.085 95.715 -12.755 96.045 ;
        RECT -13.085 94.355 -12.755 94.685 ;
        RECT -13.085 92.995 -12.755 93.325 ;
        RECT -13.085 91.635 -12.755 91.965 ;
        RECT -13.085 90.275 -12.755 90.605 ;
        RECT -13.085 88.915 -12.755 89.245 ;
        RECT -13.085 87.555 -12.755 87.885 ;
        RECT -13.085 86.195 -12.755 86.525 ;
        RECT -13.085 84.835 -12.755 85.165 ;
        RECT -13.085 83.475 -12.755 83.805 ;
        RECT -13.085 82.115 -12.755 82.445 ;
        RECT -13.085 80.755 -12.755 81.085 ;
        RECT -13.085 79.395 -12.755 79.725 ;
        RECT -13.085 78.035 -12.755 78.365 ;
        RECT -13.085 76.675 -12.755 77.005 ;
        RECT -13.085 75.315 -12.755 75.645 ;
        RECT -13.085 73.955 -12.755 74.285 ;
        RECT -13.085 72.595 -12.755 72.925 ;
        RECT -13.085 71.235 -12.755 71.565 ;
        RECT -13.085 69.875 -12.755 70.205 ;
        RECT -13.085 68.515 -12.755 68.845 ;
        RECT -13.085 67.155 -12.755 67.485 ;
        RECT -13.085 65.795 -12.755 66.125 ;
        RECT -13.085 64.435 -12.755 64.765 ;
        RECT -13.085 63.075 -12.755 63.405 ;
        RECT -13.085 61.715 -12.755 62.045 ;
        RECT -13.085 60.355 -12.755 60.685 ;
        RECT -13.085 58.995 -12.755 59.325 ;
        RECT -13.085 57.635 -12.755 57.965 ;
        RECT -13.085 56.275 -12.755 56.605 ;
        RECT -13.085 54.915 -12.755 55.245 ;
        RECT -13.085 53.555 -12.755 53.885 ;
        RECT -13.085 52.195 -12.755 52.525 ;
        RECT -13.085 50.835 -12.755 51.165 ;
        RECT -13.085 49.475 -12.755 49.805 ;
        RECT -13.085 48.115 -12.755 48.445 ;
        RECT -13.085 46.755 -12.755 47.085 ;
        RECT -13.085 45.395 -12.755 45.725 ;
        RECT -13.085 44.035 -12.755 44.365 ;
        RECT -13.085 42.675 -12.755 43.005 ;
        RECT -13.085 41.315 -12.755 41.645 ;
        RECT -13.085 39.955 -12.755 40.285 ;
        RECT -13.085 38.595 -12.755 38.925 ;
        RECT -13.085 37.235 -12.755 37.565 ;
        RECT -13.085 35.875 -12.755 36.205 ;
        RECT -13.085 34.515 -12.755 34.845 ;
        RECT -13.085 33.155 -12.755 33.485 ;
        RECT -13.085 31.795 -12.755 32.125 ;
        RECT -13.085 30.435 -12.755 30.765 ;
        RECT -13.085 29.075 -12.755 29.405 ;
        RECT -13.085 27.715 -12.755 28.045 ;
        RECT -13.085 26.355 -12.755 26.685 ;
        RECT -13.085 24.995 -12.755 25.325 ;
        RECT -13.085 23.635 -12.755 23.965 ;
        RECT -13.085 22.275 -12.755 22.605 ;
        RECT -13.085 20.915 -12.755 21.245 ;
        RECT -13.085 19.555 -12.755 19.885 ;
        RECT -13.085 18.195 -12.755 18.525 ;
        RECT -13.085 16.835 -12.755 17.165 ;
        RECT -13.085 15.475 -12.755 15.805 ;
        RECT -13.085 14.115 -12.755 14.445 ;
        RECT -13.085 12.755 -12.755 13.085 ;
        RECT -13.085 11.395 -12.755 11.725 ;
        RECT -13.085 10.035 -12.755 10.365 ;
        RECT -13.085 8.675 -12.755 9.005 ;
        RECT -13.085 7.315 -12.755 7.645 ;
        RECT -13.085 5.955 -12.755 6.285 ;
        RECT -13.085 4.595 -12.755 4.925 ;
        RECT -13.085 3.235 -12.755 3.565 ;
        RECT -13.085 1.875 -12.755 2.205 ;
        RECT -13.085 0.515 -12.755 0.845 ;
        RECT -13.085 -0.845 -12.755 -0.515 ;
        RECT -13.085 -2.205 -12.755 -1.875 ;
        RECT -13.085 -3.565 -12.755 -3.235 ;
        RECT -13.085 -4.925 -12.755 -4.595 ;
        RECT -13.085 -7.645 -12.755 -7.315 ;
        RECT -13.085 -9.005 -12.755 -8.675 ;
        RECT -13.085 -10.73 -12.755 -10.4 ;
        RECT -13.085 -11.725 -12.755 -11.395 ;
        RECT -13.085 -13.085 -12.755 -12.755 ;
        RECT -13.085 -15.805 -12.755 -15.475 ;
        RECT -13.085 -16.77 -12.755 -16.44 ;
        RECT -13.08 -17.84 -12.76 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -13.085 -112.365 -12.755 -112.035 ;
        RECT -13.085 -113.725 -12.755 -113.395 ;
        RECT -13.085 -115.085 -12.755 -114.755 ;
        RECT -13.085 -116.445 -12.755 -116.115 ;
        RECT -13.085 -117.805 -12.755 -117.475 ;
        RECT -13.085 -119.165 -12.755 -118.835 ;
        RECT -13.085 -134.125 -12.755 -133.795 ;
        RECT -13.085 -136.845 -12.755 -136.515 ;
        RECT -13.085 -140.925 -12.755 -140.595 ;
        RECT -13.085 -142.285 -12.755 -141.955 ;
        RECT -13.085 -146.365 -12.755 -146.035 ;
        RECT -13.085 -147.725 -12.755 -147.395 ;
        RECT -13.085 -149.085 -12.755 -148.755 ;
        RECT -13.085 -151.805 -12.755 -151.475 ;
        RECT -13.085 -153.165 -12.755 -152.835 ;
        RECT -13.085 -154.525 -12.755 -154.195 ;
        RECT -13.085 -155.885 -12.755 -155.555 ;
        RECT -13.085 -157.245 -12.755 -156.915 ;
        RECT -13.085 -158.605 -12.755 -158.275 ;
        RECT -13.085 -159.965 -12.755 -159.635 ;
        RECT -13.085 -161.325 -12.755 -160.995 ;
        RECT -13.085 -162.685 -12.755 -162.355 ;
        RECT -13.085 -164.045 -12.755 -163.715 ;
        RECT -13.085 -165.405 -12.755 -165.075 ;
        RECT -13.085 -166.765 -12.755 -166.435 ;
        RECT -13.085 -168.655 -12.755 -168.325 ;
        RECT -13.085 -169.485 -12.755 -169.155 ;
        RECT -13.085 -170.845 -12.755 -170.515 ;
        RECT -13.085 -172.205 -12.755 -171.875 ;
        RECT -13.085 -173.565 -12.755 -173.235 ;
        RECT -13.085 -174.925 -12.755 -174.595 ;
        RECT -13.085 -177.645 -12.755 -177.315 ;
        RECT -13.085 -183.29 -12.755 -182.16 ;
        RECT -13.08 -183.405 -12.76 -108.64 ;
    END
    PORT
      LAYER met3 ;
        RECT -11.725 244.04 -11.395 245.17 ;
        RECT -11.725 239.875 -11.395 240.205 ;
        RECT -11.725 238.515 -11.395 238.845 ;
        RECT -11.725 237.155 -11.395 237.485 ;
        RECT -11.725 235.795 -11.395 236.125 ;
        RECT -11.725 234.435 -11.395 234.765 ;
        RECT -11.725 233.075 -11.395 233.405 ;
        RECT -11.725 231.715 -11.395 232.045 ;
        RECT -11.725 230.355 -11.395 230.685 ;
        RECT -11.725 228.995 -11.395 229.325 ;
        RECT -11.725 227.635 -11.395 227.965 ;
        RECT -11.725 226.275 -11.395 226.605 ;
        RECT -11.725 224.915 -11.395 225.245 ;
        RECT -11.725 223.555 -11.395 223.885 ;
        RECT -11.725 222.195 -11.395 222.525 ;
        RECT -11.725 220.835 -11.395 221.165 ;
        RECT -11.725 219.475 -11.395 219.805 ;
        RECT -11.725 218.115 -11.395 218.445 ;
        RECT -11.725 216.755 -11.395 217.085 ;
        RECT -11.725 215.395 -11.395 215.725 ;
        RECT -11.725 214.035 -11.395 214.365 ;
        RECT -11.725 212.675 -11.395 213.005 ;
        RECT -11.725 211.315 -11.395 211.645 ;
        RECT -11.725 209.955 -11.395 210.285 ;
        RECT -11.725 208.595 -11.395 208.925 ;
        RECT -11.725 207.235 -11.395 207.565 ;
        RECT -11.725 205.875 -11.395 206.205 ;
        RECT -11.725 204.515 -11.395 204.845 ;
        RECT -11.725 203.155 -11.395 203.485 ;
        RECT -11.725 201.795 -11.395 202.125 ;
        RECT -11.725 200.435 -11.395 200.765 ;
        RECT -11.725 199.075 -11.395 199.405 ;
        RECT -11.725 197.715 -11.395 198.045 ;
        RECT -11.725 196.355 -11.395 196.685 ;
        RECT -11.725 194.995 -11.395 195.325 ;
        RECT -11.725 193.635 -11.395 193.965 ;
        RECT -11.725 192.275 -11.395 192.605 ;
        RECT -11.725 190.915 -11.395 191.245 ;
        RECT -11.725 189.555 -11.395 189.885 ;
        RECT -11.725 188.195 -11.395 188.525 ;
        RECT -11.725 186.835 -11.395 187.165 ;
        RECT -11.725 185.475 -11.395 185.805 ;
        RECT -11.725 184.115 -11.395 184.445 ;
        RECT -11.725 182.755 -11.395 183.085 ;
        RECT -11.725 181.395 -11.395 181.725 ;
        RECT -11.725 180.035 -11.395 180.365 ;
        RECT -11.725 178.675 -11.395 179.005 ;
        RECT -11.725 177.315 -11.395 177.645 ;
        RECT -11.725 175.955 -11.395 176.285 ;
        RECT -11.725 174.595 -11.395 174.925 ;
        RECT -11.725 173.235 -11.395 173.565 ;
        RECT -11.725 171.875 -11.395 172.205 ;
        RECT -11.725 170.515 -11.395 170.845 ;
        RECT -11.725 169.155 -11.395 169.485 ;
        RECT -11.725 167.795 -11.395 168.125 ;
        RECT -11.725 166.435 -11.395 166.765 ;
        RECT -11.725 165.075 -11.395 165.405 ;
        RECT -11.725 163.715 -11.395 164.045 ;
        RECT -11.725 162.355 -11.395 162.685 ;
        RECT -11.725 160.995 -11.395 161.325 ;
        RECT -11.725 159.635 -11.395 159.965 ;
        RECT -11.725 158.275 -11.395 158.605 ;
        RECT -11.725 156.915 -11.395 157.245 ;
        RECT -11.725 155.555 -11.395 155.885 ;
        RECT -11.725 154.195 -11.395 154.525 ;
        RECT -11.725 152.835 -11.395 153.165 ;
        RECT -11.725 151.475 -11.395 151.805 ;
        RECT -11.725 150.115 -11.395 150.445 ;
        RECT -11.725 148.755 -11.395 149.085 ;
        RECT -11.725 147.395 -11.395 147.725 ;
        RECT -11.725 146.035 -11.395 146.365 ;
        RECT -11.725 144.675 -11.395 145.005 ;
        RECT -11.725 143.315 -11.395 143.645 ;
        RECT -11.725 141.955 -11.395 142.285 ;
        RECT -11.725 140.595 -11.395 140.925 ;
        RECT -11.725 139.235 -11.395 139.565 ;
        RECT -11.725 137.875 -11.395 138.205 ;
        RECT -11.725 136.515 -11.395 136.845 ;
        RECT -11.725 135.155 -11.395 135.485 ;
        RECT -11.725 133.795 -11.395 134.125 ;
        RECT -11.725 132.435 -11.395 132.765 ;
        RECT -11.725 131.075 -11.395 131.405 ;
        RECT -11.725 129.715 -11.395 130.045 ;
        RECT -11.725 128.355 -11.395 128.685 ;
        RECT -11.725 126.995 -11.395 127.325 ;
        RECT -11.725 125.635 -11.395 125.965 ;
        RECT -11.725 124.275 -11.395 124.605 ;
        RECT -11.725 122.915 -11.395 123.245 ;
        RECT -11.725 121.555 -11.395 121.885 ;
        RECT -11.725 120.195 -11.395 120.525 ;
        RECT -11.725 118.835 -11.395 119.165 ;
        RECT -11.725 117.475 -11.395 117.805 ;
        RECT -11.725 116.115 -11.395 116.445 ;
        RECT -11.725 114.755 -11.395 115.085 ;
        RECT -11.725 113.395 -11.395 113.725 ;
        RECT -11.725 112.035 -11.395 112.365 ;
        RECT -11.725 110.675 -11.395 111.005 ;
        RECT -11.725 109.315 -11.395 109.645 ;
        RECT -11.725 107.955 -11.395 108.285 ;
        RECT -11.725 106.595 -11.395 106.925 ;
        RECT -11.725 105.235 -11.395 105.565 ;
        RECT -11.725 103.875 -11.395 104.205 ;
        RECT -11.725 102.515 -11.395 102.845 ;
        RECT -11.725 101.155 -11.395 101.485 ;
        RECT -11.725 99.795 -11.395 100.125 ;
        RECT -11.725 98.435 -11.395 98.765 ;
        RECT -11.725 97.075 -11.395 97.405 ;
        RECT -11.725 95.715 -11.395 96.045 ;
        RECT -11.725 94.355 -11.395 94.685 ;
        RECT -11.725 92.995 -11.395 93.325 ;
        RECT -11.725 91.635 -11.395 91.965 ;
        RECT -11.725 90.275 -11.395 90.605 ;
        RECT -11.725 88.915 -11.395 89.245 ;
        RECT -11.725 87.555 -11.395 87.885 ;
        RECT -11.725 86.195 -11.395 86.525 ;
        RECT -11.725 84.835 -11.395 85.165 ;
        RECT -11.725 83.475 -11.395 83.805 ;
        RECT -11.725 82.115 -11.395 82.445 ;
        RECT -11.725 80.755 -11.395 81.085 ;
        RECT -11.725 79.395 -11.395 79.725 ;
        RECT -11.725 78.035 -11.395 78.365 ;
        RECT -11.725 76.675 -11.395 77.005 ;
        RECT -11.725 75.315 -11.395 75.645 ;
        RECT -11.725 73.955 -11.395 74.285 ;
        RECT -11.725 72.595 -11.395 72.925 ;
        RECT -11.725 71.235 -11.395 71.565 ;
        RECT -11.725 69.875 -11.395 70.205 ;
        RECT -11.725 68.515 -11.395 68.845 ;
        RECT -11.725 67.155 -11.395 67.485 ;
        RECT -11.725 65.795 -11.395 66.125 ;
        RECT -11.725 64.435 -11.395 64.765 ;
        RECT -11.725 63.075 -11.395 63.405 ;
        RECT -11.725 61.715 -11.395 62.045 ;
        RECT -11.725 60.355 -11.395 60.685 ;
        RECT -11.725 58.995 -11.395 59.325 ;
        RECT -11.725 57.635 -11.395 57.965 ;
        RECT -11.725 56.275 -11.395 56.605 ;
        RECT -11.725 54.915 -11.395 55.245 ;
        RECT -11.725 53.555 -11.395 53.885 ;
        RECT -11.725 52.195 -11.395 52.525 ;
        RECT -11.725 50.835 -11.395 51.165 ;
        RECT -11.725 49.475 -11.395 49.805 ;
        RECT -11.725 48.115 -11.395 48.445 ;
        RECT -11.725 46.755 -11.395 47.085 ;
        RECT -11.725 45.395 -11.395 45.725 ;
        RECT -11.725 44.035 -11.395 44.365 ;
        RECT -11.725 42.675 -11.395 43.005 ;
        RECT -11.725 41.315 -11.395 41.645 ;
        RECT -11.725 39.955 -11.395 40.285 ;
        RECT -11.725 38.595 -11.395 38.925 ;
        RECT -11.725 37.235 -11.395 37.565 ;
        RECT -11.725 35.875 -11.395 36.205 ;
        RECT -11.725 34.515 -11.395 34.845 ;
        RECT -11.725 33.155 -11.395 33.485 ;
        RECT -11.725 31.795 -11.395 32.125 ;
        RECT -11.725 30.435 -11.395 30.765 ;
        RECT -11.725 29.075 -11.395 29.405 ;
        RECT -11.725 27.715 -11.395 28.045 ;
        RECT -11.725 26.355 -11.395 26.685 ;
        RECT -11.725 24.995 -11.395 25.325 ;
        RECT -11.725 23.635 -11.395 23.965 ;
        RECT -11.725 22.275 -11.395 22.605 ;
        RECT -11.725 20.915 -11.395 21.245 ;
        RECT -11.725 19.555 -11.395 19.885 ;
        RECT -11.725 18.195 -11.395 18.525 ;
        RECT -11.725 16.835 -11.395 17.165 ;
        RECT -11.725 15.475 -11.395 15.805 ;
        RECT -11.725 14.115 -11.395 14.445 ;
        RECT -11.725 12.755 -11.395 13.085 ;
        RECT -11.725 11.395 -11.395 11.725 ;
        RECT -11.725 10.035 -11.395 10.365 ;
        RECT -11.725 8.675 -11.395 9.005 ;
        RECT -11.725 7.315 -11.395 7.645 ;
        RECT -11.725 5.955 -11.395 6.285 ;
        RECT -11.725 4.595 -11.395 4.925 ;
        RECT -11.725 3.235 -11.395 3.565 ;
        RECT -11.725 1.875 -11.395 2.205 ;
        RECT -11.725 0.515 -11.395 0.845 ;
        RECT -11.725 -0.845 -11.395 -0.515 ;
        RECT -11.725 -2.205 -11.395 -1.875 ;
        RECT -11.725 -3.565 -11.395 -3.235 ;
        RECT -11.725 -4.925 -11.395 -4.595 ;
        RECT -11.725 -6.285 -11.395 -5.955 ;
        RECT -11.725 -7.645 -11.395 -7.315 ;
        RECT -11.725 -9.005 -11.395 -8.675 ;
        RECT -11.725 -10.73 -11.395 -10.4 ;
        RECT -11.725 -11.725 -11.395 -11.395 ;
        RECT -11.725 -13.085 -11.395 -12.755 ;
        RECT -11.725 -15.805 -11.395 -15.475 ;
        RECT -11.725 -16.77 -11.395 -16.44 ;
        RECT -11.725 -21.245 -11.395 -20.915 ;
        RECT -11.725 -26.685 -11.395 -26.355 ;
        RECT -11.725 -28.045 -11.395 -27.715 ;
        RECT -11.725 -29.405 -11.395 -29.075 ;
        RECT -11.725 -30.765 -11.395 -30.435 ;
        RECT -11.725 -32.125 -11.395 -31.795 ;
        RECT -11.725 -33.71 -11.395 -33.38 ;
        RECT -11.725 -36.205 -11.395 -35.875 ;
        RECT -11.725 -38.925 -11.395 -38.595 ;
        RECT -11.725 -39.75 -11.395 -39.42 ;
        RECT -11.725 -41.645 -11.395 -41.315 ;
        RECT -11.725 -44.365 -11.395 -44.035 ;
        RECT -11.725 -51.165 -11.395 -50.835 ;
        RECT -11.725 -52.525 -11.395 -52.195 ;
        RECT -11.725 -53.885 -11.395 -53.555 ;
        RECT -11.725 -55.245 -11.395 -54.915 ;
        RECT -11.725 -56.605 -11.395 -56.275 ;
        RECT -11.725 -57.965 -11.395 -57.635 ;
        RECT -11.725 -59.325 -11.395 -58.995 ;
        RECT -11.725 -60.685 -11.395 -60.355 ;
        RECT -11.725 -62.045 -11.395 -61.715 ;
        RECT -11.725 -63.405 -11.395 -63.075 ;
        RECT -11.725 -64.765 -11.395 -64.435 ;
        RECT -11.725 -66.125 -11.395 -65.795 ;
        RECT -11.725 -67.485 -11.395 -67.155 ;
        RECT -11.725 -68.845 -11.395 -68.515 ;
        RECT -11.725 -70.205 -11.395 -69.875 ;
        RECT -11.725 -71.565 -11.395 -71.235 ;
        RECT -11.725 -73.19 -11.395 -72.86 ;
        RECT -11.725 -74.285 -11.395 -73.955 ;
        RECT -11.725 -75.645 -11.395 -75.315 ;
        RECT -11.725 -78.365 -11.395 -78.035 ;
        RECT -11.725 -79.725 -11.395 -79.395 ;
        RECT -11.725 -80.73 -11.395 -80.4 ;
        RECT -11.725 -82.445 -11.395 -82.115 ;
        RECT -11.725 -83.805 -11.395 -83.475 ;
        RECT -11.725 -86.525 -11.395 -86.195 ;
        RECT -11.725 -89.245 -11.395 -88.915 ;
        RECT -11.725 -90.605 -11.395 -90.275 ;
        RECT -11.725 -91.965 -11.395 -91.635 ;
        RECT -11.725 -93.325 -11.395 -92.995 ;
        RECT -11.725 -94.685 -11.395 -94.355 ;
        RECT -11.725 -95.37 -11.395 -95.04 ;
        RECT -11.725 -97.405 -11.395 -97.075 ;
        RECT -11.725 -100.125 -11.395 -99.795 ;
        RECT -11.725 -102.91 -11.395 -102.58 ;
        RECT -11.725 -104.205 -11.395 -103.875 ;
        RECT -11.725 -105.565 -11.395 -105.235 ;
        RECT -11.725 -108.285 -11.395 -107.955 ;
        RECT -11.725 -112.365 -11.395 -112.035 ;
        RECT -11.725 -113.725 -11.395 -113.395 ;
        RECT -11.725 -115.085 -11.395 -114.755 ;
        RECT -11.725 -116.445 -11.395 -116.115 ;
        RECT -11.725 -117.805 -11.395 -117.475 ;
        RECT -11.725 -119.165 -11.395 -118.835 ;
        RECT -11.725 -125.965 -11.395 -125.635 ;
        RECT -11.725 -127.325 -11.395 -126.995 ;
        RECT -11.725 -130.045 -11.395 -129.715 ;
        RECT -11.725 -131.405 -11.395 -131.075 ;
        RECT -11.725 -134.125 -11.395 -133.795 ;
        RECT -11.725 -135.485 -11.395 -135.155 ;
        RECT -11.725 -136.845 -11.395 -136.515 ;
        RECT -11.725 -138.205 -11.395 -137.875 ;
        RECT -11.725 -139.565 -11.395 -139.235 ;
        RECT -11.725 -140.925 -11.395 -140.595 ;
        RECT -11.725 -142.285 -11.395 -141.955 ;
        RECT -11.725 -146.365 -11.395 -146.035 ;
        RECT -11.725 -147.725 -11.395 -147.395 ;
        RECT -11.725 -149.085 -11.395 -148.755 ;
        RECT -11.725 -150.445 -11.395 -150.115 ;
        RECT -11.725 -151.805 -11.395 -151.475 ;
        RECT -11.725 -153.165 -11.395 -152.835 ;
        RECT -11.725 -154.525 -11.395 -154.195 ;
        RECT -11.725 -155.885 -11.395 -155.555 ;
        RECT -11.725 -157.245 -11.395 -156.915 ;
        RECT -11.725 -158.605 -11.395 -158.275 ;
        RECT -11.725 -159.965 -11.395 -159.635 ;
        RECT -11.725 -161.325 -11.395 -160.995 ;
        RECT -11.725 -162.685 -11.395 -162.355 ;
        RECT -11.725 -164.045 -11.395 -163.715 ;
        RECT -11.725 -165.405 -11.395 -165.075 ;
        RECT -11.725 -166.765 -11.395 -166.435 ;
        RECT -11.725 -168.655 -11.395 -168.325 ;
        RECT -11.725 -169.485 -11.395 -169.155 ;
        RECT -11.725 -170.845 -11.395 -170.515 ;
        RECT -11.725 -172.205 -11.395 -171.875 ;
        RECT -11.725 -173.565 -11.395 -173.235 ;
        RECT -11.725 -174.925 -11.395 -174.595 ;
        RECT -11.725 -177.645 -11.395 -177.315 ;
        RECT -11.725 -183.29 -11.395 -182.16 ;
        RECT -11.72 -183.405 -11.4 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -10.365 46.755 -10.035 47.085 ;
        RECT -10.365 42.675 -10.035 43.005 ;
        RECT -10.365 39.955 -10.035 40.285 ;
        RECT -10.365 33.155 -10.035 33.485 ;
        RECT -10.365 31.795 -10.035 32.125 ;
        RECT -10.365 29.075 -10.035 29.405 ;
        RECT -10.365 22.275 -10.035 22.605 ;
        RECT -10.365 19.555 -10.035 19.885 ;
        RECT -10.365 18.195 -10.035 18.525 ;
        RECT -10.365 11.395 -10.035 11.725 ;
        RECT -10.365 4.595 -10.035 4.925 ;
        RECT -10.365 3.235 -10.035 3.565 ;
        RECT -10.365 1.875 -10.035 2.205 ;
        RECT -10.365 0.515 -10.035 0.845 ;
        RECT -10.365 -0.845 -10.035 -0.515 ;
        RECT -10.365 -2.205 -10.035 -1.875 ;
        RECT -10.365 -3.565 -10.035 -3.235 ;
        RECT -10.365 -4.925 -10.035 -4.595 ;
        RECT -10.365 -6.285 -10.035 -5.955 ;
        RECT -10.365 -7.645 -10.035 -7.315 ;
        RECT -10.365 -9.005 -10.035 -8.675 ;
        RECT -10.365 -10.73 -10.035 -10.4 ;
        RECT -10.365 -11.725 -10.035 -11.395 ;
        RECT -10.365 -13.085 -10.035 -12.755 ;
        RECT -10.365 -15.805 -10.035 -15.475 ;
        RECT -10.365 -16.77 -10.035 -16.44 ;
        RECT -10.365 -21.245 -10.035 -20.915 ;
        RECT -10.365 -26.685 -10.035 -26.355 ;
        RECT -10.365 -28.045 -10.035 -27.715 ;
        RECT -10.365 -29.405 -10.035 -29.075 ;
        RECT -10.365 -30.765 -10.035 -30.435 ;
        RECT -10.365 -32.125 -10.035 -31.795 ;
        RECT -10.365 -33.71 -10.035 -33.38 ;
        RECT -10.365 -36.205 -10.035 -35.875 ;
        RECT -10.365 -38.925 -10.035 -38.595 ;
        RECT -10.365 -39.75 -10.035 -39.42 ;
        RECT -10.365 -41.645 -10.035 -41.315 ;
        RECT -10.365 -44.365 -10.035 -44.035 ;
        RECT -10.365 -51.165 -10.035 -50.835 ;
        RECT -10.365 -52.525 -10.035 -52.195 ;
        RECT -10.365 -53.885 -10.035 -53.555 ;
        RECT -10.365 -55.245 -10.035 -54.915 ;
        RECT -10.365 -56.605 -10.035 -56.275 ;
        RECT -10.365 -57.965 -10.035 -57.635 ;
        RECT -10.365 -59.325 -10.035 -58.995 ;
        RECT -10.365 -60.685 -10.035 -60.355 ;
        RECT -10.365 -62.045 -10.035 -61.715 ;
        RECT -10.365 -63.405 -10.035 -63.075 ;
        RECT -10.365 -64.765 -10.035 -64.435 ;
        RECT -10.365 -66.125 -10.035 -65.795 ;
        RECT -10.365 -67.485 -10.035 -67.155 ;
        RECT -10.365 -68.845 -10.035 -68.515 ;
        RECT -10.365 -70.205 -10.035 -69.875 ;
        RECT -10.365 -71.565 -10.035 -71.235 ;
        RECT -10.365 -73.19 -10.035 -72.86 ;
        RECT -10.365 -74.285 -10.035 -73.955 ;
        RECT -10.365 -75.645 -10.035 -75.315 ;
        RECT -10.365 -78.365 -10.035 -78.035 ;
        RECT -10.365 -79.725 -10.035 -79.395 ;
        RECT -10.365 -80.73 -10.035 -80.4 ;
        RECT -10.365 -82.445 -10.035 -82.115 ;
        RECT -10.365 -83.805 -10.035 -83.475 ;
        RECT -10.365 -86.525 -10.035 -86.195 ;
        RECT -10.365 -89.245 -10.035 -88.915 ;
        RECT -10.365 -90.605 -10.035 -90.275 ;
        RECT -10.365 -91.965 -10.035 -91.635 ;
        RECT -10.365 -93.325 -10.035 -92.995 ;
        RECT -10.365 -94.685 -10.035 -94.355 ;
        RECT -10.365 -95.37 -10.035 -95.04 ;
        RECT -10.365 -97.405 -10.035 -97.075 ;
        RECT -10.365 -100.125 -10.035 -99.795 ;
        RECT -10.365 -102.91 -10.035 -102.58 ;
        RECT -10.365 -104.205 -10.035 -103.875 ;
        RECT -10.365 -105.565 -10.035 -105.235 ;
        RECT -10.365 -108.285 -10.035 -107.955 ;
        RECT -10.365 -112.365 -10.035 -112.035 ;
        RECT -10.365 -113.725 -10.035 -113.395 ;
        RECT -10.365 -115.085 -10.035 -114.755 ;
        RECT -10.365 -116.445 -10.035 -116.115 ;
        RECT -10.365 -117.805 -10.035 -117.475 ;
        RECT -10.365 -119.165 -10.035 -118.835 ;
        RECT -10.365 -124.605 -10.035 -124.275 ;
        RECT -10.365 -125.965 -10.035 -125.635 ;
        RECT -10.365 -127.325 -10.035 -126.995 ;
        RECT -10.365 -128.685 -10.035 -128.355 ;
        RECT -10.365 -130.045 -10.035 -129.715 ;
        RECT -10.365 -131.405 -10.035 -131.075 ;
        RECT -10.365 -134.125 -10.035 -133.795 ;
        RECT -10.365 -135.485 -10.035 -135.155 ;
        RECT -10.365 -136.845 -10.035 -136.515 ;
        RECT -10.365 -138.205 -10.035 -137.875 ;
        RECT -10.365 -139.565 -10.035 -139.235 ;
        RECT -10.365 -140.925 -10.035 -140.595 ;
        RECT -10.365 -142.285 -10.035 -141.955 ;
        RECT -10.365 -145.005 -10.035 -144.675 ;
        RECT -10.365 -146.365 -10.035 -146.035 ;
        RECT -10.365 -147.725 -10.035 -147.395 ;
        RECT -10.365 -149.085 -10.035 -148.755 ;
        RECT -10.365 -150.445 -10.035 -150.115 ;
        RECT -10.365 -151.805 -10.035 -151.475 ;
        RECT -10.365 -153.165 -10.035 -152.835 ;
        RECT -10.365 -154.525 -10.035 -154.195 ;
        RECT -10.365 -155.885 -10.035 -155.555 ;
        RECT -10.365 -157.245 -10.035 -156.915 ;
        RECT -10.365 -158.605 -10.035 -158.275 ;
        RECT -10.365 -159.965 -10.035 -159.635 ;
        RECT -10.365 -161.325 -10.035 -160.995 ;
        RECT -10.365 -162.685 -10.035 -162.355 ;
        RECT -10.365 -164.045 -10.035 -163.715 ;
        RECT -10.365 -165.405 -10.035 -165.075 ;
        RECT -10.365 -166.765 -10.035 -166.435 ;
        RECT -10.36 -166.765 -10.04 245.285 ;
        RECT -10.365 244.04 -10.035 245.17 ;
        RECT -10.365 239.875 -10.035 240.205 ;
        RECT -10.365 238.515 -10.035 238.845 ;
        RECT -10.365 237.155 -10.035 237.485 ;
        RECT -10.365 235.795 -10.035 236.125 ;
        RECT -10.365 234.435 -10.035 234.765 ;
        RECT -10.365 233.075 -10.035 233.405 ;
        RECT -10.365 231.715 -10.035 232.045 ;
        RECT -10.365 227.635 -10.035 227.965 ;
        RECT -10.365 224.915 -10.035 225.245 ;
        RECT -10.365 218.115 -10.035 218.445 ;
        RECT -10.365 216.755 -10.035 217.085 ;
        RECT -10.365 207.235 -10.035 207.565 ;
        RECT -10.365 204.515 -10.035 204.845 ;
        RECT -10.365 203.155 -10.035 203.485 ;
        RECT -10.365 199.075 -10.035 199.405 ;
        RECT -10.365 196.355 -10.035 196.685 ;
        RECT -10.365 189.555 -10.035 189.885 ;
        RECT -10.365 188.195 -10.035 188.525 ;
        RECT -10.365 185.475 -10.035 185.805 ;
        RECT -10.365 178.675 -10.035 179.005 ;
        RECT -10.365 175.955 -10.035 176.285 ;
        RECT -10.365 174.595 -10.035 174.925 ;
        RECT -10.365 167.795 -10.035 168.125 ;
        RECT -10.365 160.995 -10.035 161.325 ;
        RECT -10.365 159.635 -10.035 159.965 ;
        RECT -10.365 156.915 -10.035 157.245 ;
        RECT -10.365 150.115 -10.035 150.445 ;
        RECT -10.365 147.395 -10.035 147.725 ;
        RECT -10.365 146.035 -10.035 146.365 ;
        RECT -10.365 139.235 -10.035 139.565 ;
        RECT -10.365 136.515 -10.035 136.845 ;
        RECT -10.365 132.435 -10.035 132.765 ;
        RECT -10.365 131.075 -10.035 131.405 ;
        RECT -10.365 128.355 -10.035 128.685 ;
        RECT -10.365 118.835 -10.035 119.165 ;
        RECT -10.365 117.475 -10.035 117.805 ;
        RECT -10.365 110.675 -10.035 111.005 ;
        RECT -10.365 107.955 -10.035 108.285 ;
        RECT -10.365 103.875 -10.035 104.205 ;
        RECT -10.365 99.795 -10.035 100.125 ;
        RECT -10.365 97.075 -10.035 97.405 ;
        RECT -10.365 90.275 -10.035 90.605 ;
        RECT -10.365 88.915 -10.035 89.245 ;
        RECT -10.365 82.115 -10.035 82.445 ;
        RECT -10.365 79.395 -10.035 79.725 ;
        RECT -10.365 75.315 -10.035 75.645 ;
        RECT -10.365 71.235 -10.035 71.565 ;
        RECT -10.365 68.515 -10.035 68.845 ;
        RECT -10.365 61.715 -10.035 62.045 ;
        RECT -10.365 60.355 -10.035 60.685 ;
        RECT -10.365 50.835 -10.035 51.165 ;
    END
    PORT
      LAYER met3 ;
        RECT -21.245 -63.405 -20.915 -63.075 ;
        RECT -21.245 -64.765 -20.915 -64.435 ;
        RECT -21.245 -66.125 -20.915 -65.795 ;
        RECT -21.245 -67.485 -20.915 -67.155 ;
        RECT -21.245 -68.845 -20.915 -68.515 ;
        RECT -21.245 -70.205 -20.915 -69.875 ;
        RECT -21.245 -71.565 -20.915 -71.235 ;
        RECT -21.245 -72.925 -20.915 -72.595 ;
        RECT -21.245 -74.285 -20.915 -73.955 ;
        RECT -21.245 -75.645 -20.915 -75.315 ;
        RECT -21.245 -77.005 -20.915 -76.675 ;
        RECT -21.245 -78.365 -20.915 -78.035 ;
        RECT -21.245 -79.725 -20.915 -79.395 ;
        RECT -21.245 -81.085 -20.915 -80.755 ;
        RECT -21.245 -82.445 -20.915 -82.115 ;
        RECT -21.245 -83.805 -20.915 -83.475 ;
        RECT -21.245 -85.165 -20.915 -84.835 ;
        RECT -21.245 -86.525 -20.915 -86.195 ;
        RECT -21.24 -87.88 -20.92 -63.075 ;
    END
    PORT
      LAYER met3 ;
        RECT -21.245 -120.525 -20.915 -120.195 ;
        RECT -21.245 -123.245 -20.915 -122.915 ;
        RECT -21.245 -124.605 -20.915 -124.275 ;
        RECT -21.245 -125.965 -20.915 -125.635 ;
        RECT -21.245 -134.125 -20.915 -133.795 ;
        RECT -21.245 -136.845 -20.915 -136.515 ;
        RECT -21.245 -140.925 -20.915 -140.595 ;
        RECT -21.245 -143.645 -20.915 -143.315 ;
        RECT -21.245 -146.365 -20.915 -146.035 ;
        RECT -21.245 -147.725 -20.915 -147.395 ;
        RECT -21.245 -151.805 -20.915 -151.475 ;
        RECT -21.245 -155.885 -20.915 -155.555 ;
        RECT -21.245 -157.245 -20.915 -156.915 ;
        RECT -21.245 -158.605 -20.915 -158.275 ;
        RECT -21.245 -159.965 -20.915 -159.635 ;
        RECT -21.245 -161.325 -20.915 -160.995 ;
        RECT -21.245 -162.685 -20.915 -162.355 ;
        RECT -21.245 -164.045 -20.915 -163.715 ;
        RECT -21.245 -165.405 -20.915 -165.075 ;
        RECT -21.245 -166.765 -20.915 -166.435 ;
        RECT -21.245 -168.655 -20.915 -168.325 ;
        RECT -21.245 -169.485 -20.915 -169.155 ;
        RECT -21.245 -170.845 -20.915 -170.515 ;
        RECT -21.245 -172.205 -20.915 -171.875 ;
        RECT -21.24 -172.205 -20.92 -119.52 ;
    END
    PORT
      LAYER met3 ;
        RECT -19.885 244.04 -19.555 245.17 ;
        RECT -19.885 239.875 -19.555 240.205 ;
        RECT -19.885 238.515 -19.555 238.845 ;
        RECT -19.885 237.155 -19.555 237.485 ;
        RECT -19.885 235.795 -19.555 236.125 ;
        RECT -19.885 234.435 -19.555 234.765 ;
        RECT -19.885 233.075 -19.555 233.405 ;
        RECT -19.885 231.715 -19.555 232.045 ;
        RECT -19.885 230.355 -19.555 230.685 ;
        RECT -19.885 228.995 -19.555 229.325 ;
        RECT -19.885 227.635 -19.555 227.965 ;
        RECT -19.885 226.275 -19.555 226.605 ;
        RECT -19.885 224.915 -19.555 225.245 ;
        RECT -19.885 223.555 -19.555 223.885 ;
        RECT -19.885 222.195 -19.555 222.525 ;
        RECT -19.885 220.835 -19.555 221.165 ;
        RECT -19.885 219.475 -19.555 219.805 ;
        RECT -19.885 218.115 -19.555 218.445 ;
        RECT -19.885 216.755 -19.555 217.085 ;
        RECT -19.885 215.395 -19.555 215.725 ;
        RECT -19.885 214.035 -19.555 214.365 ;
        RECT -19.885 212.675 -19.555 213.005 ;
        RECT -19.885 211.315 -19.555 211.645 ;
        RECT -19.885 209.955 -19.555 210.285 ;
        RECT -19.885 208.595 -19.555 208.925 ;
        RECT -19.885 207.235 -19.555 207.565 ;
        RECT -19.885 205.875 -19.555 206.205 ;
        RECT -19.885 204.515 -19.555 204.845 ;
        RECT -19.885 203.155 -19.555 203.485 ;
        RECT -19.885 201.795 -19.555 202.125 ;
        RECT -19.885 200.435 -19.555 200.765 ;
        RECT -19.885 199.075 -19.555 199.405 ;
        RECT -19.885 197.715 -19.555 198.045 ;
        RECT -19.885 196.355 -19.555 196.685 ;
        RECT -19.885 194.995 -19.555 195.325 ;
        RECT -19.885 193.635 -19.555 193.965 ;
        RECT -19.885 192.275 -19.555 192.605 ;
        RECT -19.885 190.915 -19.555 191.245 ;
        RECT -19.885 189.555 -19.555 189.885 ;
        RECT -19.885 188.195 -19.555 188.525 ;
        RECT -19.885 186.835 -19.555 187.165 ;
        RECT -19.885 185.475 -19.555 185.805 ;
        RECT -19.885 184.115 -19.555 184.445 ;
        RECT -19.885 182.755 -19.555 183.085 ;
        RECT -19.885 181.395 -19.555 181.725 ;
        RECT -19.885 180.035 -19.555 180.365 ;
        RECT -19.885 178.675 -19.555 179.005 ;
        RECT -19.885 177.315 -19.555 177.645 ;
        RECT -19.885 175.955 -19.555 176.285 ;
        RECT -19.885 174.595 -19.555 174.925 ;
        RECT -19.885 173.235 -19.555 173.565 ;
        RECT -19.885 171.875 -19.555 172.205 ;
        RECT -19.885 170.515 -19.555 170.845 ;
        RECT -19.885 169.155 -19.555 169.485 ;
        RECT -19.885 167.795 -19.555 168.125 ;
        RECT -19.885 166.435 -19.555 166.765 ;
        RECT -19.885 165.075 -19.555 165.405 ;
        RECT -19.885 163.715 -19.555 164.045 ;
        RECT -19.885 162.355 -19.555 162.685 ;
        RECT -19.885 160.995 -19.555 161.325 ;
        RECT -19.885 159.635 -19.555 159.965 ;
        RECT -19.885 158.275 -19.555 158.605 ;
        RECT -19.885 156.915 -19.555 157.245 ;
        RECT -19.885 155.555 -19.555 155.885 ;
        RECT -19.885 154.195 -19.555 154.525 ;
        RECT -19.885 152.835 -19.555 153.165 ;
        RECT -19.885 151.475 -19.555 151.805 ;
        RECT -19.885 150.115 -19.555 150.445 ;
        RECT -19.885 148.755 -19.555 149.085 ;
        RECT -19.885 147.395 -19.555 147.725 ;
        RECT -19.885 146.035 -19.555 146.365 ;
        RECT -19.885 144.675 -19.555 145.005 ;
        RECT -19.885 143.315 -19.555 143.645 ;
        RECT -19.885 141.955 -19.555 142.285 ;
        RECT -19.885 140.595 -19.555 140.925 ;
        RECT -19.885 139.235 -19.555 139.565 ;
        RECT -19.885 137.875 -19.555 138.205 ;
        RECT -19.885 136.515 -19.555 136.845 ;
        RECT -19.885 135.155 -19.555 135.485 ;
        RECT -19.885 133.795 -19.555 134.125 ;
        RECT -19.885 132.435 -19.555 132.765 ;
        RECT -19.885 131.075 -19.555 131.405 ;
        RECT -19.885 129.715 -19.555 130.045 ;
        RECT -19.885 128.355 -19.555 128.685 ;
        RECT -19.885 126.995 -19.555 127.325 ;
        RECT -19.885 125.635 -19.555 125.965 ;
        RECT -19.885 124.275 -19.555 124.605 ;
        RECT -19.885 122.915 -19.555 123.245 ;
        RECT -19.885 121.555 -19.555 121.885 ;
        RECT -19.885 120.195 -19.555 120.525 ;
        RECT -19.885 118.835 -19.555 119.165 ;
        RECT -19.885 117.475 -19.555 117.805 ;
        RECT -19.885 116.115 -19.555 116.445 ;
        RECT -19.885 114.755 -19.555 115.085 ;
        RECT -19.885 113.395 -19.555 113.725 ;
        RECT -19.885 112.035 -19.555 112.365 ;
        RECT -19.885 110.675 -19.555 111.005 ;
        RECT -19.885 109.315 -19.555 109.645 ;
        RECT -19.885 107.955 -19.555 108.285 ;
        RECT -19.885 106.595 -19.555 106.925 ;
        RECT -19.885 105.235 -19.555 105.565 ;
        RECT -19.885 103.875 -19.555 104.205 ;
        RECT -19.885 102.515 -19.555 102.845 ;
        RECT -19.885 101.155 -19.555 101.485 ;
        RECT -19.885 99.795 -19.555 100.125 ;
        RECT -19.885 98.435 -19.555 98.765 ;
        RECT -19.885 97.075 -19.555 97.405 ;
        RECT -19.885 95.715 -19.555 96.045 ;
        RECT -19.885 94.355 -19.555 94.685 ;
        RECT -19.885 92.995 -19.555 93.325 ;
        RECT -19.885 91.635 -19.555 91.965 ;
        RECT -19.885 90.275 -19.555 90.605 ;
        RECT -19.885 88.915 -19.555 89.245 ;
        RECT -19.885 87.555 -19.555 87.885 ;
        RECT -19.885 86.195 -19.555 86.525 ;
        RECT -19.885 84.835 -19.555 85.165 ;
        RECT -19.885 83.475 -19.555 83.805 ;
        RECT -19.885 82.115 -19.555 82.445 ;
        RECT -19.885 80.755 -19.555 81.085 ;
        RECT -19.885 79.395 -19.555 79.725 ;
        RECT -19.885 78.035 -19.555 78.365 ;
        RECT -19.885 76.675 -19.555 77.005 ;
        RECT -19.885 75.315 -19.555 75.645 ;
        RECT -19.885 73.955 -19.555 74.285 ;
        RECT -19.885 72.595 -19.555 72.925 ;
        RECT -19.885 71.235 -19.555 71.565 ;
        RECT -19.885 69.875 -19.555 70.205 ;
        RECT -19.885 68.515 -19.555 68.845 ;
        RECT -19.885 67.155 -19.555 67.485 ;
        RECT -19.885 65.795 -19.555 66.125 ;
        RECT -19.885 64.435 -19.555 64.765 ;
        RECT -19.885 63.075 -19.555 63.405 ;
        RECT -19.885 61.715 -19.555 62.045 ;
        RECT -19.885 60.355 -19.555 60.685 ;
        RECT -19.885 58.995 -19.555 59.325 ;
        RECT -19.885 57.635 -19.555 57.965 ;
        RECT -19.885 56.275 -19.555 56.605 ;
        RECT -19.885 54.915 -19.555 55.245 ;
        RECT -19.885 53.555 -19.555 53.885 ;
        RECT -19.885 52.195 -19.555 52.525 ;
        RECT -19.885 50.835 -19.555 51.165 ;
        RECT -19.885 49.475 -19.555 49.805 ;
        RECT -19.885 48.115 -19.555 48.445 ;
        RECT -19.885 46.755 -19.555 47.085 ;
        RECT -19.885 45.395 -19.555 45.725 ;
        RECT -19.885 44.035 -19.555 44.365 ;
        RECT -19.885 42.675 -19.555 43.005 ;
        RECT -19.885 41.315 -19.555 41.645 ;
        RECT -19.885 39.955 -19.555 40.285 ;
        RECT -19.885 38.595 -19.555 38.925 ;
        RECT -19.885 37.235 -19.555 37.565 ;
        RECT -19.885 35.875 -19.555 36.205 ;
        RECT -19.885 34.515 -19.555 34.845 ;
        RECT -19.885 33.155 -19.555 33.485 ;
        RECT -19.885 31.795 -19.555 32.125 ;
        RECT -19.885 30.435 -19.555 30.765 ;
        RECT -19.885 29.075 -19.555 29.405 ;
        RECT -19.885 27.715 -19.555 28.045 ;
        RECT -19.885 26.355 -19.555 26.685 ;
        RECT -19.885 24.995 -19.555 25.325 ;
        RECT -19.885 23.635 -19.555 23.965 ;
        RECT -19.885 22.275 -19.555 22.605 ;
        RECT -19.885 20.915 -19.555 21.245 ;
        RECT -19.885 19.555 -19.555 19.885 ;
        RECT -19.885 18.195 -19.555 18.525 ;
        RECT -19.885 16.835 -19.555 17.165 ;
        RECT -19.885 15.475 -19.555 15.805 ;
        RECT -19.885 14.115 -19.555 14.445 ;
        RECT -19.885 12.755 -19.555 13.085 ;
        RECT -19.885 11.395 -19.555 11.725 ;
        RECT -19.885 10.035 -19.555 10.365 ;
        RECT -19.885 8.675 -19.555 9.005 ;
        RECT -19.885 7.315 -19.555 7.645 ;
        RECT -19.885 5.955 -19.555 6.285 ;
        RECT -19.885 4.595 -19.555 4.925 ;
        RECT -19.885 3.235 -19.555 3.565 ;
        RECT -19.885 1.875 -19.555 2.205 ;
        RECT -19.885 0.515 -19.555 0.845 ;
        RECT -19.885 -0.845 -19.555 -0.515 ;
        RECT -19.885 -2.205 -19.555 -1.875 ;
        RECT -19.885 -3.565 -19.555 -3.235 ;
        RECT -19.885 -7.645 -19.555 -7.315 ;
        RECT -19.885 -9.005 -19.555 -8.675 ;
        RECT -19.885 -10.73 -19.555 -10.4 ;
        RECT -19.885 -15.805 -19.555 -15.475 ;
        RECT -19.885 -16.77 -19.555 -16.44 ;
        RECT -19.885 -18.525 -19.555 -18.195 ;
        RECT -19.885 -21.245 -19.555 -20.915 ;
        RECT -19.88 -22.6 -19.56 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -19.885 -28.045 -19.555 -27.715 ;
        RECT -19.885 -29.405 -19.555 -29.075 ;
        RECT -19.885 -30.765 -19.555 -30.435 ;
        RECT -19.885 -32.125 -19.555 -31.795 ;
        RECT -19.885 -33.71 -19.555 -33.38 ;
        RECT -19.885 -34.845 -19.555 -34.515 ;
        RECT -19.885 -36.205 -19.555 -35.875 ;
        RECT -19.885 -38.925 -19.555 -38.595 ;
        RECT -19.885 -39.75 -19.555 -39.42 ;
        RECT -19.885 -41.645 -19.555 -41.315 ;
        RECT -19.885 -44.365 -19.555 -44.035 ;
        RECT -19.885 -49.805 -19.555 -49.475 ;
        RECT -19.885 -51.165 -19.555 -50.835 ;
        RECT -19.885 -52.525 -19.555 -52.195 ;
        RECT -19.885 -53.885 -19.555 -53.555 ;
        RECT -19.885 -55.245 -19.555 -54.915 ;
        RECT -19.885 -56.605 -19.555 -56.275 ;
        RECT -19.885 -57.965 -19.555 -57.635 ;
        RECT -19.885 -59.325 -19.555 -58.995 ;
        RECT -19.885 -60.685 -19.555 -60.355 ;
        RECT -19.885 -62.045 -19.555 -61.715 ;
        RECT -19.885 -63.405 -19.555 -63.075 ;
        RECT -19.885 -64.765 -19.555 -64.435 ;
        RECT -19.885 -66.125 -19.555 -65.795 ;
        RECT -19.885 -67.485 -19.555 -67.155 ;
        RECT -19.885 -68.845 -19.555 -68.515 ;
        RECT -19.885 -70.205 -19.555 -69.875 ;
        RECT -19.885 -71.565 -19.555 -71.235 ;
        RECT -19.885 -73.19 -19.555 -72.86 ;
        RECT -19.885 -74.285 -19.555 -73.955 ;
        RECT -19.885 -75.645 -19.555 -75.315 ;
        RECT -19.885 -78.365 -19.555 -78.035 ;
        RECT -19.885 -79.725 -19.555 -79.395 ;
        RECT -19.885 -80.73 -19.555 -80.4 ;
        RECT -19.885 -82.445 -19.555 -82.115 ;
        RECT -19.885 -83.805 -19.555 -83.475 ;
        RECT -19.885 -86.525 -19.555 -86.195 ;
        RECT -19.885 -89.245 -19.555 -88.915 ;
        RECT -19.885 -90.605 -19.555 -90.275 ;
        RECT -19.885 -91.965 -19.555 -91.635 ;
        RECT -19.885 -93.325 -19.555 -92.995 ;
        RECT -19.885 -94.685 -19.555 -94.355 ;
        RECT -19.885 -95.37 -19.555 -95.04 ;
        RECT -19.885 -97.405 -19.555 -97.075 ;
        RECT -19.885 -100.125 -19.555 -99.795 ;
        RECT -19.885 -101.485 -19.555 -101.155 ;
        RECT -19.885 -102.91 -19.555 -102.58 ;
        RECT -19.885 -104.205 -19.555 -103.875 ;
        RECT -19.885 -105.565 -19.555 -105.235 ;
        RECT -19.885 -108.285 -19.555 -107.955 ;
        RECT -19.885 -113.725 -19.555 -113.395 ;
        RECT -19.885 -115.085 -19.555 -114.755 ;
        RECT -19.885 -116.445 -19.555 -116.115 ;
        RECT -19.885 -120.525 -19.555 -120.195 ;
        RECT -19.885 -123.245 -19.555 -122.915 ;
        RECT -19.885 -124.605 -19.555 -124.275 ;
        RECT -19.885 -125.965 -19.555 -125.635 ;
        RECT -19.885 -134.125 -19.555 -133.795 ;
        RECT -19.885 -136.845 -19.555 -136.515 ;
        RECT -19.885 -140.925 -19.555 -140.595 ;
        RECT -19.885 -143.645 -19.555 -143.315 ;
        RECT -19.885 -146.365 -19.555 -146.035 ;
        RECT -19.885 -147.725 -19.555 -147.395 ;
        RECT -19.885 -151.805 -19.555 -151.475 ;
        RECT -19.885 -155.885 -19.555 -155.555 ;
        RECT -19.885 -157.245 -19.555 -156.915 ;
        RECT -19.885 -158.605 -19.555 -158.275 ;
        RECT -19.885 -159.965 -19.555 -159.635 ;
        RECT -19.885 -161.325 -19.555 -160.995 ;
        RECT -19.885 -162.685 -19.555 -162.355 ;
        RECT -19.885 -164.045 -19.555 -163.715 ;
        RECT -19.885 -165.405 -19.555 -165.075 ;
        RECT -19.885 -166.765 -19.555 -166.435 ;
        RECT -19.885 -168.655 -19.555 -168.325 ;
        RECT -19.885 -169.485 -19.555 -169.155 ;
        RECT -19.885 -170.845 -19.555 -170.515 ;
        RECT -19.885 -174.925 -19.555 -174.595 ;
        RECT -19.885 -177.645 -19.555 -177.315 ;
        RECT -19.885 -183.29 -19.555 -182.16 ;
        RECT -19.88 -183.405 -19.56 -27.715 ;
    END
    PORT
      LAYER met3 ;
        RECT -18.525 244.04 -18.195 245.17 ;
        RECT -18.525 239.875 -18.195 240.205 ;
        RECT -18.525 238.515 -18.195 238.845 ;
        RECT -18.525 237.155 -18.195 237.485 ;
        RECT -18.525 235.795 -18.195 236.125 ;
        RECT -18.525 234.435 -18.195 234.765 ;
        RECT -18.525 233.075 -18.195 233.405 ;
        RECT -18.525 231.715 -18.195 232.045 ;
        RECT -18.525 230.355 -18.195 230.685 ;
        RECT -18.525 228.995 -18.195 229.325 ;
        RECT -18.525 227.635 -18.195 227.965 ;
        RECT -18.525 226.275 -18.195 226.605 ;
        RECT -18.525 224.915 -18.195 225.245 ;
        RECT -18.525 223.555 -18.195 223.885 ;
        RECT -18.525 222.195 -18.195 222.525 ;
        RECT -18.525 220.835 -18.195 221.165 ;
        RECT -18.525 219.475 -18.195 219.805 ;
        RECT -18.525 218.115 -18.195 218.445 ;
        RECT -18.525 216.755 -18.195 217.085 ;
        RECT -18.525 215.395 -18.195 215.725 ;
        RECT -18.525 214.035 -18.195 214.365 ;
        RECT -18.525 212.675 -18.195 213.005 ;
        RECT -18.525 211.315 -18.195 211.645 ;
        RECT -18.525 209.955 -18.195 210.285 ;
        RECT -18.525 208.595 -18.195 208.925 ;
        RECT -18.525 207.235 -18.195 207.565 ;
        RECT -18.525 205.875 -18.195 206.205 ;
        RECT -18.525 204.515 -18.195 204.845 ;
        RECT -18.525 203.155 -18.195 203.485 ;
        RECT -18.525 201.795 -18.195 202.125 ;
        RECT -18.525 200.435 -18.195 200.765 ;
        RECT -18.525 199.075 -18.195 199.405 ;
        RECT -18.525 197.715 -18.195 198.045 ;
        RECT -18.525 196.355 -18.195 196.685 ;
        RECT -18.525 194.995 -18.195 195.325 ;
        RECT -18.525 193.635 -18.195 193.965 ;
        RECT -18.525 192.275 -18.195 192.605 ;
        RECT -18.525 190.915 -18.195 191.245 ;
        RECT -18.525 189.555 -18.195 189.885 ;
        RECT -18.525 188.195 -18.195 188.525 ;
        RECT -18.525 186.835 -18.195 187.165 ;
        RECT -18.525 185.475 -18.195 185.805 ;
        RECT -18.525 184.115 -18.195 184.445 ;
        RECT -18.525 182.755 -18.195 183.085 ;
        RECT -18.525 181.395 -18.195 181.725 ;
        RECT -18.525 180.035 -18.195 180.365 ;
        RECT -18.525 178.675 -18.195 179.005 ;
        RECT -18.525 177.315 -18.195 177.645 ;
        RECT -18.525 175.955 -18.195 176.285 ;
        RECT -18.525 174.595 -18.195 174.925 ;
        RECT -18.525 173.235 -18.195 173.565 ;
        RECT -18.525 171.875 -18.195 172.205 ;
        RECT -18.525 170.515 -18.195 170.845 ;
        RECT -18.525 169.155 -18.195 169.485 ;
        RECT -18.525 167.795 -18.195 168.125 ;
        RECT -18.525 166.435 -18.195 166.765 ;
        RECT -18.525 165.075 -18.195 165.405 ;
        RECT -18.525 163.715 -18.195 164.045 ;
        RECT -18.525 162.355 -18.195 162.685 ;
        RECT -18.525 160.995 -18.195 161.325 ;
        RECT -18.525 159.635 -18.195 159.965 ;
        RECT -18.525 158.275 -18.195 158.605 ;
        RECT -18.525 156.915 -18.195 157.245 ;
        RECT -18.525 155.555 -18.195 155.885 ;
        RECT -18.525 154.195 -18.195 154.525 ;
        RECT -18.525 152.835 -18.195 153.165 ;
        RECT -18.525 151.475 -18.195 151.805 ;
        RECT -18.525 150.115 -18.195 150.445 ;
        RECT -18.525 148.755 -18.195 149.085 ;
        RECT -18.525 147.395 -18.195 147.725 ;
        RECT -18.525 146.035 -18.195 146.365 ;
        RECT -18.525 144.675 -18.195 145.005 ;
        RECT -18.525 143.315 -18.195 143.645 ;
        RECT -18.525 141.955 -18.195 142.285 ;
        RECT -18.525 140.595 -18.195 140.925 ;
        RECT -18.525 139.235 -18.195 139.565 ;
        RECT -18.525 137.875 -18.195 138.205 ;
        RECT -18.525 136.515 -18.195 136.845 ;
        RECT -18.525 135.155 -18.195 135.485 ;
        RECT -18.525 133.795 -18.195 134.125 ;
        RECT -18.525 132.435 -18.195 132.765 ;
        RECT -18.525 131.075 -18.195 131.405 ;
        RECT -18.525 129.715 -18.195 130.045 ;
        RECT -18.525 128.355 -18.195 128.685 ;
        RECT -18.525 126.995 -18.195 127.325 ;
        RECT -18.525 125.635 -18.195 125.965 ;
        RECT -18.525 124.275 -18.195 124.605 ;
        RECT -18.525 122.915 -18.195 123.245 ;
        RECT -18.525 121.555 -18.195 121.885 ;
        RECT -18.525 120.195 -18.195 120.525 ;
        RECT -18.525 118.835 -18.195 119.165 ;
        RECT -18.525 117.475 -18.195 117.805 ;
        RECT -18.525 116.115 -18.195 116.445 ;
        RECT -18.525 114.755 -18.195 115.085 ;
        RECT -18.525 113.395 -18.195 113.725 ;
        RECT -18.525 112.035 -18.195 112.365 ;
        RECT -18.525 110.675 -18.195 111.005 ;
        RECT -18.525 109.315 -18.195 109.645 ;
        RECT -18.525 107.955 -18.195 108.285 ;
        RECT -18.525 106.595 -18.195 106.925 ;
        RECT -18.525 105.235 -18.195 105.565 ;
        RECT -18.525 103.875 -18.195 104.205 ;
        RECT -18.525 102.515 -18.195 102.845 ;
        RECT -18.525 101.155 -18.195 101.485 ;
        RECT -18.525 99.795 -18.195 100.125 ;
        RECT -18.525 98.435 -18.195 98.765 ;
        RECT -18.525 97.075 -18.195 97.405 ;
        RECT -18.525 95.715 -18.195 96.045 ;
        RECT -18.525 94.355 -18.195 94.685 ;
        RECT -18.525 92.995 -18.195 93.325 ;
        RECT -18.525 91.635 -18.195 91.965 ;
        RECT -18.525 90.275 -18.195 90.605 ;
        RECT -18.525 88.915 -18.195 89.245 ;
        RECT -18.525 87.555 -18.195 87.885 ;
        RECT -18.525 86.195 -18.195 86.525 ;
        RECT -18.525 84.835 -18.195 85.165 ;
        RECT -18.525 83.475 -18.195 83.805 ;
        RECT -18.525 82.115 -18.195 82.445 ;
        RECT -18.525 80.755 -18.195 81.085 ;
        RECT -18.525 79.395 -18.195 79.725 ;
        RECT -18.525 78.035 -18.195 78.365 ;
        RECT -18.525 76.675 -18.195 77.005 ;
        RECT -18.525 75.315 -18.195 75.645 ;
        RECT -18.525 73.955 -18.195 74.285 ;
        RECT -18.525 72.595 -18.195 72.925 ;
        RECT -18.525 71.235 -18.195 71.565 ;
        RECT -18.525 69.875 -18.195 70.205 ;
        RECT -18.525 68.515 -18.195 68.845 ;
        RECT -18.525 67.155 -18.195 67.485 ;
        RECT -18.525 65.795 -18.195 66.125 ;
        RECT -18.525 64.435 -18.195 64.765 ;
        RECT -18.525 63.075 -18.195 63.405 ;
        RECT -18.525 61.715 -18.195 62.045 ;
        RECT -18.525 60.355 -18.195 60.685 ;
        RECT -18.525 58.995 -18.195 59.325 ;
        RECT -18.525 57.635 -18.195 57.965 ;
        RECT -18.525 56.275 -18.195 56.605 ;
        RECT -18.525 54.915 -18.195 55.245 ;
        RECT -18.525 53.555 -18.195 53.885 ;
        RECT -18.525 52.195 -18.195 52.525 ;
        RECT -18.525 50.835 -18.195 51.165 ;
        RECT -18.525 49.475 -18.195 49.805 ;
        RECT -18.525 48.115 -18.195 48.445 ;
        RECT -18.525 46.755 -18.195 47.085 ;
        RECT -18.525 45.395 -18.195 45.725 ;
        RECT -18.525 44.035 -18.195 44.365 ;
        RECT -18.525 42.675 -18.195 43.005 ;
        RECT -18.525 41.315 -18.195 41.645 ;
        RECT -18.525 39.955 -18.195 40.285 ;
        RECT -18.525 38.595 -18.195 38.925 ;
        RECT -18.525 37.235 -18.195 37.565 ;
        RECT -18.525 35.875 -18.195 36.205 ;
        RECT -18.525 34.515 -18.195 34.845 ;
        RECT -18.525 33.155 -18.195 33.485 ;
        RECT -18.525 31.795 -18.195 32.125 ;
        RECT -18.525 30.435 -18.195 30.765 ;
        RECT -18.525 29.075 -18.195 29.405 ;
        RECT -18.525 27.715 -18.195 28.045 ;
        RECT -18.525 26.355 -18.195 26.685 ;
        RECT -18.525 24.995 -18.195 25.325 ;
        RECT -18.525 23.635 -18.195 23.965 ;
        RECT -18.525 22.275 -18.195 22.605 ;
        RECT -18.525 20.915 -18.195 21.245 ;
        RECT -18.525 19.555 -18.195 19.885 ;
        RECT -18.525 18.195 -18.195 18.525 ;
        RECT -18.525 16.835 -18.195 17.165 ;
        RECT -18.525 15.475 -18.195 15.805 ;
        RECT -18.525 14.115 -18.195 14.445 ;
        RECT -18.525 12.755 -18.195 13.085 ;
        RECT -18.525 11.395 -18.195 11.725 ;
        RECT -18.525 10.035 -18.195 10.365 ;
        RECT -18.525 8.675 -18.195 9.005 ;
        RECT -18.525 7.315 -18.195 7.645 ;
        RECT -18.525 5.955 -18.195 6.285 ;
        RECT -18.525 4.595 -18.195 4.925 ;
        RECT -18.525 3.235 -18.195 3.565 ;
        RECT -18.525 1.875 -18.195 2.205 ;
        RECT -18.525 0.515 -18.195 0.845 ;
        RECT -18.525 -0.845 -18.195 -0.515 ;
        RECT -18.525 -2.205 -18.195 -1.875 ;
        RECT -18.525 -3.565 -18.195 -3.235 ;
        RECT -18.525 -7.645 -18.195 -7.315 ;
        RECT -18.525 -9.005 -18.195 -8.675 ;
        RECT -18.525 -10.73 -18.195 -10.4 ;
        RECT -18.525 -15.805 -18.195 -15.475 ;
        RECT -18.525 -16.77 -18.195 -16.44 ;
        RECT -18.525 -18.525 -18.195 -18.195 ;
        RECT -18.525 -21.245 -18.195 -20.915 ;
        RECT -18.52 -21.245 -18.2 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -18.525 -26.685 -18.195 -26.355 ;
        RECT -18.525 -28.045 -18.195 -27.715 ;
        RECT -18.525 -29.405 -18.195 -29.075 ;
        RECT -18.525 -30.765 -18.195 -30.435 ;
        RECT -18.525 -32.125 -18.195 -31.795 ;
        RECT -18.525 -33.71 -18.195 -33.38 ;
        RECT -18.525 -34.845 -18.195 -34.515 ;
        RECT -18.525 -36.205 -18.195 -35.875 ;
        RECT -18.525 -38.925 -18.195 -38.595 ;
        RECT -18.525 -39.75 -18.195 -39.42 ;
        RECT -18.525 -41.645 -18.195 -41.315 ;
        RECT -18.525 -44.365 -18.195 -44.035 ;
        RECT -18.525 -49.805 -18.195 -49.475 ;
        RECT -18.525 -51.165 -18.195 -50.835 ;
        RECT -18.525 -52.525 -18.195 -52.195 ;
        RECT -18.525 -53.885 -18.195 -53.555 ;
        RECT -18.525 -55.245 -18.195 -54.915 ;
        RECT -18.525 -56.605 -18.195 -56.275 ;
        RECT -18.525 -57.965 -18.195 -57.635 ;
        RECT -18.525 -59.325 -18.195 -58.995 ;
        RECT -18.525 -60.685 -18.195 -60.355 ;
        RECT -18.525 -62.045 -18.195 -61.715 ;
        RECT -18.525 -63.405 -18.195 -63.075 ;
        RECT -18.525 -64.765 -18.195 -64.435 ;
        RECT -18.525 -66.125 -18.195 -65.795 ;
        RECT -18.525 -67.485 -18.195 -67.155 ;
        RECT -18.525 -68.845 -18.195 -68.515 ;
        RECT -18.525 -70.205 -18.195 -69.875 ;
        RECT -18.525 -71.565 -18.195 -71.235 ;
        RECT -18.525 -73.19 -18.195 -72.86 ;
        RECT -18.525 -74.285 -18.195 -73.955 ;
        RECT -18.525 -75.645 -18.195 -75.315 ;
        RECT -18.525 -78.365 -18.195 -78.035 ;
        RECT -18.525 -79.725 -18.195 -79.395 ;
        RECT -18.525 -80.73 -18.195 -80.4 ;
        RECT -18.525 -82.445 -18.195 -82.115 ;
        RECT -18.525 -83.805 -18.195 -83.475 ;
        RECT -18.525 -86.525 -18.195 -86.195 ;
        RECT -18.525 -89.245 -18.195 -88.915 ;
        RECT -18.525 -90.605 -18.195 -90.275 ;
        RECT -18.525 -91.965 -18.195 -91.635 ;
        RECT -18.525 -93.325 -18.195 -92.995 ;
        RECT -18.525 -94.685 -18.195 -94.355 ;
        RECT -18.525 -95.37 -18.195 -95.04 ;
        RECT -18.525 -97.405 -18.195 -97.075 ;
        RECT -18.525 -100.125 -18.195 -99.795 ;
        RECT -18.525 -101.485 -18.195 -101.155 ;
        RECT -18.525 -102.91 -18.195 -102.58 ;
        RECT -18.525 -104.205 -18.195 -103.875 ;
        RECT -18.525 -105.565 -18.195 -105.235 ;
        RECT -18.525 -108.285 -18.195 -107.955 ;
        RECT -18.52 -112.36 -18.2 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT -18.525 -174.925 -18.195 -174.595 ;
        RECT -18.525 -177.645 -18.195 -177.315 ;
        RECT -18.525 -183.29 -18.195 -182.16 ;
        RECT -18.52 -183.405 -18.2 -173.92 ;
    END
    PORT
      LAYER met3 ;
        RECT -17.165 244.04 -16.835 245.17 ;
        RECT -17.165 239.875 -16.835 240.205 ;
        RECT -17.165 238.515 -16.835 238.845 ;
        RECT -17.165 237.155 -16.835 237.485 ;
        RECT -17.165 235.795 -16.835 236.125 ;
        RECT -17.165 234.435 -16.835 234.765 ;
        RECT -17.165 233.075 -16.835 233.405 ;
        RECT -17.165 231.715 -16.835 232.045 ;
        RECT -17.165 230.355 -16.835 230.685 ;
        RECT -17.165 228.995 -16.835 229.325 ;
        RECT -17.165 227.635 -16.835 227.965 ;
        RECT -17.165 226.275 -16.835 226.605 ;
        RECT -17.165 224.915 -16.835 225.245 ;
        RECT -17.165 223.555 -16.835 223.885 ;
        RECT -17.165 222.195 -16.835 222.525 ;
        RECT -17.165 220.835 -16.835 221.165 ;
        RECT -17.165 219.475 -16.835 219.805 ;
        RECT -17.165 218.115 -16.835 218.445 ;
        RECT -17.165 216.755 -16.835 217.085 ;
        RECT -17.165 215.395 -16.835 215.725 ;
        RECT -17.165 214.035 -16.835 214.365 ;
        RECT -17.165 212.675 -16.835 213.005 ;
        RECT -17.165 211.315 -16.835 211.645 ;
        RECT -17.165 209.955 -16.835 210.285 ;
        RECT -17.165 208.595 -16.835 208.925 ;
        RECT -17.165 207.235 -16.835 207.565 ;
        RECT -17.165 205.875 -16.835 206.205 ;
        RECT -17.165 204.515 -16.835 204.845 ;
        RECT -17.165 203.155 -16.835 203.485 ;
        RECT -17.165 201.795 -16.835 202.125 ;
        RECT -17.165 200.435 -16.835 200.765 ;
        RECT -17.165 199.075 -16.835 199.405 ;
        RECT -17.165 197.715 -16.835 198.045 ;
        RECT -17.165 196.355 -16.835 196.685 ;
        RECT -17.165 194.995 -16.835 195.325 ;
        RECT -17.165 193.635 -16.835 193.965 ;
        RECT -17.165 192.275 -16.835 192.605 ;
        RECT -17.165 190.915 -16.835 191.245 ;
        RECT -17.165 189.555 -16.835 189.885 ;
        RECT -17.165 188.195 -16.835 188.525 ;
        RECT -17.165 186.835 -16.835 187.165 ;
        RECT -17.165 185.475 -16.835 185.805 ;
        RECT -17.165 184.115 -16.835 184.445 ;
        RECT -17.165 182.755 -16.835 183.085 ;
        RECT -17.165 181.395 -16.835 181.725 ;
        RECT -17.165 180.035 -16.835 180.365 ;
        RECT -17.165 178.675 -16.835 179.005 ;
        RECT -17.165 177.315 -16.835 177.645 ;
        RECT -17.165 175.955 -16.835 176.285 ;
        RECT -17.165 174.595 -16.835 174.925 ;
        RECT -17.165 173.235 -16.835 173.565 ;
        RECT -17.165 171.875 -16.835 172.205 ;
        RECT -17.165 170.515 -16.835 170.845 ;
        RECT -17.165 169.155 -16.835 169.485 ;
        RECT -17.165 167.795 -16.835 168.125 ;
        RECT -17.165 166.435 -16.835 166.765 ;
        RECT -17.165 165.075 -16.835 165.405 ;
        RECT -17.165 163.715 -16.835 164.045 ;
        RECT -17.165 162.355 -16.835 162.685 ;
        RECT -17.165 160.995 -16.835 161.325 ;
        RECT -17.165 159.635 -16.835 159.965 ;
        RECT -17.165 158.275 -16.835 158.605 ;
        RECT -17.165 156.915 -16.835 157.245 ;
        RECT -17.165 155.555 -16.835 155.885 ;
        RECT -17.165 154.195 -16.835 154.525 ;
        RECT -17.165 152.835 -16.835 153.165 ;
        RECT -17.165 151.475 -16.835 151.805 ;
        RECT -17.165 150.115 -16.835 150.445 ;
        RECT -17.165 148.755 -16.835 149.085 ;
        RECT -17.165 147.395 -16.835 147.725 ;
        RECT -17.165 146.035 -16.835 146.365 ;
        RECT -17.165 144.675 -16.835 145.005 ;
        RECT -17.165 143.315 -16.835 143.645 ;
        RECT -17.165 141.955 -16.835 142.285 ;
        RECT -17.165 140.595 -16.835 140.925 ;
        RECT -17.165 139.235 -16.835 139.565 ;
        RECT -17.165 137.875 -16.835 138.205 ;
        RECT -17.165 136.515 -16.835 136.845 ;
        RECT -17.165 135.155 -16.835 135.485 ;
        RECT -17.165 133.795 -16.835 134.125 ;
        RECT -17.165 132.435 -16.835 132.765 ;
        RECT -17.165 131.075 -16.835 131.405 ;
        RECT -17.165 129.715 -16.835 130.045 ;
        RECT -17.165 128.355 -16.835 128.685 ;
        RECT -17.165 126.995 -16.835 127.325 ;
        RECT -17.165 125.635 -16.835 125.965 ;
        RECT -17.165 124.275 -16.835 124.605 ;
        RECT -17.165 122.915 -16.835 123.245 ;
        RECT -17.165 121.555 -16.835 121.885 ;
        RECT -17.165 120.195 -16.835 120.525 ;
        RECT -17.165 118.835 -16.835 119.165 ;
        RECT -17.165 117.475 -16.835 117.805 ;
        RECT -17.165 116.115 -16.835 116.445 ;
        RECT -17.165 114.755 -16.835 115.085 ;
        RECT -17.165 113.395 -16.835 113.725 ;
        RECT -17.165 112.035 -16.835 112.365 ;
        RECT -17.165 110.675 -16.835 111.005 ;
        RECT -17.165 109.315 -16.835 109.645 ;
        RECT -17.165 107.955 -16.835 108.285 ;
        RECT -17.165 106.595 -16.835 106.925 ;
        RECT -17.165 105.235 -16.835 105.565 ;
        RECT -17.165 103.875 -16.835 104.205 ;
        RECT -17.165 102.515 -16.835 102.845 ;
        RECT -17.165 101.155 -16.835 101.485 ;
        RECT -17.165 99.795 -16.835 100.125 ;
        RECT -17.165 98.435 -16.835 98.765 ;
        RECT -17.165 97.075 -16.835 97.405 ;
        RECT -17.165 95.715 -16.835 96.045 ;
        RECT -17.165 94.355 -16.835 94.685 ;
        RECT -17.165 92.995 -16.835 93.325 ;
        RECT -17.165 91.635 -16.835 91.965 ;
        RECT -17.165 90.275 -16.835 90.605 ;
        RECT -17.165 88.915 -16.835 89.245 ;
        RECT -17.165 87.555 -16.835 87.885 ;
        RECT -17.165 86.195 -16.835 86.525 ;
        RECT -17.165 84.835 -16.835 85.165 ;
        RECT -17.165 83.475 -16.835 83.805 ;
        RECT -17.165 82.115 -16.835 82.445 ;
        RECT -17.165 80.755 -16.835 81.085 ;
        RECT -17.165 79.395 -16.835 79.725 ;
        RECT -17.165 78.035 -16.835 78.365 ;
        RECT -17.165 76.675 -16.835 77.005 ;
        RECT -17.165 75.315 -16.835 75.645 ;
        RECT -17.165 73.955 -16.835 74.285 ;
        RECT -17.165 72.595 -16.835 72.925 ;
        RECT -17.165 71.235 -16.835 71.565 ;
        RECT -17.165 69.875 -16.835 70.205 ;
        RECT -17.165 68.515 -16.835 68.845 ;
        RECT -17.165 67.155 -16.835 67.485 ;
        RECT -17.165 65.795 -16.835 66.125 ;
        RECT -17.165 64.435 -16.835 64.765 ;
        RECT -17.165 63.075 -16.835 63.405 ;
        RECT -17.165 61.715 -16.835 62.045 ;
        RECT -17.165 60.355 -16.835 60.685 ;
        RECT -17.165 58.995 -16.835 59.325 ;
        RECT -17.165 57.635 -16.835 57.965 ;
        RECT -17.165 56.275 -16.835 56.605 ;
        RECT -17.165 54.915 -16.835 55.245 ;
        RECT -17.165 53.555 -16.835 53.885 ;
        RECT -17.165 52.195 -16.835 52.525 ;
        RECT -17.165 50.835 -16.835 51.165 ;
        RECT -17.165 49.475 -16.835 49.805 ;
        RECT -17.165 48.115 -16.835 48.445 ;
        RECT -17.165 46.755 -16.835 47.085 ;
        RECT -17.165 45.395 -16.835 45.725 ;
        RECT -17.165 44.035 -16.835 44.365 ;
        RECT -17.165 42.675 -16.835 43.005 ;
        RECT -17.165 41.315 -16.835 41.645 ;
        RECT -17.165 39.955 -16.835 40.285 ;
        RECT -17.165 38.595 -16.835 38.925 ;
        RECT -17.165 37.235 -16.835 37.565 ;
        RECT -17.165 35.875 -16.835 36.205 ;
        RECT -17.165 34.515 -16.835 34.845 ;
        RECT -17.165 33.155 -16.835 33.485 ;
        RECT -17.165 31.795 -16.835 32.125 ;
        RECT -17.165 30.435 -16.835 30.765 ;
        RECT -17.165 29.075 -16.835 29.405 ;
        RECT -17.165 27.715 -16.835 28.045 ;
        RECT -17.165 26.355 -16.835 26.685 ;
        RECT -17.165 24.995 -16.835 25.325 ;
        RECT -17.165 23.635 -16.835 23.965 ;
        RECT -17.165 22.275 -16.835 22.605 ;
        RECT -17.165 20.915 -16.835 21.245 ;
        RECT -17.165 19.555 -16.835 19.885 ;
        RECT -17.165 18.195 -16.835 18.525 ;
        RECT -17.165 16.835 -16.835 17.165 ;
        RECT -17.165 15.475 -16.835 15.805 ;
        RECT -17.165 14.115 -16.835 14.445 ;
        RECT -17.165 12.755 -16.835 13.085 ;
        RECT -17.165 11.395 -16.835 11.725 ;
        RECT -17.165 10.035 -16.835 10.365 ;
        RECT -17.165 8.675 -16.835 9.005 ;
        RECT -17.165 7.315 -16.835 7.645 ;
        RECT -17.165 5.955 -16.835 6.285 ;
        RECT -17.165 4.595 -16.835 4.925 ;
        RECT -17.165 3.235 -16.835 3.565 ;
        RECT -17.165 1.875 -16.835 2.205 ;
        RECT -17.165 0.515 -16.835 0.845 ;
        RECT -17.165 -0.845 -16.835 -0.515 ;
        RECT -17.165 -2.205 -16.835 -1.875 ;
        RECT -17.165 -3.565 -16.835 -3.235 ;
        RECT -17.165 -4.925 -16.835 -4.595 ;
        RECT -17.165 -7.645 -16.835 -7.315 ;
        RECT -17.165 -9.005 -16.835 -8.675 ;
        RECT -17.165 -10.73 -16.835 -10.4 ;
        RECT -17.165 -11.725 -16.835 -11.395 ;
        RECT -17.16 -11.725 -16.84 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -17.165 -26.685 -16.835 -26.355 ;
        RECT -17.165 -28.045 -16.835 -27.715 ;
        RECT -17.165 -29.405 -16.835 -29.075 ;
        RECT -17.165 -30.765 -16.835 -30.435 ;
        RECT -17.165 -32.125 -16.835 -31.795 ;
        RECT -17.165 -33.71 -16.835 -33.38 ;
        RECT -17.165 -34.845 -16.835 -34.515 ;
        RECT -17.165 -36.205 -16.835 -35.875 ;
        RECT -17.165 -38.925 -16.835 -38.595 ;
        RECT -17.165 -39.75 -16.835 -39.42 ;
        RECT -17.165 -41.645 -16.835 -41.315 ;
        RECT -17.165 -44.365 -16.835 -44.035 ;
        RECT -17.165 -51.165 -16.835 -50.835 ;
        RECT -17.165 -52.525 -16.835 -52.195 ;
        RECT -17.165 -53.885 -16.835 -53.555 ;
        RECT -17.165 -55.245 -16.835 -54.915 ;
        RECT -17.165 -56.605 -16.835 -56.275 ;
        RECT -17.165 -57.965 -16.835 -57.635 ;
        RECT -17.165 -59.325 -16.835 -58.995 ;
        RECT -17.165 -60.685 -16.835 -60.355 ;
        RECT -17.165 -62.045 -16.835 -61.715 ;
        RECT -17.165 -63.405 -16.835 -63.075 ;
        RECT -17.165 -64.765 -16.835 -64.435 ;
        RECT -17.165 -66.125 -16.835 -65.795 ;
        RECT -17.165 -67.485 -16.835 -67.155 ;
        RECT -17.165 -68.845 -16.835 -68.515 ;
        RECT -17.165 -70.205 -16.835 -69.875 ;
        RECT -17.165 -71.565 -16.835 -71.235 ;
        RECT -17.165 -73.19 -16.835 -72.86 ;
        RECT -17.165 -74.285 -16.835 -73.955 ;
        RECT -17.165 -75.645 -16.835 -75.315 ;
        RECT -17.165 -78.365 -16.835 -78.035 ;
        RECT -17.165 -79.725 -16.835 -79.395 ;
        RECT -17.165 -80.73 -16.835 -80.4 ;
        RECT -17.165 -82.445 -16.835 -82.115 ;
        RECT -17.165 -83.805 -16.835 -83.475 ;
        RECT -17.165 -86.525 -16.835 -86.195 ;
        RECT -17.165 -89.245 -16.835 -88.915 ;
        RECT -17.165 -90.605 -16.835 -90.275 ;
        RECT -17.165 -91.965 -16.835 -91.635 ;
        RECT -17.165 -93.325 -16.835 -92.995 ;
        RECT -17.165 -94.685 -16.835 -94.355 ;
        RECT -17.165 -95.37 -16.835 -95.04 ;
        RECT -17.165 -97.405 -16.835 -97.075 ;
        RECT -17.165 -100.125 -16.835 -99.795 ;
        RECT -17.165 -102.91 -16.835 -102.58 ;
        RECT -17.165 -104.205 -16.835 -103.875 ;
        RECT -17.165 -105.565 -16.835 -105.235 ;
        RECT -17.165 -108.285 -16.835 -107.955 ;
        RECT -17.16 -113.04 -16.84 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT -17.165 -174.925 -16.835 -174.595 ;
        RECT -17.165 -177.645 -16.835 -177.315 ;
        RECT -17.165 -183.29 -16.835 -182.16 ;
        RECT -17.16 -183.405 -16.84 -172.56 ;
    END
    PORT
      LAYER met3 ;
        RECT -15.805 129.715 -15.475 130.045 ;
        RECT -15.805 128.355 -15.475 128.685 ;
        RECT -15.805 126.995 -15.475 127.325 ;
        RECT -15.805 125.635 -15.475 125.965 ;
        RECT -15.805 124.275 -15.475 124.605 ;
        RECT -15.805 122.915 -15.475 123.245 ;
        RECT -15.805 121.555 -15.475 121.885 ;
        RECT -15.805 120.195 -15.475 120.525 ;
        RECT -15.805 118.835 -15.475 119.165 ;
        RECT -15.805 117.475 -15.475 117.805 ;
        RECT -15.805 116.115 -15.475 116.445 ;
        RECT -15.805 114.755 -15.475 115.085 ;
        RECT -15.805 113.395 -15.475 113.725 ;
        RECT -15.805 112.035 -15.475 112.365 ;
        RECT -15.805 110.675 -15.475 111.005 ;
        RECT -15.805 109.315 -15.475 109.645 ;
        RECT -15.805 107.955 -15.475 108.285 ;
        RECT -15.805 106.595 -15.475 106.925 ;
        RECT -15.805 105.235 -15.475 105.565 ;
        RECT -15.805 103.875 -15.475 104.205 ;
        RECT -15.805 102.515 -15.475 102.845 ;
        RECT -15.805 101.155 -15.475 101.485 ;
        RECT -15.805 99.795 -15.475 100.125 ;
        RECT -15.805 98.435 -15.475 98.765 ;
        RECT -15.805 97.075 -15.475 97.405 ;
        RECT -15.805 95.715 -15.475 96.045 ;
        RECT -15.805 94.355 -15.475 94.685 ;
        RECT -15.805 92.995 -15.475 93.325 ;
        RECT -15.805 91.635 -15.475 91.965 ;
        RECT -15.805 90.275 -15.475 90.605 ;
        RECT -15.805 88.915 -15.475 89.245 ;
        RECT -15.805 87.555 -15.475 87.885 ;
        RECT -15.805 86.195 -15.475 86.525 ;
        RECT -15.805 84.835 -15.475 85.165 ;
        RECT -15.805 83.475 -15.475 83.805 ;
        RECT -15.805 82.115 -15.475 82.445 ;
        RECT -15.805 80.755 -15.475 81.085 ;
        RECT -15.805 79.395 -15.475 79.725 ;
        RECT -15.805 78.035 -15.475 78.365 ;
        RECT -15.805 76.675 -15.475 77.005 ;
        RECT -15.805 75.315 -15.475 75.645 ;
        RECT -15.805 73.955 -15.475 74.285 ;
        RECT -15.805 72.595 -15.475 72.925 ;
        RECT -15.805 71.235 -15.475 71.565 ;
        RECT -15.805 69.875 -15.475 70.205 ;
        RECT -15.805 68.515 -15.475 68.845 ;
        RECT -15.805 67.155 -15.475 67.485 ;
        RECT -15.805 65.795 -15.475 66.125 ;
        RECT -15.805 64.435 -15.475 64.765 ;
        RECT -15.805 63.075 -15.475 63.405 ;
        RECT -15.805 61.715 -15.475 62.045 ;
        RECT -15.805 60.355 -15.475 60.685 ;
        RECT -15.805 58.995 -15.475 59.325 ;
        RECT -15.805 57.635 -15.475 57.965 ;
        RECT -15.805 56.275 -15.475 56.605 ;
        RECT -15.805 54.915 -15.475 55.245 ;
        RECT -15.805 53.555 -15.475 53.885 ;
        RECT -15.805 52.195 -15.475 52.525 ;
        RECT -15.805 50.835 -15.475 51.165 ;
        RECT -15.805 49.475 -15.475 49.805 ;
        RECT -15.805 48.115 -15.475 48.445 ;
        RECT -15.805 46.755 -15.475 47.085 ;
        RECT -15.805 45.395 -15.475 45.725 ;
        RECT -15.805 44.035 -15.475 44.365 ;
        RECT -15.805 42.675 -15.475 43.005 ;
        RECT -15.805 41.315 -15.475 41.645 ;
        RECT -15.805 39.955 -15.475 40.285 ;
        RECT -15.805 38.595 -15.475 38.925 ;
        RECT -15.805 37.235 -15.475 37.565 ;
        RECT -15.805 35.875 -15.475 36.205 ;
        RECT -15.805 34.515 -15.475 34.845 ;
        RECT -15.805 33.155 -15.475 33.485 ;
        RECT -15.805 31.795 -15.475 32.125 ;
        RECT -15.805 30.435 -15.475 30.765 ;
        RECT -15.805 29.075 -15.475 29.405 ;
        RECT -15.805 27.715 -15.475 28.045 ;
        RECT -15.805 26.355 -15.475 26.685 ;
        RECT -15.805 24.995 -15.475 25.325 ;
        RECT -15.805 23.635 -15.475 23.965 ;
        RECT -15.805 22.275 -15.475 22.605 ;
        RECT -15.805 20.915 -15.475 21.245 ;
        RECT -15.805 19.555 -15.475 19.885 ;
        RECT -15.805 18.195 -15.475 18.525 ;
        RECT -15.805 16.835 -15.475 17.165 ;
        RECT -15.805 15.475 -15.475 15.805 ;
        RECT -15.805 14.115 -15.475 14.445 ;
        RECT -15.805 12.755 -15.475 13.085 ;
        RECT -15.805 11.395 -15.475 11.725 ;
        RECT -15.805 10.035 -15.475 10.365 ;
        RECT -15.805 8.675 -15.475 9.005 ;
        RECT -15.805 7.315 -15.475 7.645 ;
        RECT -15.805 5.955 -15.475 6.285 ;
        RECT -15.805 4.595 -15.475 4.925 ;
        RECT -15.805 3.235 -15.475 3.565 ;
        RECT -15.805 1.875 -15.475 2.205 ;
        RECT -15.805 0.515 -15.475 0.845 ;
        RECT -15.805 -0.845 -15.475 -0.515 ;
        RECT -15.805 -2.205 -15.475 -1.875 ;
        RECT -15.805 -3.565 -15.475 -3.235 ;
        RECT -15.805 -4.925 -15.475 -4.595 ;
        RECT -15.805 -7.645 -15.475 -7.315 ;
        RECT -15.805 -9.005 -15.475 -8.675 ;
        RECT -15.805 -10.73 -15.475 -10.4 ;
        RECT -15.805 -11.725 -15.475 -11.395 ;
        RECT -15.805 -13.085 -15.475 -12.755 ;
        RECT -15.805 -15.805 -15.475 -15.475 ;
        RECT -15.805 -16.77 -15.475 -16.44 ;
        RECT -15.805 -18.525 -15.475 -18.195 ;
        RECT -15.8 -19.88 -15.48 245.285 ;
        RECT -15.805 244.04 -15.475 245.17 ;
        RECT -15.805 239.875 -15.475 240.205 ;
        RECT -15.805 238.515 -15.475 238.845 ;
        RECT -15.805 237.155 -15.475 237.485 ;
        RECT -15.805 235.795 -15.475 236.125 ;
        RECT -15.805 234.435 -15.475 234.765 ;
        RECT -15.805 233.075 -15.475 233.405 ;
        RECT -15.805 231.715 -15.475 232.045 ;
        RECT -15.805 230.355 -15.475 230.685 ;
        RECT -15.805 228.995 -15.475 229.325 ;
        RECT -15.805 227.635 -15.475 227.965 ;
        RECT -15.805 226.275 -15.475 226.605 ;
        RECT -15.805 224.915 -15.475 225.245 ;
        RECT -15.805 223.555 -15.475 223.885 ;
        RECT -15.805 222.195 -15.475 222.525 ;
        RECT -15.805 220.835 -15.475 221.165 ;
        RECT -15.805 219.475 -15.475 219.805 ;
        RECT -15.805 218.115 -15.475 218.445 ;
        RECT -15.805 216.755 -15.475 217.085 ;
        RECT -15.805 215.395 -15.475 215.725 ;
        RECT -15.805 214.035 -15.475 214.365 ;
        RECT -15.805 212.675 -15.475 213.005 ;
        RECT -15.805 211.315 -15.475 211.645 ;
        RECT -15.805 209.955 -15.475 210.285 ;
        RECT -15.805 208.595 -15.475 208.925 ;
        RECT -15.805 207.235 -15.475 207.565 ;
        RECT -15.805 205.875 -15.475 206.205 ;
        RECT -15.805 204.515 -15.475 204.845 ;
        RECT -15.805 203.155 -15.475 203.485 ;
        RECT -15.805 201.795 -15.475 202.125 ;
        RECT -15.805 200.435 -15.475 200.765 ;
        RECT -15.805 199.075 -15.475 199.405 ;
        RECT -15.805 197.715 -15.475 198.045 ;
        RECT -15.805 196.355 -15.475 196.685 ;
        RECT -15.805 194.995 -15.475 195.325 ;
        RECT -15.805 193.635 -15.475 193.965 ;
        RECT -15.805 192.275 -15.475 192.605 ;
        RECT -15.805 190.915 -15.475 191.245 ;
        RECT -15.805 189.555 -15.475 189.885 ;
        RECT -15.805 188.195 -15.475 188.525 ;
        RECT -15.805 186.835 -15.475 187.165 ;
        RECT -15.805 185.475 -15.475 185.805 ;
        RECT -15.805 184.115 -15.475 184.445 ;
        RECT -15.805 182.755 -15.475 183.085 ;
        RECT -15.805 181.395 -15.475 181.725 ;
        RECT -15.805 180.035 -15.475 180.365 ;
        RECT -15.805 178.675 -15.475 179.005 ;
        RECT -15.805 177.315 -15.475 177.645 ;
        RECT -15.805 175.955 -15.475 176.285 ;
        RECT -15.805 174.595 -15.475 174.925 ;
        RECT -15.805 173.235 -15.475 173.565 ;
        RECT -15.805 171.875 -15.475 172.205 ;
        RECT -15.805 170.515 -15.475 170.845 ;
        RECT -15.805 169.155 -15.475 169.485 ;
        RECT -15.805 167.795 -15.475 168.125 ;
        RECT -15.805 166.435 -15.475 166.765 ;
        RECT -15.805 165.075 -15.475 165.405 ;
        RECT -15.805 163.715 -15.475 164.045 ;
        RECT -15.805 162.355 -15.475 162.685 ;
        RECT -15.805 160.995 -15.475 161.325 ;
        RECT -15.805 159.635 -15.475 159.965 ;
        RECT -15.805 158.275 -15.475 158.605 ;
        RECT -15.805 156.915 -15.475 157.245 ;
        RECT -15.805 155.555 -15.475 155.885 ;
        RECT -15.805 154.195 -15.475 154.525 ;
        RECT -15.805 152.835 -15.475 153.165 ;
        RECT -15.805 151.475 -15.475 151.805 ;
        RECT -15.805 150.115 -15.475 150.445 ;
        RECT -15.805 148.755 -15.475 149.085 ;
        RECT -15.805 147.395 -15.475 147.725 ;
        RECT -15.805 146.035 -15.475 146.365 ;
        RECT -15.805 144.675 -15.475 145.005 ;
        RECT -15.805 143.315 -15.475 143.645 ;
        RECT -15.805 141.955 -15.475 142.285 ;
        RECT -15.805 140.595 -15.475 140.925 ;
        RECT -15.805 139.235 -15.475 139.565 ;
        RECT -15.805 137.875 -15.475 138.205 ;
        RECT -15.805 136.515 -15.475 136.845 ;
        RECT -15.805 135.155 -15.475 135.485 ;
        RECT -15.805 133.795 -15.475 134.125 ;
        RECT -15.805 132.435 -15.475 132.765 ;
        RECT -15.805 131.075 -15.475 131.405 ;
    END
    PORT
      LAYER met3 ;
        RECT -25.325 244.04 -24.995 245.17 ;
        RECT -25.325 239.875 -24.995 240.205 ;
        RECT -25.325 238.515 -24.995 238.845 ;
        RECT -25.325 237.155 -24.995 237.485 ;
        RECT -25.325 235.795 -24.995 236.125 ;
        RECT -25.325 234.435 -24.995 234.765 ;
        RECT -25.325 233.075 -24.995 233.405 ;
        RECT -25.325 231.715 -24.995 232.045 ;
        RECT -25.325 230.355 -24.995 230.685 ;
        RECT -25.325 228.995 -24.995 229.325 ;
        RECT -25.325 227.635 -24.995 227.965 ;
        RECT -25.325 226.275 -24.995 226.605 ;
        RECT -25.325 224.915 -24.995 225.245 ;
        RECT -25.325 223.555 -24.995 223.885 ;
        RECT -25.325 222.195 -24.995 222.525 ;
        RECT -25.325 220.835 -24.995 221.165 ;
        RECT -25.325 219.475 -24.995 219.805 ;
        RECT -25.325 218.115 -24.995 218.445 ;
        RECT -25.325 216.755 -24.995 217.085 ;
        RECT -25.325 215.395 -24.995 215.725 ;
        RECT -25.325 214.035 -24.995 214.365 ;
        RECT -25.325 212.675 -24.995 213.005 ;
        RECT -25.325 211.315 -24.995 211.645 ;
        RECT -25.325 209.955 -24.995 210.285 ;
        RECT -25.325 208.595 -24.995 208.925 ;
        RECT -25.325 207.235 -24.995 207.565 ;
        RECT -25.325 205.875 -24.995 206.205 ;
        RECT -25.325 204.515 -24.995 204.845 ;
        RECT -25.325 203.155 -24.995 203.485 ;
        RECT -25.325 201.795 -24.995 202.125 ;
        RECT -25.325 200.435 -24.995 200.765 ;
        RECT -25.325 199.075 -24.995 199.405 ;
        RECT -25.325 197.715 -24.995 198.045 ;
        RECT -25.325 196.355 -24.995 196.685 ;
        RECT -25.325 194.995 -24.995 195.325 ;
        RECT -25.325 193.635 -24.995 193.965 ;
        RECT -25.325 192.275 -24.995 192.605 ;
        RECT -25.325 190.915 -24.995 191.245 ;
        RECT -25.325 189.555 -24.995 189.885 ;
        RECT -25.325 188.195 -24.995 188.525 ;
        RECT -25.325 186.835 -24.995 187.165 ;
        RECT -25.325 185.475 -24.995 185.805 ;
        RECT -25.325 184.115 -24.995 184.445 ;
        RECT -25.325 182.755 -24.995 183.085 ;
        RECT -25.325 181.395 -24.995 181.725 ;
        RECT -25.325 180.035 -24.995 180.365 ;
        RECT -25.325 178.675 -24.995 179.005 ;
        RECT -25.325 177.315 -24.995 177.645 ;
        RECT -25.325 175.955 -24.995 176.285 ;
        RECT -25.325 174.595 -24.995 174.925 ;
        RECT -25.325 173.235 -24.995 173.565 ;
        RECT -25.325 171.875 -24.995 172.205 ;
        RECT -25.325 170.515 -24.995 170.845 ;
        RECT -25.325 169.155 -24.995 169.485 ;
        RECT -25.325 167.795 -24.995 168.125 ;
        RECT -25.325 166.435 -24.995 166.765 ;
        RECT -25.325 165.075 -24.995 165.405 ;
        RECT -25.325 163.715 -24.995 164.045 ;
        RECT -25.325 162.355 -24.995 162.685 ;
        RECT -25.325 160.995 -24.995 161.325 ;
        RECT -25.325 159.635 -24.995 159.965 ;
        RECT -25.325 158.275 -24.995 158.605 ;
        RECT -25.325 156.915 -24.995 157.245 ;
        RECT -25.325 155.555 -24.995 155.885 ;
        RECT -25.325 154.195 -24.995 154.525 ;
        RECT -25.325 152.835 -24.995 153.165 ;
        RECT -25.325 151.475 -24.995 151.805 ;
        RECT -25.325 150.115 -24.995 150.445 ;
        RECT -25.325 148.755 -24.995 149.085 ;
        RECT -25.325 147.395 -24.995 147.725 ;
        RECT -25.325 146.035 -24.995 146.365 ;
        RECT -25.325 144.675 -24.995 145.005 ;
        RECT -25.325 143.315 -24.995 143.645 ;
        RECT -25.325 141.955 -24.995 142.285 ;
        RECT -25.325 140.595 -24.995 140.925 ;
        RECT -25.325 139.235 -24.995 139.565 ;
        RECT -25.325 137.875 -24.995 138.205 ;
        RECT -25.325 136.515 -24.995 136.845 ;
        RECT -25.325 135.155 -24.995 135.485 ;
        RECT -25.325 133.795 -24.995 134.125 ;
        RECT -25.325 132.435 -24.995 132.765 ;
        RECT -25.325 131.075 -24.995 131.405 ;
        RECT -25.325 129.715 -24.995 130.045 ;
        RECT -25.325 128.355 -24.995 128.685 ;
        RECT -25.325 126.995 -24.995 127.325 ;
        RECT -25.325 125.635 -24.995 125.965 ;
        RECT -25.325 124.275 -24.995 124.605 ;
        RECT -25.325 122.915 -24.995 123.245 ;
        RECT -25.325 121.555 -24.995 121.885 ;
        RECT -25.325 120.195 -24.995 120.525 ;
        RECT -25.325 118.835 -24.995 119.165 ;
        RECT -25.325 117.475 -24.995 117.805 ;
        RECT -25.325 116.115 -24.995 116.445 ;
        RECT -25.325 114.755 -24.995 115.085 ;
        RECT -25.325 113.395 -24.995 113.725 ;
        RECT -25.325 112.035 -24.995 112.365 ;
        RECT -25.325 110.675 -24.995 111.005 ;
        RECT -25.325 109.315 -24.995 109.645 ;
        RECT -25.325 107.955 -24.995 108.285 ;
        RECT -25.325 106.595 -24.995 106.925 ;
        RECT -25.325 105.235 -24.995 105.565 ;
        RECT -25.325 103.875 -24.995 104.205 ;
        RECT -25.325 102.515 -24.995 102.845 ;
        RECT -25.325 101.155 -24.995 101.485 ;
        RECT -25.325 99.795 -24.995 100.125 ;
        RECT -25.325 98.435 -24.995 98.765 ;
        RECT -25.325 97.075 -24.995 97.405 ;
        RECT -25.325 95.715 -24.995 96.045 ;
        RECT -25.325 94.355 -24.995 94.685 ;
        RECT -25.325 92.995 -24.995 93.325 ;
        RECT -25.325 91.635 -24.995 91.965 ;
        RECT -25.325 90.275 -24.995 90.605 ;
        RECT -25.325 88.915 -24.995 89.245 ;
        RECT -25.325 87.555 -24.995 87.885 ;
        RECT -25.325 86.195 -24.995 86.525 ;
        RECT -25.325 84.835 -24.995 85.165 ;
        RECT -25.325 83.475 -24.995 83.805 ;
        RECT -25.325 82.115 -24.995 82.445 ;
        RECT -25.325 80.755 -24.995 81.085 ;
        RECT -25.325 79.395 -24.995 79.725 ;
        RECT -25.325 78.035 -24.995 78.365 ;
        RECT -25.325 76.675 -24.995 77.005 ;
        RECT -25.325 75.315 -24.995 75.645 ;
        RECT -25.325 73.955 -24.995 74.285 ;
        RECT -25.325 72.595 -24.995 72.925 ;
        RECT -25.325 71.235 -24.995 71.565 ;
        RECT -25.325 69.875 -24.995 70.205 ;
        RECT -25.325 68.515 -24.995 68.845 ;
        RECT -25.325 67.155 -24.995 67.485 ;
        RECT -25.325 65.795 -24.995 66.125 ;
        RECT -25.325 64.435 -24.995 64.765 ;
        RECT -25.325 63.075 -24.995 63.405 ;
        RECT -25.325 61.715 -24.995 62.045 ;
        RECT -25.325 60.355 -24.995 60.685 ;
        RECT -25.325 58.995 -24.995 59.325 ;
        RECT -25.325 57.635 -24.995 57.965 ;
        RECT -25.325 56.275 -24.995 56.605 ;
        RECT -25.325 54.915 -24.995 55.245 ;
        RECT -25.325 53.555 -24.995 53.885 ;
        RECT -25.325 52.195 -24.995 52.525 ;
        RECT -25.325 50.835 -24.995 51.165 ;
        RECT -25.325 49.475 -24.995 49.805 ;
        RECT -25.325 48.115 -24.995 48.445 ;
        RECT -25.325 46.755 -24.995 47.085 ;
        RECT -25.325 45.395 -24.995 45.725 ;
        RECT -25.325 44.035 -24.995 44.365 ;
        RECT -25.325 42.675 -24.995 43.005 ;
        RECT -25.325 41.315 -24.995 41.645 ;
        RECT -25.325 39.955 -24.995 40.285 ;
        RECT -25.325 38.595 -24.995 38.925 ;
        RECT -25.325 37.235 -24.995 37.565 ;
        RECT -25.325 35.875 -24.995 36.205 ;
        RECT -25.325 34.515 -24.995 34.845 ;
        RECT -25.325 33.155 -24.995 33.485 ;
        RECT -25.325 31.795 -24.995 32.125 ;
        RECT -25.325 30.435 -24.995 30.765 ;
        RECT -25.325 29.075 -24.995 29.405 ;
        RECT -25.325 27.715 -24.995 28.045 ;
        RECT -25.325 26.355 -24.995 26.685 ;
        RECT -25.325 24.995 -24.995 25.325 ;
        RECT -25.325 23.635 -24.995 23.965 ;
        RECT -25.325 22.275 -24.995 22.605 ;
        RECT -25.325 20.915 -24.995 21.245 ;
        RECT -25.325 19.555 -24.995 19.885 ;
        RECT -25.325 18.195 -24.995 18.525 ;
        RECT -25.325 16.835 -24.995 17.165 ;
        RECT -25.325 15.475 -24.995 15.805 ;
        RECT -25.325 14.115 -24.995 14.445 ;
        RECT -25.325 12.755 -24.995 13.085 ;
        RECT -25.325 11.395 -24.995 11.725 ;
        RECT -25.325 10.035 -24.995 10.365 ;
        RECT -25.325 8.675 -24.995 9.005 ;
        RECT -25.325 7.315 -24.995 7.645 ;
        RECT -25.325 5.955 -24.995 6.285 ;
        RECT -25.325 4.595 -24.995 4.925 ;
        RECT -25.325 3.235 -24.995 3.565 ;
        RECT -25.325 1.875 -24.995 2.205 ;
        RECT -25.325 0.515 -24.995 0.845 ;
        RECT -25.325 -0.845 -24.995 -0.515 ;
        RECT -25.325 -2.205 -24.995 -1.875 ;
        RECT -25.325 -7.645 -24.995 -7.315 ;
        RECT -25.325 -9.005 -24.995 -8.675 ;
        RECT -25.325 -10.73 -24.995 -10.4 ;
        RECT -25.325 -15.805 -24.995 -15.475 ;
        RECT -25.325 -16.77 -24.995 -16.44 ;
        RECT -25.325 -18.525 -24.995 -18.195 ;
        RECT -25.325 -21.245 -24.995 -20.915 ;
        RECT -25.325 -29.405 -24.995 -29.075 ;
        RECT -25.325 -32.125 -24.995 -31.795 ;
        RECT -25.325 -33.71 -24.995 -33.38 ;
        RECT -25.325 -34.845 -24.995 -34.515 ;
        RECT -25.325 -36.205 -24.995 -35.875 ;
        RECT -25.325 -38.925 -24.995 -38.595 ;
        RECT -25.325 -39.75 -24.995 -39.42 ;
        RECT -25.325 -41.645 -24.995 -41.315 ;
        RECT -25.325 -44.365 -24.995 -44.035 ;
        RECT -25.325 -49.805 -24.995 -49.475 ;
        RECT -25.325 -51.165 -24.995 -50.835 ;
        RECT -25.325 -53.885 -24.995 -53.555 ;
        RECT -25.325 -55.245 -24.995 -54.915 ;
        RECT -25.325 -59.325 -24.995 -58.995 ;
        RECT -25.325 -60.685 -24.995 -60.355 ;
        RECT -25.325 -67.485 -24.995 -67.155 ;
        RECT -25.325 -68.845 -24.995 -68.515 ;
        RECT -25.325 -70.205 -24.995 -69.875 ;
        RECT -25.325 -71.565 -24.995 -71.235 ;
        RECT -25.325 -72.925 -24.995 -72.595 ;
        RECT -25.325 -74.285 -24.995 -73.955 ;
        RECT -25.325 -75.645 -24.995 -75.315 ;
        RECT -25.325 -77.005 -24.995 -76.675 ;
        RECT -25.325 -78.365 -24.995 -78.035 ;
        RECT -25.325 -79.725 -24.995 -79.395 ;
        RECT -25.325 -81.085 -24.995 -80.755 ;
        RECT -25.325 -82.445 -24.995 -82.115 ;
        RECT -25.325 -83.805 -24.995 -83.475 ;
        RECT -25.325 -85.165 -24.995 -84.835 ;
        RECT -25.325 -86.525 -24.995 -86.195 ;
        RECT -25.325 -87.885 -24.995 -87.555 ;
        RECT -25.325 -89.245 -24.995 -88.915 ;
        RECT -25.325 -90.605 -24.995 -90.275 ;
        RECT -25.325 -91.965 -24.995 -91.635 ;
        RECT -25.325 -93.325 -24.995 -92.995 ;
        RECT -25.325 -94.685 -24.995 -94.355 ;
        RECT -25.325 -96.045 -24.995 -95.715 ;
        RECT -25.325 -97.405 -24.995 -97.075 ;
        RECT -25.325 -98.765 -24.995 -98.435 ;
        RECT -25.325 -100.125 -24.995 -99.795 ;
        RECT -25.325 -101.485 -24.995 -101.155 ;
        RECT -25.325 -102.845 -24.995 -102.515 ;
        RECT -25.325 -104.205 -24.995 -103.875 ;
        RECT -25.325 -105.565 -24.995 -105.235 ;
        RECT -25.325 -106.925 -24.995 -106.595 ;
        RECT -25.325 -108.285 -24.995 -107.955 ;
        RECT -25.325 -109.645 -24.995 -109.315 ;
        RECT -25.325 -111.005 -24.995 -110.675 ;
        RECT -25.325 -112.365 -24.995 -112.035 ;
        RECT -25.325 -113.725 -24.995 -113.395 ;
        RECT -25.325 -115.085 -24.995 -114.755 ;
        RECT -25.325 -116.445 -24.995 -116.115 ;
        RECT -25.325 -117.805 -24.995 -117.475 ;
        RECT -25.325 -119.165 -24.995 -118.835 ;
        RECT -25.325 -120.525 -24.995 -120.195 ;
        RECT -25.325 -121.885 -24.995 -121.555 ;
        RECT -25.325 -123.245 -24.995 -122.915 ;
        RECT -25.325 -124.605 -24.995 -124.275 ;
        RECT -25.325 -125.965 -24.995 -125.635 ;
        RECT -25.325 -127.325 -24.995 -126.995 ;
        RECT -25.325 -128.685 -24.995 -128.355 ;
        RECT -25.325 -132.765 -24.995 -132.435 ;
        RECT -25.325 -134.125 -24.995 -133.795 ;
        RECT -25.325 -135.485 -24.995 -135.155 ;
        RECT -25.325 -136.845 -24.995 -136.515 ;
        RECT -25.325 -140.925 -24.995 -140.595 ;
        RECT -25.325 -142.285 -24.995 -141.955 ;
        RECT -25.325 -143.645 -24.995 -143.315 ;
        RECT -25.325 -145.005 -24.995 -144.675 ;
        RECT -25.325 -146.365 -24.995 -146.035 ;
        RECT -25.325 -147.725 -24.995 -147.395 ;
        RECT -25.325 -151.805 -24.995 -151.475 ;
        RECT -25.325 -155.885 -24.995 -155.555 ;
        RECT -25.325 -157.245 -24.995 -156.915 ;
        RECT -25.325 -158.605 -24.995 -158.275 ;
        RECT -25.325 -159.965 -24.995 -159.635 ;
        RECT -25.325 -161.325 -24.995 -160.995 ;
        RECT -25.325 -162.685 -24.995 -162.355 ;
        RECT -25.325 -164.045 -24.995 -163.715 ;
        RECT -25.325 -165.405 -24.995 -165.075 ;
        RECT -25.325 -166.765 -24.995 -166.435 ;
        RECT -25.325 -168.655 -24.995 -168.325 ;
        RECT -25.325 -169.485 -24.995 -169.155 ;
        RECT -25.325 -170.845 -24.995 -170.515 ;
        RECT -25.325 -172.205 -24.995 -171.875 ;
        RECT -25.325 -173.565 -24.995 -173.235 ;
        RECT -25.325 -174.925 -24.995 -174.595 ;
        RECT -25.325 -177.645 -24.995 -177.315 ;
        RECT -25.325 -183.29 -24.995 -182.16 ;
        RECT -25.32 -183.405 -25 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -23.965 244.04 -23.635 245.17 ;
        RECT -23.965 239.875 -23.635 240.205 ;
        RECT -23.965 238.515 -23.635 238.845 ;
        RECT -23.965 237.155 -23.635 237.485 ;
        RECT -23.965 235.795 -23.635 236.125 ;
        RECT -23.965 234.435 -23.635 234.765 ;
        RECT -23.965 233.075 -23.635 233.405 ;
        RECT -23.965 231.715 -23.635 232.045 ;
        RECT -23.965 230.355 -23.635 230.685 ;
        RECT -23.965 228.995 -23.635 229.325 ;
        RECT -23.965 227.635 -23.635 227.965 ;
        RECT -23.965 226.275 -23.635 226.605 ;
        RECT -23.965 224.915 -23.635 225.245 ;
        RECT -23.965 223.555 -23.635 223.885 ;
        RECT -23.965 222.195 -23.635 222.525 ;
        RECT -23.965 220.835 -23.635 221.165 ;
        RECT -23.965 219.475 -23.635 219.805 ;
        RECT -23.965 218.115 -23.635 218.445 ;
        RECT -23.965 216.755 -23.635 217.085 ;
        RECT -23.965 215.395 -23.635 215.725 ;
        RECT -23.965 214.035 -23.635 214.365 ;
        RECT -23.965 212.675 -23.635 213.005 ;
        RECT -23.965 211.315 -23.635 211.645 ;
        RECT -23.965 209.955 -23.635 210.285 ;
        RECT -23.965 208.595 -23.635 208.925 ;
        RECT -23.965 207.235 -23.635 207.565 ;
        RECT -23.965 205.875 -23.635 206.205 ;
        RECT -23.965 204.515 -23.635 204.845 ;
        RECT -23.965 203.155 -23.635 203.485 ;
        RECT -23.965 201.795 -23.635 202.125 ;
        RECT -23.965 200.435 -23.635 200.765 ;
        RECT -23.965 199.075 -23.635 199.405 ;
        RECT -23.965 197.715 -23.635 198.045 ;
        RECT -23.965 196.355 -23.635 196.685 ;
        RECT -23.965 194.995 -23.635 195.325 ;
        RECT -23.965 193.635 -23.635 193.965 ;
        RECT -23.965 192.275 -23.635 192.605 ;
        RECT -23.965 190.915 -23.635 191.245 ;
        RECT -23.965 189.555 -23.635 189.885 ;
        RECT -23.965 188.195 -23.635 188.525 ;
        RECT -23.965 186.835 -23.635 187.165 ;
        RECT -23.965 185.475 -23.635 185.805 ;
        RECT -23.965 184.115 -23.635 184.445 ;
        RECT -23.965 182.755 -23.635 183.085 ;
        RECT -23.965 181.395 -23.635 181.725 ;
        RECT -23.965 180.035 -23.635 180.365 ;
        RECT -23.965 178.675 -23.635 179.005 ;
        RECT -23.965 177.315 -23.635 177.645 ;
        RECT -23.965 175.955 -23.635 176.285 ;
        RECT -23.965 174.595 -23.635 174.925 ;
        RECT -23.965 173.235 -23.635 173.565 ;
        RECT -23.965 171.875 -23.635 172.205 ;
        RECT -23.965 170.515 -23.635 170.845 ;
        RECT -23.965 169.155 -23.635 169.485 ;
        RECT -23.965 167.795 -23.635 168.125 ;
        RECT -23.965 166.435 -23.635 166.765 ;
        RECT -23.965 165.075 -23.635 165.405 ;
        RECT -23.965 163.715 -23.635 164.045 ;
        RECT -23.965 162.355 -23.635 162.685 ;
        RECT -23.965 160.995 -23.635 161.325 ;
        RECT -23.965 159.635 -23.635 159.965 ;
        RECT -23.965 158.275 -23.635 158.605 ;
        RECT -23.965 156.915 -23.635 157.245 ;
        RECT -23.965 155.555 -23.635 155.885 ;
        RECT -23.965 154.195 -23.635 154.525 ;
        RECT -23.965 152.835 -23.635 153.165 ;
        RECT -23.965 151.475 -23.635 151.805 ;
        RECT -23.965 150.115 -23.635 150.445 ;
        RECT -23.965 148.755 -23.635 149.085 ;
        RECT -23.965 147.395 -23.635 147.725 ;
        RECT -23.965 146.035 -23.635 146.365 ;
        RECT -23.965 144.675 -23.635 145.005 ;
        RECT -23.965 143.315 -23.635 143.645 ;
        RECT -23.965 141.955 -23.635 142.285 ;
        RECT -23.965 140.595 -23.635 140.925 ;
        RECT -23.965 139.235 -23.635 139.565 ;
        RECT -23.965 137.875 -23.635 138.205 ;
        RECT -23.965 136.515 -23.635 136.845 ;
        RECT -23.965 135.155 -23.635 135.485 ;
        RECT -23.965 133.795 -23.635 134.125 ;
        RECT -23.965 132.435 -23.635 132.765 ;
        RECT -23.965 131.075 -23.635 131.405 ;
        RECT -23.965 129.715 -23.635 130.045 ;
        RECT -23.965 128.355 -23.635 128.685 ;
        RECT -23.965 126.995 -23.635 127.325 ;
        RECT -23.965 125.635 -23.635 125.965 ;
        RECT -23.965 124.275 -23.635 124.605 ;
        RECT -23.965 122.915 -23.635 123.245 ;
        RECT -23.965 121.555 -23.635 121.885 ;
        RECT -23.965 120.195 -23.635 120.525 ;
        RECT -23.965 118.835 -23.635 119.165 ;
        RECT -23.965 117.475 -23.635 117.805 ;
        RECT -23.965 116.115 -23.635 116.445 ;
        RECT -23.965 114.755 -23.635 115.085 ;
        RECT -23.965 113.395 -23.635 113.725 ;
        RECT -23.965 112.035 -23.635 112.365 ;
        RECT -23.965 110.675 -23.635 111.005 ;
        RECT -23.965 109.315 -23.635 109.645 ;
        RECT -23.965 107.955 -23.635 108.285 ;
        RECT -23.965 106.595 -23.635 106.925 ;
        RECT -23.965 105.235 -23.635 105.565 ;
        RECT -23.965 103.875 -23.635 104.205 ;
        RECT -23.965 102.515 -23.635 102.845 ;
        RECT -23.965 101.155 -23.635 101.485 ;
        RECT -23.965 99.795 -23.635 100.125 ;
        RECT -23.965 98.435 -23.635 98.765 ;
        RECT -23.965 97.075 -23.635 97.405 ;
        RECT -23.965 95.715 -23.635 96.045 ;
        RECT -23.965 94.355 -23.635 94.685 ;
        RECT -23.965 92.995 -23.635 93.325 ;
        RECT -23.965 91.635 -23.635 91.965 ;
        RECT -23.965 90.275 -23.635 90.605 ;
        RECT -23.965 88.915 -23.635 89.245 ;
        RECT -23.965 87.555 -23.635 87.885 ;
        RECT -23.965 86.195 -23.635 86.525 ;
        RECT -23.965 84.835 -23.635 85.165 ;
        RECT -23.965 83.475 -23.635 83.805 ;
        RECT -23.965 82.115 -23.635 82.445 ;
        RECT -23.965 80.755 -23.635 81.085 ;
        RECT -23.965 79.395 -23.635 79.725 ;
        RECT -23.965 78.035 -23.635 78.365 ;
        RECT -23.965 76.675 -23.635 77.005 ;
        RECT -23.965 75.315 -23.635 75.645 ;
        RECT -23.965 73.955 -23.635 74.285 ;
        RECT -23.965 72.595 -23.635 72.925 ;
        RECT -23.965 71.235 -23.635 71.565 ;
        RECT -23.965 69.875 -23.635 70.205 ;
        RECT -23.965 68.515 -23.635 68.845 ;
        RECT -23.965 67.155 -23.635 67.485 ;
        RECT -23.965 65.795 -23.635 66.125 ;
        RECT -23.965 64.435 -23.635 64.765 ;
        RECT -23.965 63.075 -23.635 63.405 ;
        RECT -23.965 61.715 -23.635 62.045 ;
        RECT -23.965 60.355 -23.635 60.685 ;
        RECT -23.965 58.995 -23.635 59.325 ;
        RECT -23.965 57.635 -23.635 57.965 ;
        RECT -23.965 56.275 -23.635 56.605 ;
        RECT -23.965 54.915 -23.635 55.245 ;
        RECT -23.965 53.555 -23.635 53.885 ;
        RECT -23.965 52.195 -23.635 52.525 ;
        RECT -23.965 50.835 -23.635 51.165 ;
        RECT -23.965 49.475 -23.635 49.805 ;
        RECT -23.965 48.115 -23.635 48.445 ;
        RECT -23.965 46.755 -23.635 47.085 ;
        RECT -23.965 45.395 -23.635 45.725 ;
        RECT -23.965 44.035 -23.635 44.365 ;
        RECT -23.965 42.675 -23.635 43.005 ;
        RECT -23.965 41.315 -23.635 41.645 ;
        RECT -23.965 39.955 -23.635 40.285 ;
        RECT -23.965 38.595 -23.635 38.925 ;
        RECT -23.965 37.235 -23.635 37.565 ;
        RECT -23.965 35.875 -23.635 36.205 ;
        RECT -23.965 34.515 -23.635 34.845 ;
        RECT -23.965 33.155 -23.635 33.485 ;
        RECT -23.965 31.795 -23.635 32.125 ;
        RECT -23.965 30.435 -23.635 30.765 ;
        RECT -23.965 29.075 -23.635 29.405 ;
        RECT -23.965 27.715 -23.635 28.045 ;
        RECT -23.965 26.355 -23.635 26.685 ;
        RECT -23.965 24.995 -23.635 25.325 ;
        RECT -23.965 23.635 -23.635 23.965 ;
        RECT -23.965 22.275 -23.635 22.605 ;
        RECT -23.965 20.915 -23.635 21.245 ;
        RECT -23.965 19.555 -23.635 19.885 ;
        RECT -23.965 18.195 -23.635 18.525 ;
        RECT -23.965 16.835 -23.635 17.165 ;
        RECT -23.965 15.475 -23.635 15.805 ;
        RECT -23.965 14.115 -23.635 14.445 ;
        RECT -23.965 12.755 -23.635 13.085 ;
        RECT -23.965 11.395 -23.635 11.725 ;
        RECT -23.965 10.035 -23.635 10.365 ;
        RECT -23.965 8.675 -23.635 9.005 ;
        RECT -23.965 7.315 -23.635 7.645 ;
        RECT -23.965 5.955 -23.635 6.285 ;
        RECT -23.965 4.595 -23.635 4.925 ;
        RECT -23.965 3.235 -23.635 3.565 ;
        RECT -23.965 1.875 -23.635 2.205 ;
        RECT -23.965 0.515 -23.635 0.845 ;
        RECT -23.965 -0.845 -23.635 -0.515 ;
        RECT -23.965 -2.205 -23.635 -1.875 ;
        RECT -23.965 -7.645 -23.635 -7.315 ;
        RECT -23.965 -9.005 -23.635 -8.675 ;
        RECT -23.965 -10.73 -23.635 -10.4 ;
        RECT -23.965 -15.805 -23.635 -15.475 ;
        RECT -23.965 -16.77 -23.635 -16.44 ;
        RECT -23.965 -18.525 -23.635 -18.195 ;
        RECT -23.965 -21.245 -23.635 -20.915 ;
        RECT -23.965 -29.405 -23.635 -29.075 ;
        RECT -23.965 -32.125 -23.635 -31.795 ;
        RECT -23.965 -33.71 -23.635 -33.38 ;
        RECT -23.965 -34.845 -23.635 -34.515 ;
        RECT -23.965 -36.205 -23.635 -35.875 ;
        RECT -23.965 -38.925 -23.635 -38.595 ;
        RECT -23.965 -39.75 -23.635 -39.42 ;
        RECT -23.965 -41.645 -23.635 -41.315 ;
        RECT -23.965 -44.365 -23.635 -44.035 ;
        RECT -23.965 -49.805 -23.635 -49.475 ;
        RECT -23.965 -51.165 -23.635 -50.835 ;
        RECT -23.965 -52.525 -23.635 -52.195 ;
        RECT -23.965 -53.885 -23.635 -53.555 ;
        RECT -23.965 -55.245 -23.635 -54.915 ;
        RECT -23.965 -56.605 -23.635 -56.275 ;
        RECT -23.965 -57.965 -23.635 -57.635 ;
        RECT -23.965 -59.325 -23.635 -58.995 ;
        RECT -23.965 -60.685 -23.635 -60.355 ;
        RECT -23.965 -62.045 -23.635 -61.715 ;
        RECT -23.965 -64.765 -23.635 -64.435 ;
        RECT -23.965 -66.125 -23.635 -65.795 ;
        RECT -23.965 -67.485 -23.635 -67.155 ;
        RECT -23.965 -68.845 -23.635 -68.515 ;
        RECT -23.965 -70.205 -23.635 -69.875 ;
        RECT -23.965 -71.565 -23.635 -71.235 ;
        RECT -23.965 -72.925 -23.635 -72.595 ;
        RECT -23.965 -74.285 -23.635 -73.955 ;
        RECT -23.965 -75.645 -23.635 -75.315 ;
        RECT -23.965 -77.005 -23.635 -76.675 ;
        RECT -23.965 -78.365 -23.635 -78.035 ;
        RECT -23.965 -79.725 -23.635 -79.395 ;
        RECT -23.965 -81.085 -23.635 -80.755 ;
        RECT -23.965 -82.445 -23.635 -82.115 ;
        RECT -23.965 -83.805 -23.635 -83.475 ;
        RECT -23.965 -85.165 -23.635 -84.835 ;
        RECT -23.965 -86.525 -23.635 -86.195 ;
        RECT -23.965 -87.885 -23.635 -87.555 ;
        RECT -23.965 -89.245 -23.635 -88.915 ;
        RECT -23.965 -90.605 -23.635 -90.275 ;
        RECT -23.965 -91.965 -23.635 -91.635 ;
        RECT -23.965 -93.325 -23.635 -92.995 ;
        RECT -23.965 -94.685 -23.635 -94.355 ;
        RECT -23.965 -96.045 -23.635 -95.715 ;
        RECT -23.965 -97.405 -23.635 -97.075 ;
        RECT -23.965 -98.765 -23.635 -98.435 ;
        RECT -23.965 -100.125 -23.635 -99.795 ;
        RECT -23.965 -101.485 -23.635 -101.155 ;
        RECT -23.965 -102.845 -23.635 -102.515 ;
        RECT -23.965 -104.205 -23.635 -103.875 ;
        RECT -23.965 -105.565 -23.635 -105.235 ;
        RECT -23.965 -106.925 -23.635 -106.595 ;
        RECT -23.965 -108.285 -23.635 -107.955 ;
        RECT -23.965 -109.645 -23.635 -109.315 ;
        RECT -23.965 -111.005 -23.635 -110.675 ;
        RECT -23.965 -112.365 -23.635 -112.035 ;
        RECT -23.965 -113.725 -23.635 -113.395 ;
        RECT -23.965 -115.085 -23.635 -114.755 ;
        RECT -23.965 -116.445 -23.635 -116.115 ;
        RECT -23.965 -117.805 -23.635 -117.475 ;
        RECT -23.965 -119.165 -23.635 -118.835 ;
        RECT -23.965 -120.525 -23.635 -120.195 ;
        RECT -23.965 -121.885 -23.635 -121.555 ;
        RECT -23.965 -123.245 -23.635 -122.915 ;
        RECT -23.965 -124.605 -23.635 -124.275 ;
        RECT -23.965 -125.965 -23.635 -125.635 ;
        RECT -23.965 -127.325 -23.635 -126.995 ;
        RECT -23.965 -134.125 -23.635 -133.795 ;
        RECT -23.965 -135.485 -23.635 -135.155 ;
        RECT -23.965 -136.845 -23.635 -136.515 ;
        RECT -23.965 -140.925 -23.635 -140.595 ;
        RECT -23.965 -142.285 -23.635 -141.955 ;
        RECT -23.965 -146.365 -23.635 -146.035 ;
        RECT -23.965 -147.725 -23.635 -147.395 ;
        RECT -23.965 -151.805 -23.635 -151.475 ;
        RECT -23.965 -157.245 -23.635 -156.915 ;
        RECT -23.965 -158.605 -23.635 -158.275 ;
        RECT -23.965 -159.965 -23.635 -159.635 ;
        RECT -23.965 -161.325 -23.635 -160.995 ;
        RECT -23.965 -162.685 -23.635 -162.355 ;
        RECT -23.965 -164.045 -23.635 -163.715 ;
        RECT -23.965 -165.405 -23.635 -165.075 ;
        RECT -23.965 -166.765 -23.635 -166.435 ;
        RECT -23.965 -168.655 -23.635 -168.325 ;
        RECT -23.965 -169.485 -23.635 -169.155 ;
        RECT -23.965 -170.845 -23.635 -170.515 ;
        RECT -23.965 -172.205 -23.635 -171.875 ;
        RECT -23.965 -174.925 -23.635 -174.595 ;
        RECT -23.965 -177.645 -23.635 -177.315 ;
        RECT -23.965 -183.29 -23.635 -182.16 ;
        RECT -23.96 -183.405 -23.64 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -22.605 244.04 -22.275 245.17 ;
        RECT -22.605 239.875 -22.275 240.205 ;
        RECT -22.605 238.515 -22.275 238.845 ;
        RECT -22.605 237.155 -22.275 237.485 ;
        RECT -22.605 235.795 -22.275 236.125 ;
        RECT -22.605 234.435 -22.275 234.765 ;
        RECT -22.605 233.075 -22.275 233.405 ;
        RECT -22.605 231.715 -22.275 232.045 ;
        RECT -22.605 230.355 -22.275 230.685 ;
        RECT -22.605 228.995 -22.275 229.325 ;
        RECT -22.605 227.635 -22.275 227.965 ;
        RECT -22.605 226.275 -22.275 226.605 ;
        RECT -22.605 224.915 -22.275 225.245 ;
        RECT -22.605 223.555 -22.275 223.885 ;
        RECT -22.605 222.195 -22.275 222.525 ;
        RECT -22.605 220.835 -22.275 221.165 ;
        RECT -22.605 219.475 -22.275 219.805 ;
        RECT -22.605 218.115 -22.275 218.445 ;
        RECT -22.605 216.755 -22.275 217.085 ;
        RECT -22.605 215.395 -22.275 215.725 ;
        RECT -22.605 214.035 -22.275 214.365 ;
        RECT -22.605 212.675 -22.275 213.005 ;
        RECT -22.605 211.315 -22.275 211.645 ;
        RECT -22.605 209.955 -22.275 210.285 ;
        RECT -22.605 208.595 -22.275 208.925 ;
        RECT -22.605 207.235 -22.275 207.565 ;
        RECT -22.605 205.875 -22.275 206.205 ;
        RECT -22.605 204.515 -22.275 204.845 ;
        RECT -22.605 203.155 -22.275 203.485 ;
        RECT -22.605 201.795 -22.275 202.125 ;
        RECT -22.605 200.435 -22.275 200.765 ;
        RECT -22.605 199.075 -22.275 199.405 ;
        RECT -22.605 197.715 -22.275 198.045 ;
        RECT -22.605 196.355 -22.275 196.685 ;
        RECT -22.605 194.995 -22.275 195.325 ;
        RECT -22.605 193.635 -22.275 193.965 ;
        RECT -22.605 192.275 -22.275 192.605 ;
        RECT -22.605 190.915 -22.275 191.245 ;
        RECT -22.605 189.555 -22.275 189.885 ;
        RECT -22.605 188.195 -22.275 188.525 ;
        RECT -22.605 186.835 -22.275 187.165 ;
        RECT -22.605 185.475 -22.275 185.805 ;
        RECT -22.605 184.115 -22.275 184.445 ;
        RECT -22.605 182.755 -22.275 183.085 ;
        RECT -22.605 181.395 -22.275 181.725 ;
        RECT -22.605 180.035 -22.275 180.365 ;
        RECT -22.605 178.675 -22.275 179.005 ;
        RECT -22.605 177.315 -22.275 177.645 ;
        RECT -22.605 175.955 -22.275 176.285 ;
        RECT -22.605 174.595 -22.275 174.925 ;
        RECT -22.605 173.235 -22.275 173.565 ;
        RECT -22.605 171.875 -22.275 172.205 ;
        RECT -22.605 170.515 -22.275 170.845 ;
        RECT -22.605 169.155 -22.275 169.485 ;
        RECT -22.605 167.795 -22.275 168.125 ;
        RECT -22.605 166.435 -22.275 166.765 ;
        RECT -22.605 165.075 -22.275 165.405 ;
        RECT -22.605 163.715 -22.275 164.045 ;
        RECT -22.605 162.355 -22.275 162.685 ;
        RECT -22.605 160.995 -22.275 161.325 ;
        RECT -22.605 159.635 -22.275 159.965 ;
        RECT -22.605 158.275 -22.275 158.605 ;
        RECT -22.605 156.915 -22.275 157.245 ;
        RECT -22.605 155.555 -22.275 155.885 ;
        RECT -22.605 154.195 -22.275 154.525 ;
        RECT -22.605 152.835 -22.275 153.165 ;
        RECT -22.605 151.475 -22.275 151.805 ;
        RECT -22.605 150.115 -22.275 150.445 ;
        RECT -22.605 148.755 -22.275 149.085 ;
        RECT -22.605 147.395 -22.275 147.725 ;
        RECT -22.605 146.035 -22.275 146.365 ;
        RECT -22.605 144.675 -22.275 145.005 ;
        RECT -22.605 143.315 -22.275 143.645 ;
        RECT -22.605 141.955 -22.275 142.285 ;
        RECT -22.605 140.595 -22.275 140.925 ;
        RECT -22.605 139.235 -22.275 139.565 ;
        RECT -22.605 137.875 -22.275 138.205 ;
        RECT -22.605 136.515 -22.275 136.845 ;
        RECT -22.605 135.155 -22.275 135.485 ;
        RECT -22.605 133.795 -22.275 134.125 ;
        RECT -22.605 132.435 -22.275 132.765 ;
        RECT -22.605 131.075 -22.275 131.405 ;
        RECT -22.605 129.715 -22.275 130.045 ;
        RECT -22.605 128.355 -22.275 128.685 ;
        RECT -22.605 126.995 -22.275 127.325 ;
        RECT -22.605 125.635 -22.275 125.965 ;
        RECT -22.605 124.275 -22.275 124.605 ;
        RECT -22.605 122.915 -22.275 123.245 ;
        RECT -22.605 121.555 -22.275 121.885 ;
        RECT -22.605 120.195 -22.275 120.525 ;
        RECT -22.605 118.835 -22.275 119.165 ;
        RECT -22.605 117.475 -22.275 117.805 ;
        RECT -22.605 116.115 -22.275 116.445 ;
        RECT -22.605 114.755 -22.275 115.085 ;
        RECT -22.605 113.395 -22.275 113.725 ;
        RECT -22.605 112.035 -22.275 112.365 ;
        RECT -22.605 110.675 -22.275 111.005 ;
        RECT -22.605 109.315 -22.275 109.645 ;
        RECT -22.605 107.955 -22.275 108.285 ;
        RECT -22.605 106.595 -22.275 106.925 ;
        RECT -22.605 105.235 -22.275 105.565 ;
        RECT -22.605 103.875 -22.275 104.205 ;
        RECT -22.605 102.515 -22.275 102.845 ;
        RECT -22.605 101.155 -22.275 101.485 ;
        RECT -22.605 99.795 -22.275 100.125 ;
        RECT -22.605 98.435 -22.275 98.765 ;
        RECT -22.605 97.075 -22.275 97.405 ;
        RECT -22.605 95.715 -22.275 96.045 ;
        RECT -22.605 94.355 -22.275 94.685 ;
        RECT -22.605 92.995 -22.275 93.325 ;
        RECT -22.605 91.635 -22.275 91.965 ;
        RECT -22.605 90.275 -22.275 90.605 ;
        RECT -22.605 88.915 -22.275 89.245 ;
        RECT -22.605 87.555 -22.275 87.885 ;
        RECT -22.605 86.195 -22.275 86.525 ;
        RECT -22.605 84.835 -22.275 85.165 ;
        RECT -22.605 83.475 -22.275 83.805 ;
        RECT -22.605 82.115 -22.275 82.445 ;
        RECT -22.605 80.755 -22.275 81.085 ;
        RECT -22.605 79.395 -22.275 79.725 ;
        RECT -22.605 78.035 -22.275 78.365 ;
        RECT -22.605 76.675 -22.275 77.005 ;
        RECT -22.605 75.315 -22.275 75.645 ;
        RECT -22.605 73.955 -22.275 74.285 ;
        RECT -22.605 72.595 -22.275 72.925 ;
        RECT -22.605 71.235 -22.275 71.565 ;
        RECT -22.605 69.875 -22.275 70.205 ;
        RECT -22.605 68.515 -22.275 68.845 ;
        RECT -22.605 67.155 -22.275 67.485 ;
        RECT -22.605 65.795 -22.275 66.125 ;
        RECT -22.605 64.435 -22.275 64.765 ;
        RECT -22.605 63.075 -22.275 63.405 ;
        RECT -22.605 61.715 -22.275 62.045 ;
        RECT -22.605 60.355 -22.275 60.685 ;
        RECT -22.605 58.995 -22.275 59.325 ;
        RECT -22.605 57.635 -22.275 57.965 ;
        RECT -22.605 56.275 -22.275 56.605 ;
        RECT -22.605 54.915 -22.275 55.245 ;
        RECT -22.605 53.555 -22.275 53.885 ;
        RECT -22.605 52.195 -22.275 52.525 ;
        RECT -22.605 50.835 -22.275 51.165 ;
        RECT -22.605 49.475 -22.275 49.805 ;
        RECT -22.605 48.115 -22.275 48.445 ;
        RECT -22.605 46.755 -22.275 47.085 ;
        RECT -22.605 45.395 -22.275 45.725 ;
        RECT -22.605 44.035 -22.275 44.365 ;
        RECT -22.605 42.675 -22.275 43.005 ;
        RECT -22.605 41.315 -22.275 41.645 ;
        RECT -22.605 39.955 -22.275 40.285 ;
        RECT -22.605 38.595 -22.275 38.925 ;
        RECT -22.605 37.235 -22.275 37.565 ;
        RECT -22.605 35.875 -22.275 36.205 ;
        RECT -22.605 34.515 -22.275 34.845 ;
        RECT -22.605 33.155 -22.275 33.485 ;
        RECT -22.605 31.795 -22.275 32.125 ;
        RECT -22.605 30.435 -22.275 30.765 ;
        RECT -22.605 29.075 -22.275 29.405 ;
        RECT -22.605 27.715 -22.275 28.045 ;
        RECT -22.605 26.355 -22.275 26.685 ;
        RECT -22.605 24.995 -22.275 25.325 ;
        RECT -22.605 23.635 -22.275 23.965 ;
        RECT -22.605 22.275 -22.275 22.605 ;
        RECT -22.605 20.915 -22.275 21.245 ;
        RECT -22.605 19.555 -22.275 19.885 ;
        RECT -22.605 18.195 -22.275 18.525 ;
        RECT -22.605 16.835 -22.275 17.165 ;
        RECT -22.605 15.475 -22.275 15.805 ;
        RECT -22.605 14.115 -22.275 14.445 ;
        RECT -22.605 12.755 -22.275 13.085 ;
        RECT -22.605 11.395 -22.275 11.725 ;
        RECT -22.605 10.035 -22.275 10.365 ;
        RECT -22.605 8.675 -22.275 9.005 ;
        RECT -22.605 7.315 -22.275 7.645 ;
        RECT -22.605 5.955 -22.275 6.285 ;
        RECT -22.605 4.595 -22.275 4.925 ;
        RECT -22.605 3.235 -22.275 3.565 ;
        RECT -22.605 1.875 -22.275 2.205 ;
        RECT -22.605 0.515 -22.275 0.845 ;
        RECT -22.605 -0.845 -22.275 -0.515 ;
        RECT -22.605 -2.205 -22.275 -1.875 ;
        RECT -22.605 -7.645 -22.275 -7.315 ;
        RECT -22.605 -9.005 -22.275 -8.675 ;
        RECT -22.605 -10.73 -22.275 -10.4 ;
        RECT -22.605 -15.805 -22.275 -15.475 ;
        RECT -22.605 -16.77 -22.275 -16.44 ;
        RECT -22.605 -18.525 -22.275 -18.195 ;
        RECT -22.605 -21.245 -22.275 -20.915 ;
        RECT -22.605 -29.405 -22.275 -29.075 ;
        RECT -22.605 -32.125 -22.275 -31.795 ;
        RECT -22.605 -33.71 -22.275 -33.38 ;
        RECT -22.605 -34.845 -22.275 -34.515 ;
        RECT -22.605 -36.205 -22.275 -35.875 ;
        RECT -22.605 -38.925 -22.275 -38.595 ;
        RECT -22.605 -39.75 -22.275 -39.42 ;
        RECT -22.605 -41.645 -22.275 -41.315 ;
        RECT -22.605 -44.365 -22.275 -44.035 ;
        RECT -22.605 -49.805 -22.275 -49.475 ;
        RECT -22.605 -51.165 -22.275 -50.835 ;
        RECT -22.605 -52.525 -22.275 -52.195 ;
        RECT -22.605 -53.885 -22.275 -53.555 ;
        RECT -22.605 -55.245 -22.275 -54.915 ;
        RECT -22.605 -56.605 -22.275 -56.275 ;
        RECT -22.605 -57.965 -22.275 -57.635 ;
        RECT -22.605 -59.325 -22.275 -58.995 ;
        RECT -22.605 -60.685 -22.275 -60.355 ;
        RECT -22.605 -62.045 -22.275 -61.715 ;
        RECT -22.605 -64.765 -22.275 -64.435 ;
        RECT -22.605 -66.125 -22.275 -65.795 ;
        RECT -22.605 -67.485 -22.275 -67.155 ;
        RECT -22.605 -68.845 -22.275 -68.515 ;
        RECT -22.605 -70.205 -22.275 -69.875 ;
        RECT -22.605 -71.565 -22.275 -71.235 ;
        RECT -22.605 -72.925 -22.275 -72.595 ;
        RECT -22.605 -74.285 -22.275 -73.955 ;
        RECT -22.605 -75.645 -22.275 -75.315 ;
        RECT -22.605 -77.005 -22.275 -76.675 ;
        RECT -22.605 -78.365 -22.275 -78.035 ;
        RECT -22.605 -79.725 -22.275 -79.395 ;
        RECT -22.605 -81.085 -22.275 -80.755 ;
        RECT -22.605 -82.445 -22.275 -82.115 ;
        RECT -22.605 -83.805 -22.275 -83.475 ;
        RECT -22.605 -85.165 -22.275 -84.835 ;
        RECT -22.605 -86.525 -22.275 -86.195 ;
        RECT -22.605 -87.885 -22.275 -87.555 ;
        RECT -22.605 -89.245 -22.275 -88.915 ;
        RECT -22.605 -90.605 -22.275 -90.275 ;
        RECT -22.605 -91.965 -22.275 -91.635 ;
        RECT -22.605 -93.325 -22.275 -92.995 ;
        RECT -22.605 -94.685 -22.275 -94.355 ;
        RECT -22.605 -96.045 -22.275 -95.715 ;
        RECT -22.605 -97.405 -22.275 -97.075 ;
        RECT -22.605 -98.765 -22.275 -98.435 ;
        RECT -22.605 -100.125 -22.275 -99.795 ;
        RECT -22.605 -101.485 -22.275 -101.155 ;
        RECT -22.605 -102.845 -22.275 -102.515 ;
        RECT -22.605 -104.205 -22.275 -103.875 ;
        RECT -22.605 -105.565 -22.275 -105.235 ;
        RECT -22.605 -106.925 -22.275 -106.595 ;
        RECT -22.605 -108.285 -22.275 -107.955 ;
        RECT -22.605 -109.645 -22.275 -109.315 ;
        RECT -22.605 -111.005 -22.275 -110.675 ;
        RECT -22.605 -113.725 -22.275 -113.395 ;
        RECT -22.605 -115.085 -22.275 -114.755 ;
        RECT -22.605 -116.445 -22.275 -116.115 ;
        RECT -22.605 -117.805 -22.275 -117.475 ;
        RECT -22.605 -119.165 -22.275 -118.835 ;
        RECT -22.605 -120.525 -22.275 -120.195 ;
        RECT -22.605 -121.885 -22.275 -121.555 ;
        RECT -22.605 -123.245 -22.275 -122.915 ;
        RECT -22.605 -124.605 -22.275 -124.275 ;
        RECT -22.605 -125.965 -22.275 -125.635 ;
        RECT -22.605 -127.325 -22.275 -126.995 ;
        RECT -22.605 -134.125 -22.275 -133.795 ;
        RECT -22.605 -135.485 -22.275 -135.155 ;
        RECT -22.605 -136.845 -22.275 -136.515 ;
        RECT -22.605 -140.925 -22.275 -140.595 ;
        RECT -22.605 -142.285 -22.275 -141.955 ;
        RECT -22.605 -143.645 -22.275 -143.315 ;
        RECT -22.605 -146.365 -22.275 -146.035 ;
        RECT -22.605 -147.725 -22.275 -147.395 ;
        RECT -22.605 -151.805 -22.275 -151.475 ;
        RECT -22.605 -155.885 -22.275 -155.555 ;
        RECT -22.605 -157.245 -22.275 -156.915 ;
        RECT -22.605 -158.605 -22.275 -158.275 ;
        RECT -22.605 -159.965 -22.275 -159.635 ;
        RECT -22.605 -161.325 -22.275 -160.995 ;
        RECT -22.605 -162.685 -22.275 -162.355 ;
        RECT -22.605 -164.045 -22.275 -163.715 ;
        RECT -22.605 -165.405 -22.275 -165.075 ;
        RECT -22.605 -166.765 -22.275 -166.435 ;
        RECT -22.605 -169.485 -22.275 -169.155 ;
        RECT -22.605 -170.845 -22.275 -170.515 ;
        RECT -22.605 -174.925 -22.275 -174.595 ;
        RECT -22.605 -177.645 -22.275 -177.315 ;
        RECT -22.605 -183.29 -22.275 -182.16 ;
        RECT -22.6 -183.405 -22.28 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -21.245 116.115 -20.915 116.445 ;
        RECT -21.245 114.755 -20.915 115.085 ;
        RECT -21.245 113.395 -20.915 113.725 ;
        RECT -21.245 112.035 -20.915 112.365 ;
        RECT -21.245 110.675 -20.915 111.005 ;
        RECT -21.245 109.315 -20.915 109.645 ;
        RECT -21.245 107.955 -20.915 108.285 ;
        RECT -21.245 106.595 -20.915 106.925 ;
        RECT -21.245 105.235 -20.915 105.565 ;
        RECT -21.245 103.875 -20.915 104.205 ;
        RECT -21.245 102.515 -20.915 102.845 ;
        RECT -21.245 101.155 -20.915 101.485 ;
        RECT -21.245 99.795 -20.915 100.125 ;
        RECT -21.245 98.435 -20.915 98.765 ;
        RECT -21.245 97.075 -20.915 97.405 ;
        RECT -21.245 95.715 -20.915 96.045 ;
        RECT -21.245 94.355 -20.915 94.685 ;
        RECT -21.245 92.995 -20.915 93.325 ;
        RECT -21.245 91.635 -20.915 91.965 ;
        RECT -21.245 90.275 -20.915 90.605 ;
        RECT -21.245 88.915 -20.915 89.245 ;
        RECT -21.245 87.555 -20.915 87.885 ;
        RECT -21.245 86.195 -20.915 86.525 ;
        RECT -21.245 84.835 -20.915 85.165 ;
        RECT -21.245 83.475 -20.915 83.805 ;
        RECT -21.245 82.115 -20.915 82.445 ;
        RECT -21.245 80.755 -20.915 81.085 ;
        RECT -21.245 79.395 -20.915 79.725 ;
        RECT -21.245 78.035 -20.915 78.365 ;
        RECT -21.245 76.675 -20.915 77.005 ;
        RECT -21.245 75.315 -20.915 75.645 ;
        RECT -21.245 73.955 -20.915 74.285 ;
        RECT -21.245 72.595 -20.915 72.925 ;
        RECT -21.245 71.235 -20.915 71.565 ;
        RECT -21.245 69.875 -20.915 70.205 ;
        RECT -21.245 68.515 -20.915 68.845 ;
        RECT -21.245 67.155 -20.915 67.485 ;
        RECT -21.245 65.795 -20.915 66.125 ;
        RECT -21.245 64.435 -20.915 64.765 ;
        RECT -21.245 63.075 -20.915 63.405 ;
        RECT -21.245 61.715 -20.915 62.045 ;
        RECT -21.245 60.355 -20.915 60.685 ;
        RECT -21.245 58.995 -20.915 59.325 ;
        RECT -21.245 57.635 -20.915 57.965 ;
        RECT -21.245 56.275 -20.915 56.605 ;
        RECT -21.245 54.915 -20.915 55.245 ;
        RECT -21.245 53.555 -20.915 53.885 ;
        RECT -21.245 52.195 -20.915 52.525 ;
        RECT -21.245 50.835 -20.915 51.165 ;
        RECT -21.245 49.475 -20.915 49.805 ;
        RECT -21.245 48.115 -20.915 48.445 ;
        RECT -21.245 46.755 -20.915 47.085 ;
        RECT -21.245 45.395 -20.915 45.725 ;
        RECT -21.245 44.035 -20.915 44.365 ;
        RECT -21.245 42.675 -20.915 43.005 ;
        RECT -21.245 41.315 -20.915 41.645 ;
        RECT -21.245 39.955 -20.915 40.285 ;
        RECT -21.245 38.595 -20.915 38.925 ;
        RECT -21.245 37.235 -20.915 37.565 ;
        RECT -21.245 35.875 -20.915 36.205 ;
        RECT -21.245 34.515 -20.915 34.845 ;
        RECT -21.245 33.155 -20.915 33.485 ;
        RECT -21.245 31.795 -20.915 32.125 ;
        RECT -21.245 30.435 -20.915 30.765 ;
        RECT -21.245 29.075 -20.915 29.405 ;
        RECT -21.245 27.715 -20.915 28.045 ;
        RECT -21.245 26.355 -20.915 26.685 ;
        RECT -21.245 24.995 -20.915 25.325 ;
        RECT -21.245 23.635 -20.915 23.965 ;
        RECT -21.245 22.275 -20.915 22.605 ;
        RECT -21.245 20.915 -20.915 21.245 ;
        RECT -21.245 19.555 -20.915 19.885 ;
        RECT -21.245 18.195 -20.915 18.525 ;
        RECT -21.245 16.835 -20.915 17.165 ;
        RECT -21.245 15.475 -20.915 15.805 ;
        RECT -21.245 14.115 -20.915 14.445 ;
        RECT -21.245 12.755 -20.915 13.085 ;
        RECT -21.245 11.395 -20.915 11.725 ;
        RECT -21.245 10.035 -20.915 10.365 ;
        RECT -21.245 8.675 -20.915 9.005 ;
        RECT -21.245 7.315 -20.915 7.645 ;
        RECT -21.245 5.955 -20.915 6.285 ;
        RECT -21.245 4.595 -20.915 4.925 ;
        RECT -21.245 3.235 -20.915 3.565 ;
        RECT -21.245 1.875 -20.915 2.205 ;
        RECT -21.245 0.515 -20.915 0.845 ;
        RECT -21.245 -0.845 -20.915 -0.515 ;
        RECT -21.245 -2.205 -20.915 -1.875 ;
        RECT -21.245 -3.565 -20.915 -3.235 ;
        RECT -21.245 -7.645 -20.915 -7.315 ;
        RECT -21.245 -9.005 -20.915 -8.675 ;
        RECT -21.245 -10.73 -20.915 -10.4 ;
        RECT -21.245 -15.805 -20.915 -15.475 ;
        RECT -21.245 -16.77 -20.915 -16.44 ;
        RECT -21.245 -18.525 -20.915 -18.195 ;
        RECT -21.245 -21.245 -20.915 -20.915 ;
        RECT -21.24 -23.28 -20.92 245.285 ;
        RECT -21.245 244.04 -20.915 245.17 ;
        RECT -21.245 239.875 -20.915 240.205 ;
        RECT -21.245 238.515 -20.915 238.845 ;
        RECT -21.245 237.155 -20.915 237.485 ;
        RECT -21.245 235.795 -20.915 236.125 ;
        RECT -21.245 234.435 -20.915 234.765 ;
        RECT -21.245 233.075 -20.915 233.405 ;
        RECT -21.245 231.715 -20.915 232.045 ;
        RECT -21.245 230.355 -20.915 230.685 ;
        RECT -21.245 228.995 -20.915 229.325 ;
        RECT -21.245 227.635 -20.915 227.965 ;
        RECT -21.245 226.275 -20.915 226.605 ;
        RECT -21.245 224.915 -20.915 225.245 ;
        RECT -21.245 223.555 -20.915 223.885 ;
        RECT -21.245 222.195 -20.915 222.525 ;
        RECT -21.245 220.835 -20.915 221.165 ;
        RECT -21.245 219.475 -20.915 219.805 ;
        RECT -21.245 218.115 -20.915 218.445 ;
        RECT -21.245 216.755 -20.915 217.085 ;
        RECT -21.245 215.395 -20.915 215.725 ;
        RECT -21.245 214.035 -20.915 214.365 ;
        RECT -21.245 212.675 -20.915 213.005 ;
        RECT -21.245 211.315 -20.915 211.645 ;
        RECT -21.245 209.955 -20.915 210.285 ;
        RECT -21.245 208.595 -20.915 208.925 ;
        RECT -21.245 207.235 -20.915 207.565 ;
        RECT -21.245 205.875 -20.915 206.205 ;
        RECT -21.245 204.515 -20.915 204.845 ;
        RECT -21.245 203.155 -20.915 203.485 ;
        RECT -21.245 201.795 -20.915 202.125 ;
        RECT -21.245 200.435 -20.915 200.765 ;
        RECT -21.245 199.075 -20.915 199.405 ;
        RECT -21.245 197.715 -20.915 198.045 ;
        RECT -21.245 196.355 -20.915 196.685 ;
        RECT -21.245 194.995 -20.915 195.325 ;
        RECT -21.245 193.635 -20.915 193.965 ;
        RECT -21.245 192.275 -20.915 192.605 ;
        RECT -21.245 190.915 -20.915 191.245 ;
        RECT -21.245 189.555 -20.915 189.885 ;
        RECT -21.245 188.195 -20.915 188.525 ;
        RECT -21.245 186.835 -20.915 187.165 ;
        RECT -21.245 185.475 -20.915 185.805 ;
        RECT -21.245 184.115 -20.915 184.445 ;
        RECT -21.245 182.755 -20.915 183.085 ;
        RECT -21.245 181.395 -20.915 181.725 ;
        RECT -21.245 180.035 -20.915 180.365 ;
        RECT -21.245 178.675 -20.915 179.005 ;
        RECT -21.245 177.315 -20.915 177.645 ;
        RECT -21.245 175.955 -20.915 176.285 ;
        RECT -21.245 174.595 -20.915 174.925 ;
        RECT -21.245 173.235 -20.915 173.565 ;
        RECT -21.245 171.875 -20.915 172.205 ;
        RECT -21.245 170.515 -20.915 170.845 ;
        RECT -21.245 169.155 -20.915 169.485 ;
        RECT -21.245 167.795 -20.915 168.125 ;
        RECT -21.245 166.435 -20.915 166.765 ;
        RECT -21.245 165.075 -20.915 165.405 ;
        RECT -21.245 163.715 -20.915 164.045 ;
        RECT -21.245 162.355 -20.915 162.685 ;
        RECT -21.245 160.995 -20.915 161.325 ;
        RECT -21.245 159.635 -20.915 159.965 ;
        RECT -21.245 158.275 -20.915 158.605 ;
        RECT -21.245 156.915 -20.915 157.245 ;
        RECT -21.245 155.555 -20.915 155.885 ;
        RECT -21.245 154.195 -20.915 154.525 ;
        RECT -21.245 152.835 -20.915 153.165 ;
        RECT -21.245 151.475 -20.915 151.805 ;
        RECT -21.245 150.115 -20.915 150.445 ;
        RECT -21.245 148.755 -20.915 149.085 ;
        RECT -21.245 147.395 -20.915 147.725 ;
        RECT -21.245 146.035 -20.915 146.365 ;
        RECT -21.245 144.675 -20.915 145.005 ;
        RECT -21.245 143.315 -20.915 143.645 ;
        RECT -21.245 141.955 -20.915 142.285 ;
        RECT -21.245 140.595 -20.915 140.925 ;
        RECT -21.245 139.235 -20.915 139.565 ;
        RECT -21.245 137.875 -20.915 138.205 ;
        RECT -21.245 136.515 -20.915 136.845 ;
        RECT -21.245 135.155 -20.915 135.485 ;
        RECT -21.245 133.795 -20.915 134.125 ;
        RECT -21.245 132.435 -20.915 132.765 ;
        RECT -21.245 131.075 -20.915 131.405 ;
        RECT -21.245 129.715 -20.915 130.045 ;
        RECT -21.245 128.355 -20.915 128.685 ;
        RECT -21.245 126.995 -20.915 127.325 ;
        RECT -21.245 125.635 -20.915 125.965 ;
        RECT -21.245 124.275 -20.915 124.605 ;
        RECT -21.245 122.915 -20.915 123.245 ;
        RECT -21.245 121.555 -20.915 121.885 ;
        RECT -21.245 120.195 -20.915 120.525 ;
        RECT -21.245 118.835 -20.915 119.165 ;
        RECT -21.245 117.475 -20.915 117.805 ;
    END
    PORT
      LAYER met3 ;
        RECT -30.765 244.04 -30.435 245.17 ;
        RECT -30.765 239.875 -30.435 240.205 ;
        RECT -30.765 238.515 -30.435 238.845 ;
        RECT -30.765 237.155 -30.435 237.485 ;
        RECT -30.765 235.795 -30.435 236.125 ;
        RECT -30.765 234.435 -30.435 234.765 ;
        RECT -30.765 233.075 -30.435 233.405 ;
        RECT -30.765 231.715 -30.435 232.045 ;
        RECT -30.765 230.355 -30.435 230.685 ;
        RECT -30.765 228.995 -30.435 229.325 ;
        RECT -30.765 227.635 -30.435 227.965 ;
        RECT -30.765 226.275 -30.435 226.605 ;
        RECT -30.765 224.915 -30.435 225.245 ;
        RECT -30.765 223.555 -30.435 223.885 ;
        RECT -30.765 222.195 -30.435 222.525 ;
        RECT -30.765 220.835 -30.435 221.165 ;
        RECT -30.765 219.475 -30.435 219.805 ;
        RECT -30.765 218.115 -30.435 218.445 ;
        RECT -30.765 216.755 -30.435 217.085 ;
        RECT -30.765 215.395 -30.435 215.725 ;
        RECT -30.765 214.035 -30.435 214.365 ;
        RECT -30.765 212.675 -30.435 213.005 ;
        RECT -30.765 211.315 -30.435 211.645 ;
        RECT -30.765 209.955 -30.435 210.285 ;
        RECT -30.765 208.595 -30.435 208.925 ;
        RECT -30.765 207.235 -30.435 207.565 ;
        RECT -30.765 205.875 -30.435 206.205 ;
        RECT -30.765 204.515 -30.435 204.845 ;
        RECT -30.765 203.155 -30.435 203.485 ;
        RECT -30.765 201.795 -30.435 202.125 ;
        RECT -30.765 200.435 -30.435 200.765 ;
        RECT -30.765 199.075 -30.435 199.405 ;
        RECT -30.765 197.715 -30.435 198.045 ;
        RECT -30.765 196.355 -30.435 196.685 ;
        RECT -30.765 194.995 -30.435 195.325 ;
        RECT -30.765 193.635 -30.435 193.965 ;
        RECT -30.765 192.275 -30.435 192.605 ;
        RECT -30.765 190.915 -30.435 191.245 ;
        RECT -30.765 189.555 -30.435 189.885 ;
        RECT -30.765 188.195 -30.435 188.525 ;
        RECT -30.765 186.835 -30.435 187.165 ;
        RECT -30.765 185.475 -30.435 185.805 ;
        RECT -30.765 184.115 -30.435 184.445 ;
        RECT -30.765 182.755 -30.435 183.085 ;
        RECT -30.765 181.395 -30.435 181.725 ;
        RECT -30.765 180.035 -30.435 180.365 ;
        RECT -30.765 178.675 -30.435 179.005 ;
        RECT -30.765 177.315 -30.435 177.645 ;
        RECT -30.765 175.955 -30.435 176.285 ;
        RECT -30.765 174.595 -30.435 174.925 ;
        RECT -30.765 173.235 -30.435 173.565 ;
        RECT -30.765 171.875 -30.435 172.205 ;
        RECT -30.765 170.515 -30.435 170.845 ;
        RECT -30.765 169.155 -30.435 169.485 ;
        RECT -30.765 167.795 -30.435 168.125 ;
        RECT -30.765 166.435 -30.435 166.765 ;
        RECT -30.765 165.075 -30.435 165.405 ;
        RECT -30.765 163.715 -30.435 164.045 ;
        RECT -30.765 162.355 -30.435 162.685 ;
        RECT -30.765 160.995 -30.435 161.325 ;
        RECT -30.765 159.635 -30.435 159.965 ;
        RECT -30.765 158.275 -30.435 158.605 ;
        RECT -30.765 156.915 -30.435 157.245 ;
        RECT -30.765 155.555 -30.435 155.885 ;
        RECT -30.765 154.195 -30.435 154.525 ;
        RECT -30.765 152.835 -30.435 153.165 ;
        RECT -30.765 151.475 -30.435 151.805 ;
        RECT -30.765 150.115 -30.435 150.445 ;
        RECT -30.765 148.755 -30.435 149.085 ;
        RECT -30.765 147.395 -30.435 147.725 ;
        RECT -30.765 146.035 -30.435 146.365 ;
        RECT -30.765 144.675 -30.435 145.005 ;
        RECT -30.765 143.315 -30.435 143.645 ;
        RECT -30.765 141.955 -30.435 142.285 ;
        RECT -30.765 140.595 -30.435 140.925 ;
        RECT -30.765 139.235 -30.435 139.565 ;
        RECT -30.765 137.875 -30.435 138.205 ;
        RECT -30.765 136.515 -30.435 136.845 ;
        RECT -30.765 135.155 -30.435 135.485 ;
        RECT -30.765 133.795 -30.435 134.125 ;
        RECT -30.765 132.435 -30.435 132.765 ;
        RECT -30.765 131.075 -30.435 131.405 ;
        RECT -30.765 129.715 -30.435 130.045 ;
        RECT -30.765 128.355 -30.435 128.685 ;
        RECT -30.765 126.995 -30.435 127.325 ;
        RECT -30.765 125.635 -30.435 125.965 ;
        RECT -30.765 124.275 -30.435 124.605 ;
        RECT -30.765 122.915 -30.435 123.245 ;
        RECT -30.765 121.555 -30.435 121.885 ;
        RECT -30.765 120.195 -30.435 120.525 ;
        RECT -30.765 118.835 -30.435 119.165 ;
        RECT -30.765 117.475 -30.435 117.805 ;
        RECT -30.765 116.115 -30.435 116.445 ;
        RECT -30.765 114.755 -30.435 115.085 ;
        RECT -30.765 113.395 -30.435 113.725 ;
        RECT -30.765 112.035 -30.435 112.365 ;
        RECT -30.765 110.675 -30.435 111.005 ;
        RECT -30.765 109.315 -30.435 109.645 ;
        RECT -30.765 107.955 -30.435 108.285 ;
        RECT -30.765 106.595 -30.435 106.925 ;
        RECT -30.765 105.235 -30.435 105.565 ;
        RECT -30.765 103.875 -30.435 104.205 ;
        RECT -30.765 102.515 -30.435 102.845 ;
        RECT -30.765 101.155 -30.435 101.485 ;
        RECT -30.765 99.795 -30.435 100.125 ;
        RECT -30.765 98.435 -30.435 98.765 ;
        RECT -30.765 97.075 -30.435 97.405 ;
        RECT -30.765 95.715 -30.435 96.045 ;
        RECT -30.765 94.355 -30.435 94.685 ;
        RECT -30.765 92.995 -30.435 93.325 ;
        RECT -30.765 91.635 -30.435 91.965 ;
        RECT -30.765 90.275 -30.435 90.605 ;
        RECT -30.765 88.915 -30.435 89.245 ;
        RECT -30.765 87.555 -30.435 87.885 ;
        RECT -30.765 86.195 -30.435 86.525 ;
        RECT -30.765 84.835 -30.435 85.165 ;
        RECT -30.765 83.475 -30.435 83.805 ;
        RECT -30.765 82.115 -30.435 82.445 ;
        RECT -30.765 80.755 -30.435 81.085 ;
        RECT -30.765 79.395 -30.435 79.725 ;
        RECT -30.765 78.035 -30.435 78.365 ;
        RECT -30.765 76.675 -30.435 77.005 ;
        RECT -30.765 75.315 -30.435 75.645 ;
        RECT -30.765 73.955 -30.435 74.285 ;
        RECT -30.765 72.595 -30.435 72.925 ;
        RECT -30.765 71.235 -30.435 71.565 ;
        RECT -30.765 69.875 -30.435 70.205 ;
        RECT -30.765 68.515 -30.435 68.845 ;
        RECT -30.765 67.155 -30.435 67.485 ;
        RECT -30.765 65.795 -30.435 66.125 ;
        RECT -30.765 64.435 -30.435 64.765 ;
        RECT -30.765 63.075 -30.435 63.405 ;
        RECT -30.765 61.715 -30.435 62.045 ;
        RECT -30.765 60.355 -30.435 60.685 ;
        RECT -30.765 58.995 -30.435 59.325 ;
        RECT -30.765 57.635 -30.435 57.965 ;
        RECT -30.765 56.275 -30.435 56.605 ;
        RECT -30.765 54.915 -30.435 55.245 ;
        RECT -30.765 53.555 -30.435 53.885 ;
        RECT -30.765 52.195 -30.435 52.525 ;
        RECT -30.765 50.835 -30.435 51.165 ;
        RECT -30.765 49.475 -30.435 49.805 ;
        RECT -30.765 48.115 -30.435 48.445 ;
        RECT -30.765 46.755 -30.435 47.085 ;
        RECT -30.765 45.395 -30.435 45.725 ;
        RECT -30.765 44.035 -30.435 44.365 ;
        RECT -30.765 42.675 -30.435 43.005 ;
        RECT -30.765 41.315 -30.435 41.645 ;
        RECT -30.765 39.955 -30.435 40.285 ;
        RECT -30.765 38.595 -30.435 38.925 ;
        RECT -30.765 37.235 -30.435 37.565 ;
        RECT -30.765 35.875 -30.435 36.205 ;
        RECT -30.765 34.515 -30.435 34.845 ;
        RECT -30.765 33.155 -30.435 33.485 ;
        RECT -30.765 31.795 -30.435 32.125 ;
        RECT -30.765 30.435 -30.435 30.765 ;
        RECT -30.765 29.075 -30.435 29.405 ;
        RECT -30.765 27.715 -30.435 28.045 ;
        RECT -30.765 26.355 -30.435 26.685 ;
        RECT -30.765 24.995 -30.435 25.325 ;
        RECT -30.765 23.635 -30.435 23.965 ;
        RECT -30.765 22.275 -30.435 22.605 ;
        RECT -30.765 20.915 -30.435 21.245 ;
        RECT -30.765 19.555 -30.435 19.885 ;
        RECT -30.765 18.195 -30.435 18.525 ;
        RECT -30.765 16.835 -30.435 17.165 ;
        RECT -30.765 15.475 -30.435 15.805 ;
        RECT -30.765 14.115 -30.435 14.445 ;
        RECT -30.765 12.755 -30.435 13.085 ;
        RECT -30.765 11.395 -30.435 11.725 ;
        RECT -30.765 10.035 -30.435 10.365 ;
        RECT -30.765 8.675 -30.435 9.005 ;
        RECT -30.765 7.315 -30.435 7.645 ;
        RECT -30.765 5.955 -30.435 6.285 ;
        RECT -30.765 4.595 -30.435 4.925 ;
        RECT -30.765 3.235 -30.435 3.565 ;
        RECT -30.765 1.875 -30.435 2.205 ;
        RECT -30.765 0.515 -30.435 0.845 ;
        RECT -30.765 -0.845 -30.435 -0.515 ;
        RECT -30.765 -7.645 -30.435 -7.315 ;
        RECT -30.765 -9.005 -30.435 -8.675 ;
        RECT -30.765 -10.365 -30.435 -10.035 ;
        RECT -30.765 -14.445 -30.435 -14.115 ;
        RECT -30.765 -15.805 -30.435 -15.475 ;
        RECT -30.765 -17.165 -30.435 -16.835 ;
        RECT -30.765 -18.525 -30.435 -18.195 ;
        RECT -30.765 -19.885 -30.435 -19.555 ;
        RECT -30.765 -21.245 -30.435 -20.915 ;
        RECT -30.765 -22.605 -30.435 -22.275 ;
        RECT -30.765 -23.965 -30.435 -23.635 ;
        RECT -30.765 -25.325 -30.435 -24.995 ;
        RECT -30.765 -32.125 -30.435 -31.795 ;
        RECT -30.765 -33.71 -30.435 -33.38 ;
        RECT -30.765 -34.845 -30.435 -34.515 ;
        RECT -30.765 -36.205 -30.435 -35.875 ;
        RECT -30.765 -38.925 -30.435 -38.595 ;
        RECT -30.765 -39.75 -30.435 -39.42 ;
        RECT -30.765 -41.645 -30.435 -41.315 ;
        RECT -30.765 -44.365 -30.435 -44.035 ;
        RECT -30.765 -49.805 -30.435 -49.475 ;
        RECT -30.765 -51.165 -30.435 -50.835 ;
        RECT -30.765 -53.885 -30.435 -53.555 ;
        RECT -30.765 -55.245 -30.435 -54.915 ;
        RECT -30.765 -59.325 -30.435 -58.995 ;
        RECT -30.765 -60.685 -30.435 -60.355 ;
        RECT -30.76 -64.76 -30.44 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -30.765 -70.205 -30.435 -69.875 ;
        RECT -30.765 -71.565 -30.435 -71.235 ;
        RECT -30.765 -72.925 -30.435 -72.595 ;
        RECT -30.765 -74.285 -30.435 -73.955 ;
        RECT -30.765 -75.645 -30.435 -75.315 ;
        RECT -30.765 -77.005 -30.435 -76.675 ;
        RECT -30.765 -78.365 -30.435 -78.035 ;
        RECT -30.765 -79.725 -30.435 -79.395 ;
        RECT -30.765 -81.085 -30.435 -80.755 ;
        RECT -30.765 -82.445 -30.435 -82.115 ;
        RECT -30.765 -83.805 -30.435 -83.475 ;
        RECT -30.765 -85.165 -30.435 -84.835 ;
        RECT -30.765 -86.525 -30.435 -86.195 ;
        RECT -30.765 -87.885 -30.435 -87.555 ;
        RECT -30.765 -89.245 -30.435 -88.915 ;
        RECT -30.765 -90.81 -30.435 -90.48 ;
        RECT -30.765 -91.965 -30.435 -91.635 ;
        RECT -30.765 -93.325 -30.435 -92.995 ;
        RECT -30.765 -94.685 -30.435 -94.355 ;
        RECT -30.765 -96.045 -30.435 -95.715 ;
        RECT -30.765 -97.405 -30.435 -97.075 ;
        RECT -30.765 -100.125 -30.435 -99.795 ;
        RECT -30.765 -101.35 -30.435 -101.02 ;
        RECT -30.765 -102.845 -30.435 -102.515 ;
        RECT -30.765 -104.205 -30.435 -103.875 ;
        RECT -30.765 -105.565 -30.435 -105.235 ;
        RECT -30.765 -108.285 -30.435 -107.955 ;
        RECT -30.765 -109.645 -30.435 -109.315 ;
        RECT -30.765 -112.365 -30.435 -112.035 ;
        RECT -30.765 -113.725 -30.435 -113.395 ;
        RECT -30.765 -115.085 -30.435 -114.755 ;
        RECT -30.765 -116.445 -30.435 -116.115 ;
        RECT -30.765 -117.805 -30.435 -117.475 ;
        RECT -30.765 -119.165 -30.435 -118.835 ;
        RECT -30.765 -120.525 -30.435 -120.195 ;
        RECT -30.765 -121.885 -30.435 -121.555 ;
        RECT -30.765 -123.245 -30.435 -122.915 ;
        RECT -30.765 -124.605 -30.435 -124.275 ;
        RECT -30.765 -125.965 -30.435 -125.635 ;
        RECT -30.765 -127.325 -30.435 -126.995 ;
        RECT -30.765 -128.685 -30.435 -128.355 ;
        RECT -30.765 -132.765 -30.435 -132.435 ;
        RECT -30.765 -134.125 -30.435 -133.795 ;
        RECT -30.765 -135.485 -30.435 -135.155 ;
        RECT -30.765 -136.845 -30.435 -136.515 ;
        RECT -30.765 -140.925 -30.435 -140.595 ;
        RECT -30.765 -142.285 -30.435 -141.955 ;
        RECT -30.765 -143.645 -30.435 -143.315 ;
        RECT -30.765 -145.005 -30.435 -144.675 ;
        RECT -30.765 -146.365 -30.435 -146.035 ;
        RECT -30.765 -147.725 -30.435 -147.395 ;
        RECT -30.765 -150.445 -30.435 -150.115 ;
        RECT -30.765 -151.805 -30.435 -151.475 ;
        RECT -30.765 -155.885 -30.435 -155.555 ;
        RECT -30.765 -157.245 -30.435 -156.915 ;
        RECT -30.765 -158.605 -30.435 -158.275 ;
        RECT -30.765 -159.965 -30.435 -159.635 ;
        RECT -30.765 -161.325 -30.435 -160.995 ;
        RECT -30.765 -162.685 -30.435 -162.355 ;
        RECT -30.765 -164.045 -30.435 -163.715 ;
        RECT -30.765 -165.405 -30.435 -165.075 ;
        RECT -30.765 -166.765 -30.435 -166.435 ;
        RECT -30.765 -168.655 -30.435 -168.325 ;
        RECT -30.765 -169.485 -30.435 -169.155 ;
        RECT -30.765 -170.845 -30.435 -170.515 ;
        RECT -30.765 -172.205 -30.435 -171.875 ;
        RECT -30.765 -173.565 -30.435 -173.235 ;
        RECT -30.765 -174.925 -30.435 -174.595 ;
        RECT -30.765 -177.645 -30.435 -177.315 ;
        RECT -30.765 -183.29 -30.435 -182.16 ;
        RECT -30.76 -183.405 -30.44 -69.2 ;
    END
    PORT
      LAYER met3 ;
        RECT -29.405 244.04 -29.075 245.17 ;
        RECT -29.405 239.875 -29.075 240.205 ;
        RECT -29.405 238.515 -29.075 238.845 ;
        RECT -29.405 237.155 -29.075 237.485 ;
        RECT -29.405 235.795 -29.075 236.125 ;
        RECT -29.405 234.435 -29.075 234.765 ;
        RECT -29.405 233.075 -29.075 233.405 ;
        RECT -29.405 231.715 -29.075 232.045 ;
        RECT -29.405 230.355 -29.075 230.685 ;
        RECT -29.405 228.995 -29.075 229.325 ;
        RECT -29.405 227.635 -29.075 227.965 ;
        RECT -29.405 226.275 -29.075 226.605 ;
        RECT -29.405 224.915 -29.075 225.245 ;
        RECT -29.405 223.555 -29.075 223.885 ;
        RECT -29.405 222.195 -29.075 222.525 ;
        RECT -29.405 220.835 -29.075 221.165 ;
        RECT -29.405 219.475 -29.075 219.805 ;
        RECT -29.405 218.115 -29.075 218.445 ;
        RECT -29.405 216.755 -29.075 217.085 ;
        RECT -29.405 215.395 -29.075 215.725 ;
        RECT -29.405 214.035 -29.075 214.365 ;
        RECT -29.405 212.675 -29.075 213.005 ;
        RECT -29.405 211.315 -29.075 211.645 ;
        RECT -29.405 209.955 -29.075 210.285 ;
        RECT -29.405 208.595 -29.075 208.925 ;
        RECT -29.405 207.235 -29.075 207.565 ;
        RECT -29.405 205.875 -29.075 206.205 ;
        RECT -29.405 204.515 -29.075 204.845 ;
        RECT -29.405 203.155 -29.075 203.485 ;
        RECT -29.405 201.795 -29.075 202.125 ;
        RECT -29.405 200.435 -29.075 200.765 ;
        RECT -29.405 199.075 -29.075 199.405 ;
        RECT -29.405 197.715 -29.075 198.045 ;
        RECT -29.405 196.355 -29.075 196.685 ;
        RECT -29.405 194.995 -29.075 195.325 ;
        RECT -29.405 193.635 -29.075 193.965 ;
        RECT -29.405 192.275 -29.075 192.605 ;
        RECT -29.405 190.915 -29.075 191.245 ;
        RECT -29.405 189.555 -29.075 189.885 ;
        RECT -29.405 188.195 -29.075 188.525 ;
        RECT -29.405 186.835 -29.075 187.165 ;
        RECT -29.405 185.475 -29.075 185.805 ;
        RECT -29.405 184.115 -29.075 184.445 ;
        RECT -29.405 182.755 -29.075 183.085 ;
        RECT -29.405 181.395 -29.075 181.725 ;
        RECT -29.405 180.035 -29.075 180.365 ;
        RECT -29.405 178.675 -29.075 179.005 ;
        RECT -29.405 177.315 -29.075 177.645 ;
        RECT -29.405 175.955 -29.075 176.285 ;
        RECT -29.405 174.595 -29.075 174.925 ;
        RECT -29.405 173.235 -29.075 173.565 ;
        RECT -29.405 171.875 -29.075 172.205 ;
        RECT -29.405 170.515 -29.075 170.845 ;
        RECT -29.405 169.155 -29.075 169.485 ;
        RECT -29.405 167.795 -29.075 168.125 ;
        RECT -29.405 166.435 -29.075 166.765 ;
        RECT -29.405 165.075 -29.075 165.405 ;
        RECT -29.405 163.715 -29.075 164.045 ;
        RECT -29.405 162.355 -29.075 162.685 ;
        RECT -29.405 160.995 -29.075 161.325 ;
        RECT -29.405 159.635 -29.075 159.965 ;
        RECT -29.405 158.275 -29.075 158.605 ;
        RECT -29.405 156.915 -29.075 157.245 ;
        RECT -29.405 155.555 -29.075 155.885 ;
        RECT -29.405 154.195 -29.075 154.525 ;
        RECT -29.405 152.835 -29.075 153.165 ;
        RECT -29.405 151.475 -29.075 151.805 ;
        RECT -29.405 150.115 -29.075 150.445 ;
        RECT -29.405 148.755 -29.075 149.085 ;
        RECT -29.405 147.395 -29.075 147.725 ;
        RECT -29.405 146.035 -29.075 146.365 ;
        RECT -29.405 144.675 -29.075 145.005 ;
        RECT -29.405 143.315 -29.075 143.645 ;
        RECT -29.405 141.955 -29.075 142.285 ;
        RECT -29.405 140.595 -29.075 140.925 ;
        RECT -29.405 139.235 -29.075 139.565 ;
        RECT -29.405 137.875 -29.075 138.205 ;
        RECT -29.405 136.515 -29.075 136.845 ;
        RECT -29.405 135.155 -29.075 135.485 ;
        RECT -29.405 133.795 -29.075 134.125 ;
        RECT -29.405 132.435 -29.075 132.765 ;
        RECT -29.405 131.075 -29.075 131.405 ;
        RECT -29.405 129.715 -29.075 130.045 ;
        RECT -29.405 128.355 -29.075 128.685 ;
        RECT -29.405 126.995 -29.075 127.325 ;
        RECT -29.405 125.635 -29.075 125.965 ;
        RECT -29.405 124.275 -29.075 124.605 ;
        RECT -29.405 122.915 -29.075 123.245 ;
        RECT -29.405 121.555 -29.075 121.885 ;
        RECT -29.405 120.195 -29.075 120.525 ;
        RECT -29.405 118.835 -29.075 119.165 ;
        RECT -29.405 117.475 -29.075 117.805 ;
        RECT -29.405 116.115 -29.075 116.445 ;
        RECT -29.405 114.755 -29.075 115.085 ;
        RECT -29.405 113.395 -29.075 113.725 ;
        RECT -29.405 112.035 -29.075 112.365 ;
        RECT -29.405 110.675 -29.075 111.005 ;
        RECT -29.405 109.315 -29.075 109.645 ;
        RECT -29.405 107.955 -29.075 108.285 ;
        RECT -29.405 106.595 -29.075 106.925 ;
        RECT -29.405 105.235 -29.075 105.565 ;
        RECT -29.405 103.875 -29.075 104.205 ;
        RECT -29.405 102.515 -29.075 102.845 ;
        RECT -29.405 101.155 -29.075 101.485 ;
        RECT -29.405 99.795 -29.075 100.125 ;
        RECT -29.405 98.435 -29.075 98.765 ;
        RECT -29.405 97.075 -29.075 97.405 ;
        RECT -29.405 95.715 -29.075 96.045 ;
        RECT -29.405 94.355 -29.075 94.685 ;
        RECT -29.405 92.995 -29.075 93.325 ;
        RECT -29.405 91.635 -29.075 91.965 ;
        RECT -29.405 90.275 -29.075 90.605 ;
        RECT -29.405 88.915 -29.075 89.245 ;
        RECT -29.405 87.555 -29.075 87.885 ;
        RECT -29.405 86.195 -29.075 86.525 ;
        RECT -29.405 84.835 -29.075 85.165 ;
        RECT -29.405 83.475 -29.075 83.805 ;
        RECT -29.405 82.115 -29.075 82.445 ;
        RECT -29.405 80.755 -29.075 81.085 ;
        RECT -29.405 79.395 -29.075 79.725 ;
        RECT -29.405 78.035 -29.075 78.365 ;
        RECT -29.405 76.675 -29.075 77.005 ;
        RECT -29.405 75.315 -29.075 75.645 ;
        RECT -29.405 73.955 -29.075 74.285 ;
        RECT -29.405 72.595 -29.075 72.925 ;
        RECT -29.405 71.235 -29.075 71.565 ;
        RECT -29.405 69.875 -29.075 70.205 ;
        RECT -29.405 68.515 -29.075 68.845 ;
        RECT -29.405 67.155 -29.075 67.485 ;
        RECT -29.405 65.795 -29.075 66.125 ;
        RECT -29.405 64.435 -29.075 64.765 ;
        RECT -29.405 63.075 -29.075 63.405 ;
        RECT -29.405 61.715 -29.075 62.045 ;
        RECT -29.405 60.355 -29.075 60.685 ;
        RECT -29.405 58.995 -29.075 59.325 ;
        RECT -29.405 57.635 -29.075 57.965 ;
        RECT -29.405 56.275 -29.075 56.605 ;
        RECT -29.405 54.915 -29.075 55.245 ;
        RECT -29.405 53.555 -29.075 53.885 ;
        RECT -29.405 52.195 -29.075 52.525 ;
        RECT -29.405 50.835 -29.075 51.165 ;
        RECT -29.405 49.475 -29.075 49.805 ;
        RECT -29.405 48.115 -29.075 48.445 ;
        RECT -29.405 46.755 -29.075 47.085 ;
        RECT -29.405 45.395 -29.075 45.725 ;
        RECT -29.405 44.035 -29.075 44.365 ;
        RECT -29.405 42.675 -29.075 43.005 ;
        RECT -29.405 41.315 -29.075 41.645 ;
        RECT -29.405 39.955 -29.075 40.285 ;
        RECT -29.405 38.595 -29.075 38.925 ;
        RECT -29.405 37.235 -29.075 37.565 ;
        RECT -29.405 35.875 -29.075 36.205 ;
        RECT -29.405 34.515 -29.075 34.845 ;
        RECT -29.405 33.155 -29.075 33.485 ;
        RECT -29.405 31.795 -29.075 32.125 ;
        RECT -29.405 30.435 -29.075 30.765 ;
        RECT -29.405 29.075 -29.075 29.405 ;
        RECT -29.405 27.715 -29.075 28.045 ;
        RECT -29.405 26.355 -29.075 26.685 ;
        RECT -29.405 24.995 -29.075 25.325 ;
        RECT -29.405 23.635 -29.075 23.965 ;
        RECT -29.405 22.275 -29.075 22.605 ;
        RECT -29.405 20.915 -29.075 21.245 ;
        RECT -29.405 19.555 -29.075 19.885 ;
        RECT -29.405 18.195 -29.075 18.525 ;
        RECT -29.405 16.835 -29.075 17.165 ;
        RECT -29.405 15.475 -29.075 15.805 ;
        RECT -29.405 14.115 -29.075 14.445 ;
        RECT -29.405 12.755 -29.075 13.085 ;
        RECT -29.405 11.395 -29.075 11.725 ;
        RECT -29.405 10.035 -29.075 10.365 ;
        RECT -29.405 8.675 -29.075 9.005 ;
        RECT -29.405 7.315 -29.075 7.645 ;
        RECT -29.405 5.955 -29.075 6.285 ;
        RECT -29.405 4.595 -29.075 4.925 ;
        RECT -29.405 3.235 -29.075 3.565 ;
        RECT -29.405 1.875 -29.075 2.205 ;
        RECT -29.405 0.515 -29.075 0.845 ;
        RECT -29.405 -0.845 -29.075 -0.515 ;
        RECT -29.405 -7.645 -29.075 -7.315 ;
        RECT -29.405 -9.005 -29.075 -8.675 ;
        RECT -29.405 -10.73 -29.075 -10.4 ;
        RECT -29.405 -15.805 -29.075 -15.475 ;
        RECT -29.405 -16.77 -29.075 -16.44 ;
        RECT -29.405 -18.525 -29.075 -18.195 ;
        RECT -29.405 -21.245 -29.075 -20.915 ;
        RECT -29.405 -32.125 -29.075 -31.795 ;
        RECT -29.405 -33.71 -29.075 -33.38 ;
        RECT -29.405 -34.845 -29.075 -34.515 ;
        RECT -29.405 -36.205 -29.075 -35.875 ;
        RECT -29.405 -38.925 -29.075 -38.595 ;
        RECT -29.405 -39.75 -29.075 -39.42 ;
        RECT -29.405 -41.645 -29.075 -41.315 ;
        RECT -29.405 -44.365 -29.075 -44.035 ;
        RECT -29.405 -49.805 -29.075 -49.475 ;
        RECT -29.405 -51.165 -29.075 -50.835 ;
        RECT -29.405 -53.885 -29.075 -53.555 ;
        RECT -29.405 -55.245 -29.075 -54.915 ;
        RECT -29.405 -59.325 -29.075 -58.995 ;
        RECT -29.405 -60.685 -29.075 -60.355 ;
        RECT -29.4 -64.08 -29.08 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -29.405 -70.205 -29.075 -69.875 ;
        RECT -29.405 -71.565 -29.075 -71.235 ;
        RECT -29.405 -72.925 -29.075 -72.595 ;
        RECT -29.405 -74.285 -29.075 -73.955 ;
        RECT -29.405 -75.645 -29.075 -75.315 ;
        RECT -29.405 -77.005 -29.075 -76.675 ;
        RECT -29.405 -78.365 -29.075 -78.035 ;
        RECT -29.405 -79.725 -29.075 -79.395 ;
        RECT -29.405 -81.085 -29.075 -80.755 ;
        RECT -29.405 -82.445 -29.075 -82.115 ;
        RECT -29.405 -83.805 -29.075 -83.475 ;
        RECT -29.405 -85.165 -29.075 -84.835 ;
        RECT -29.405 -86.525 -29.075 -86.195 ;
        RECT -29.405 -87.885 -29.075 -87.555 ;
        RECT -29.405 -89.245 -29.075 -88.915 ;
        RECT -29.405 -90.81 -29.075 -90.48 ;
        RECT -29.405 -91.965 -29.075 -91.635 ;
        RECT -29.405 -93.325 -29.075 -92.995 ;
        RECT -29.405 -94.685 -29.075 -94.355 ;
        RECT -29.405 -96.045 -29.075 -95.715 ;
        RECT -29.405 -97.405 -29.075 -97.075 ;
        RECT -29.405 -100.125 -29.075 -99.795 ;
        RECT -29.405 -101.35 -29.075 -101.02 ;
        RECT -29.405 -102.845 -29.075 -102.515 ;
        RECT -29.405 -104.205 -29.075 -103.875 ;
        RECT -29.405 -105.565 -29.075 -105.235 ;
        RECT -29.405 -108.285 -29.075 -107.955 ;
        RECT -29.405 -109.645 -29.075 -109.315 ;
        RECT -29.4 -111.68 -29.08 -67.84 ;
    END
    PORT
      LAYER met3 ;
        RECT -29.405 -174.925 -29.075 -174.595 ;
        RECT -29.405 -177.645 -29.075 -177.315 ;
        RECT -29.405 -183.29 -29.075 -182.16 ;
        RECT -29.4 -183.405 -29.08 -173.92 ;
    END
    PORT
      LAYER met3 ;
        RECT -28.045 244.04 -27.715 245.17 ;
        RECT -28.045 239.875 -27.715 240.205 ;
        RECT -28.045 238.515 -27.715 238.845 ;
        RECT -28.045 237.155 -27.715 237.485 ;
        RECT -28.045 235.795 -27.715 236.125 ;
        RECT -28.045 234.435 -27.715 234.765 ;
        RECT -28.045 233.075 -27.715 233.405 ;
        RECT -28.045 231.715 -27.715 232.045 ;
        RECT -28.045 230.355 -27.715 230.685 ;
        RECT -28.045 228.995 -27.715 229.325 ;
        RECT -28.045 227.635 -27.715 227.965 ;
        RECT -28.045 226.275 -27.715 226.605 ;
        RECT -28.045 224.915 -27.715 225.245 ;
        RECT -28.045 223.555 -27.715 223.885 ;
        RECT -28.045 222.195 -27.715 222.525 ;
        RECT -28.045 220.835 -27.715 221.165 ;
        RECT -28.045 219.475 -27.715 219.805 ;
        RECT -28.045 218.115 -27.715 218.445 ;
        RECT -28.045 216.755 -27.715 217.085 ;
        RECT -28.045 215.395 -27.715 215.725 ;
        RECT -28.045 214.035 -27.715 214.365 ;
        RECT -28.045 212.675 -27.715 213.005 ;
        RECT -28.045 211.315 -27.715 211.645 ;
        RECT -28.045 209.955 -27.715 210.285 ;
        RECT -28.045 208.595 -27.715 208.925 ;
        RECT -28.045 207.235 -27.715 207.565 ;
        RECT -28.045 205.875 -27.715 206.205 ;
        RECT -28.045 204.515 -27.715 204.845 ;
        RECT -28.045 203.155 -27.715 203.485 ;
        RECT -28.045 201.795 -27.715 202.125 ;
        RECT -28.045 200.435 -27.715 200.765 ;
        RECT -28.045 199.075 -27.715 199.405 ;
        RECT -28.045 197.715 -27.715 198.045 ;
        RECT -28.045 196.355 -27.715 196.685 ;
        RECT -28.045 194.995 -27.715 195.325 ;
        RECT -28.045 193.635 -27.715 193.965 ;
        RECT -28.045 192.275 -27.715 192.605 ;
        RECT -28.045 190.915 -27.715 191.245 ;
        RECT -28.045 189.555 -27.715 189.885 ;
        RECT -28.045 188.195 -27.715 188.525 ;
        RECT -28.045 186.835 -27.715 187.165 ;
        RECT -28.045 185.475 -27.715 185.805 ;
        RECT -28.045 184.115 -27.715 184.445 ;
        RECT -28.045 182.755 -27.715 183.085 ;
        RECT -28.045 181.395 -27.715 181.725 ;
        RECT -28.045 180.035 -27.715 180.365 ;
        RECT -28.045 178.675 -27.715 179.005 ;
        RECT -28.045 177.315 -27.715 177.645 ;
        RECT -28.045 175.955 -27.715 176.285 ;
        RECT -28.045 174.595 -27.715 174.925 ;
        RECT -28.045 173.235 -27.715 173.565 ;
        RECT -28.045 171.875 -27.715 172.205 ;
        RECT -28.045 170.515 -27.715 170.845 ;
        RECT -28.045 169.155 -27.715 169.485 ;
        RECT -28.045 167.795 -27.715 168.125 ;
        RECT -28.045 166.435 -27.715 166.765 ;
        RECT -28.045 165.075 -27.715 165.405 ;
        RECT -28.045 163.715 -27.715 164.045 ;
        RECT -28.045 162.355 -27.715 162.685 ;
        RECT -28.045 160.995 -27.715 161.325 ;
        RECT -28.045 159.635 -27.715 159.965 ;
        RECT -28.045 158.275 -27.715 158.605 ;
        RECT -28.045 156.915 -27.715 157.245 ;
        RECT -28.045 155.555 -27.715 155.885 ;
        RECT -28.045 154.195 -27.715 154.525 ;
        RECT -28.045 152.835 -27.715 153.165 ;
        RECT -28.045 151.475 -27.715 151.805 ;
        RECT -28.045 150.115 -27.715 150.445 ;
        RECT -28.045 148.755 -27.715 149.085 ;
        RECT -28.045 147.395 -27.715 147.725 ;
        RECT -28.045 146.035 -27.715 146.365 ;
        RECT -28.045 144.675 -27.715 145.005 ;
        RECT -28.045 143.315 -27.715 143.645 ;
        RECT -28.045 141.955 -27.715 142.285 ;
        RECT -28.045 140.595 -27.715 140.925 ;
        RECT -28.045 139.235 -27.715 139.565 ;
        RECT -28.045 137.875 -27.715 138.205 ;
        RECT -28.045 136.515 -27.715 136.845 ;
        RECT -28.045 135.155 -27.715 135.485 ;
        RECT -28.045 133.795 -27.715 134.125 ;
        RECT -28.045 132.435 -27.715 132.765 ;
        RECT -28.045 131.075 -27.715 131.405 ;
        RECT -28.045 129.715 -27.715 130.045 ;
        RECT -28.045 128.355 -27.715 128.685 ;
        RECT -28.045 126.995 -27.715 127.325 ;
        RECT -28.045 125.635 -27.715 125.965 ;
        RECT -28.045 124.275 -27.715 124.605 ;
        RECT -28.045 122.915 -27.715 123.245 ;
        RECT -28.045 121.555 -27.715 121.885 ;
        RECT -28.045 120.195 -27.715 120.525 ;
        RECT -28.045 118.835 -27.715 119.165 ;
        RECT -28.045 117.475 -27.715 117.805 ;
        RECT -28.045 116.115 -27.715 116.445 ;
        RECT -28.045 114.755 -27.715 115.085 ;
        RECT -28.045 113.395 -27.715 113.725 ;
        RECT -28.045 112.035 -27.715 112.365 ;
        RECT -28.045 110.675 -27.715 111.005 ;
        RECT -28.045 109.315 -27.715 109.645 ;
        RECT -28.045 107.955 -27.715 108.285 ;
        RECT -28.045 106.595 -27.715 106.925 ;
        RECT -28.045 105.235 -27.715 105.565 ;
        RECT -28.045 103.875 -27.715 104.205 ;
        RECT -28.045 102.515 -27.715 102.845 ;
        RECT -28.045 101.155 -27.715 101.485 ;
        RECT -28.045 99.795 -27.715 100.125 ;
        RECT -28.045 98.435 -27.715 98.765 ;
        RECT -28.045 97.075 -27.715 97.405 ;
        RECT -28.045 95.715 -27.715 96.045 ;
        RECT -28.045 94.355 -27.715 94.685 ;
        RECT -28.045 92.995 -27.715 93.325 ;
        RECT -28.045 91.635 -27.715 91.965 ;
        RECT -28.045 90.275 -27.715 90.605 ;
        RECT -28.045 88.915 -27.715 89.245 ;
        RECT -28.045 87.555 -27.715 87.885 ;
        RECT -28.045 86.195 -27.715 86.525 ;
        RECT -28.045 84.835 -27.715 85.165 ;
        RECT -28.045 83.475 -27.715 83.805 ;
        RECT -28.045 82.115 -27.715 82.445 ;
        RECT -28.045 80.755 -27.715 81.085 ;
        RECT -28.045 79.395 -27.715 79.725 ;
        RECT -28.045 78.035 -27.715 78.365 ;
        RECT -28.045 76.675 -27.715 77.005 ;
        RECT -28.045 75.315 -27.715 75.645 ;
        RECT -28.045 73.955 -27.715 74.285 ;
        RECT -28.045 72.595 -27.715 72.925 ;
        RECT -28.045 71.235 -27.715 71.565 ;
        RECT -28.045 69.875 -27.715 70.205 ;
        RECT -28.045 68.515 -27.715 68.845 ;
        RECT -28.045 67.155 -27.715 67.485 ;
        RECT -28.045 65.795 -27.715 66.125 ;
        RECT -28.045 64.435 -27.715 64.765 ;
        RECT -28.045 63.075 -27.715 63.405 ;
        RECT -28.045 61.715 -27.715 62.045 ;
        RECT -28.045 60.355 -27.715 60.685 ;
        RECT -28.045 58.995 -27.715 59.325 ;
        RECT -28.045 57.635 -27.715 57.965 ;
        RECT -28.045 56.275 -27.715 56.605 ;
        RECT -28.045 54.915 -27.715 55.245 ;
        RECT -28.045 53.555 -27.715 53.885 ;
        RECT -28.045 52.195 -27.715 52.525 ;
        RECT -28.045 50.835 -27.715 51.165 ;
        RECT -28.045 49.475 -27.715 49.805 ;
        RECT -28.045 48.115 -27.715 48.445 ;
        RECT -28.045 46.755 -27.715 47.085 ;
        RECT -28.045 45.395 -27.715 45.725 ;
        RECT -28.045 44.035 -27.715 44.365 ;
        RECT -28.045 42.675 -27.715 43.005 ;
        RECT -28.045 41.315 -27.715 41.645 ;
        RECT -28.045 39.955 -27.715 40.285 ;
        RECT -28.045 38.595 -27.715 38.925 ;
        RECT -28.045 37.235 -27.715 37.565 ;
        RECT -28.045 35.875 -27.715 36.205 ;
        RECT -28.045 34.515 -27.715 34.845 ;
        RECT -28.045 33.155 -27.715 33.485 ;
        RECT -28.045 31.795 -27.715 32.125 ;
        RECT -28.045 30.435 -27.715 30.765 ;
        RECT -28.045 29.075 -27.715 29.405 ;
        RECT -28.045 27.715 -27.715 28.045 ;
        RECT -28.045 26.355 -27.715 26.685 ;
        RECT -28.045 24.995 -27.715 25.325 ;
        RECT -28.045 23.635 -27.715 23.965 ;
        RECT -28.045 22.275 -27.715 22.605 ;
        RECT -28.045 20.915 -27.715 21.245 ;
        RECT -28.045 19.555 -27.715 19.885 ;
        RECT -28.045 18.195 -27.715 18.525 ;
        RECT -28.045 16.835 -27.715 17.165 ;
        RECT -28.045 15.475 -27.715 15.805 ;
        RECT -28.045 14.115 -27.715 14.445 ;
        RECT -28.045 12.755 -27.715 13.085 ;
        RECT -28.045 11.395 -27.715 11.725 ;
        RECT -28.045 10.035 -27.715 10.365 ;
        RECT -28.045 8.675 -27.715 9.005 ;
        RECT -28.045 7.315 -27.715 7.645 ;
        RECT -28.045 5.955 -27.715 6.285 ;
        RECT -28.045 4.595 -27.715 4.925 ;
        RECT -28.045 3.235 -27.715 3.565 ;
        RECT -28.045 1.875 -27.715 2.205 ;
        RECT -28.045 0.515 -27.715 0.845 ;
        RECT -28.045 -0.845 -27.715 -0.515 ;
        RECT -28.045 -7.645 -27.715 -7.315 ;
        RECT -28.045 -9.005 -27.715 -8.675 ;
        RECT -28.045 -10.73 -27.715 -10.4 ;
        RECT -28.045 -15.805 -27.715 -15.475 ;
        RECT -28.045 -16.77 -27.715 -16.44 ;
        RECT -28.045 -18.525 -27.715 -18.195 ;
        RECT -28.045 -21.245 -27.715 -20.915 ;
        RECT -28.045 -32.125 -27.715 -31.795 ;
        RECT -28.045 -33.71 -27.715 -33.38 ;
        RECT -28.045 -34.845 -27.715 -34.515 ;
        RECT -28.045 -36.205 -27.715 -35.875 ;
        RECT -28.045 -38.925 -27.715 -38.595 ;
        RECT -28.045 -39.75 -27.715 -39.42 ;
        RECT -28.045 -41.645 -27.715 -41.315 ;
        RECT -28.045 -44.365 -27.715 -44.035 ;
        RECT -28.045 -49.805 -27.715 -49.475 ;
        RECT -28.045 -51.165 -27.715 -50.835 ;
        RECT -28.045 -53.885 -27.715 -53.555 ;
        RECT -28.045 -55.245 -27.715 -54.915 ;
        RECT -28.045 -59.325 -27.715 -58.995 ;
        RECT -28.045 -60.685 -27.715 -60.355 ;
        RECT -28.045 -67.485 -27.715 -67.155 ;
        RECT -28.045 -68.845 -27.715 -68.515 ;
        RECT -28.045 -70.205 -27.715 -69.875 ;
        RECT -28.045 -71.565 -27.715 -71.235 ;
        RECT -28.045 -72.925 -27.715 -72.595 ;
        RECT -28.045 -74.285 -27.715 -73.955 ;
        RECT -28.045 -75.645 -27.715 -75.315 ;
        RECT -28.045 -77.005 -27.715 -76.675 ;
        RECT -28.045 -78.365 -27.715 -78.035 ;
        RECT -28.045 -79.725 -27.715 -79.395 ;
        RECT -28.045 -81.085 -27.715 -80.755 ;
        RECT -28.045 -82.445 -27.715 -82.115 ;
        RECT -28.045 -83.805 -27.715 -83.475 ;
        RECT -28.045 -85.165 -27.715 -84.835 ;
        RECT -28.045 -86.525 -27.715 -86.195 ;
        RECT -28.045 -87.885 -27.715 -87.555 ;
        RECT -28.045 -89.245 -27.715 -88.915 ;
        RECT -28.045 -90.81 -27.715 -90.48 ;
        RECT -28.045 -91.965 -27.715 -91.635 ;
        RECT -28.045 -93.325 -27.715 -92.995 ;
        RECT -28.045 -94.685 -27.715 -94.355 ;
        RECT -28.045 -96.045 -27.715 -95.715 ;
        RECT -28.045 -97.405 -27.715 -97.075 ;
        RECT -28.045 -100.125 -27.715 -99.795 ;
        RECT -28.045 -101.35 -27.715 -101.02 ;
        RECT -28.045 -102.845 -27.715 -102.515 ;
        RECT -28.045 -104.205 -27.715 -103.875 ;
        RECT -28.045 -105.565 -27.715 -105.235 ;
        RECT -28.045 -108.285 -27.715 -107.955 ;
        RECT -28.045 -109.645 -27.715 -109.315 ;
        RECT -28.045 -112.365 -27.715 -112.035 ;
        RECT -28.045 -113.725 -27.715 -113.395 ;
        RECT -28.045 -115.085 -27.715 -114.755 ;
        RECT -28.045 -116.445 -27.715 -116.115 ;
        RECT -28.045 -117.805 -27.715 -117.475 ;
        RECT -28.045 -119.165 -27.715 -118.835 ;
        RECT -28.045 -120.525 -27.715 -120.195 ;
        RECT -28.045 -121.885 -27.715 -121.555 ;
        RECT -28.045 -123.245 -27.715 -122.915 ;
        RECT -28.045 -125.965 -27.715 -125.635 ;
        RECT -28.045 -127.325 -27.715 -126.995 ;
        RECT -28.045 -128.685 -27.715 -128.355 ;
        RECT -28.045 -132.765 -27.715 -132.435 ;
        RECT -28.045 -134.125 -27.715 -133.795 ;
        RECT -28.045 -135.485 -27.715 -135.155 ;
        RECT -28.045 -136.845 -27.715 -136.515 ;
        RECT -28.045 -140.925 -27.715 -140.595 ;
        RECT -28.045 -142.285 -27.715 -141.955 ;
        RECT -28.045 -143.645 -27.715 -143.315 ;
        RECT -28.045 -145.005 -27.715 -144.675 ;
        RECT -28.045 -146.365 -27.715 -146.035 ;
        RECT -28.045 -147.725 -27.715 -147.395 ;
        RECT -28.045 -151.805 -27.715 -151.475 ;
        RECT -28.045 -155.885 -27.715 -155.555 ;
        RECT -28.045 -157.245 -27.715 -156.915 ;
        RECT -28.045 -158.605 -27.715 -158.275 ;
        RECT -28.045 -159.965 -27.715 -159.635 ;
        RECT -28.045 -161.325 -27.715 -160.995 ;
        RECT -28.045 -162.685 -27.715 -162.355 ;
        RECT -28.045 -164.045 -27.715 -163.715 ;
        RECT -28.045 -165.405 -27.715 -165.075 ;
        RECT -28.045 -166.765 -27.715 -166.435 ;
        RECT -28.045 -168.655 -27.715 -168.325 ;
        RECT -28.045 -169.485 -27.715 -169.155 ;
        RECT -28.045 -170.845 -27.715 -170.515 ;
        RECT -28.045 -172.205 -27.715 -171.875 ;
        RECT -28.04 -172.205 -27.72 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -26.685 141.955 -26.355 142.285 ;
        RECT -26.685 140.595 -26.355 140.925 ;
        RECT -26.685 139.235 -26.355 139.565 ;
        RECT -26.685 137.875 -26.355 138.205 ;
        RECT -26.685 136.515 -26.355 136.845 ;
        RECT -26.685 135.155 -26.355 135.485 ;
        RECT -26.685 133.795 -26.355 134.125 ;
        RECT -26.685 132.435 -26.355 132.765 ;
        RECT -26.685 131.075 -26.355 131.405 ;
        RECT -26.685 129.715 -26.355 130.045 ;
        RECT -26.685 128.355 -26.355 128.685 ;
        RECT -26.685 126.995 -26.355 127.325 ;
        RECT -26.685 125.635 -26.355 125.965 ;
        RECT -26.685 124.275 -26.355 124.605 ;
        RECT -26.685 122.915 -26.355 123.245 ;
        RECT -26.685 121.555 -26.355 121.885 ;
        RECT -26.685 120.195 -26.355 120.525 ;
        RECT -26.685 118.835 -26.355 119.165 ;
        RECT -26.685 117.475 -26.355 117.805 ;
        RECT -26.685 116.115 -26.355 116.445 ;
        RECT -26.685 114.755 -26.355 115.085 ;
        RECT -26.685 113.395 -26.355 113.725 ;
        RECT -26.685 112.035 -26.355 112.365 ;
        RECT -26.685 110.675 -26.355 111.005 ;
        RECT -26.685 109.315 -26.355 109.645 ;
        RECT -26.685 107.955 -26.355 108.285 ;
        RECT -26.685 106.595 -26.355 106.925 ;
        RECT -26.685 105.235 -26.355 105.565 ;
        RECT -26.685 103.875 -26.355 104.205 ;
        RECT -26.685 102.515 -26.355 102.845 ;
        RECT -26.685 101.155 -26.355 101.485 ;
        RECT -26.685 99.795 -26.355 100.125 ;
        RECT -26.685 98.435 -26.355 98.765 ;
        RECT -26.685 97.075 -26.355 97.405 ;
        RECT -26.685 95.715 -26.355 96.045 ;
        RECT -26.685 94.355 -26.355 94.685 ;
        RECT -26.685 92.995 -26.355 93.325 ;
        RECT -26.685 91.635 -26.355 91.965 ;
        RECT -26.685 90.275 -26.355 90.605 ;
        RECT -26.685 88.915 -26.355 89.245 ;
        RECT -26.685 87.555 -26.355 87.885 ;
        RECT -26.685 86.195 -26.355 86.525 ;
        RECT -26.685 84.835 -26.355 85.165 ;
        RECT -26.685 83.475 -26.355 83.805 ;
        RECT -26.685 82.115 -26.355 82.445 ;
        RECT -26.685 80.755 -26.355 81.085 ;
        RECT -26.685 79.395 -26.355 79.725 ;
        RECT -26.685 78.035 -26.355 78.365 ;
        RECT -26.685 76.675 -26.355 77.005 ;
        RECT -26.685 75.315 -26.355 75.645 ;
        RECT -26.685 73.955 -26.355 74.285 ;
        RECT -26.685 72.595 -26.355 72.925 ;
        RECT -26.685 71.235 -26.355 71.565 ;
        RECT -26.685 69.875 -26.355 70.205 ;
        RECT -26.685 68.515 -26.355 68.845 ;
        RECT -26.685 67.155 -26.355 67.485 ;
        RECT -26.685 65.795 -26.355 66.125 ;
        RECT -26.685 64.435 -26.355 64.765 ;
        RECT -26.685 63.075 -26.355 63.405 ;
        RECT -26.685 61.715 -26.355 62.045 ;
        RECT -26.685 60.355 -26.355 60.685 ;
        RECT -26.685 58.995 -26.355 59.325 ;
        RECT -26.685 57.635 -26.355 57.965 ;
        RECT -26.685 56.275 -26.355 56.605 ;
        RECT -26.685 54.915 -26.355 55.245 ;
        RECT -26.685 53.555 -26.355 53.885 ;
        RECT -26.685 52.195 -26.355 52.525 ;
        RECT -26.685 50.835 -26.355 51.165 ;
        RECT -26.685 49.475 -26.355 49.805 ;
        RECT -26.685 48.115 -26.355 48.445 ;
        RECT -26.685 46.755 -26.355 47.085 ;
        RECT -26.685 45.395 -26.355 45.725 ;
        RECT -26.685 44.035 -26.355 44.365 ;
        RECT -26.685 42.675 -26.355 43.005 ;
        RECT -26.685 41.315 -26.355 41.645 ;
        RECT -26.685 39.955 -26.355 40.285 ;
        RECT -26.685 38.595 -26.355 38.925 ;
        RECT -26.685 37.235 -26.355 37.565 ;
        RECT -26.685 35.875 -26.355 36.205 ;
        RECT -26.685 34.515 -26.355 34.845 ;
        RECT -26.685 33.155 -26.355 33.485 ;
        RECT -26.685 31.795 -26.355 32.125 ;
        RECT -26.685 30.435 -26.355 30.765 ;
        RECT -26.685 29.075 -26.355 29.405 ;
        RECT -26.685 27.715 -26.355 28.045 ;
        RECT -26.685 26.355 -26.355 26.685 ;
        RECT -26.685 24.995 -26.355 25.325 ;
        RECT -26.685 23.635 -26.355 23.965 ;
        RECT -26.685 22.275 -26.355 22.605 ;
        RECT -26.685 20.915 -26.355 21.245 ;
        RECT -26.685 19.555 -26.355 19.885 ;
        RECT -26.685 18.195 -26.355 18.525 ;
        RECT -26.685 16.835 -26.355 17.165 ;
        RECT -26.685 15.475 -26.355 15.805 ;
        RECT -26.685 14.115 -26.355 14.445 ;
        RECT -26.685 12.755 -26.355 13.085 ;
        RECT -26.685 11.395 -26.355 11.725 ;
        RECT -26.685 10.035 -26.355 10.365 ;
        RECT -26.685 8.675 -26.355 9.005 ;
        RECT -26.685 7.315 -26.355 7.645 ;
        RECT -26.685 5.955 -26.355 6.285 ;
        RECT -26.685 4.595 -26.355 4.925 ;
        RECT -26.685 3.235 -26.355 3.565 ;
        RECT -26.685 1.875 -26.355 2.205 ;
        RECT -26.685 0.515 -26.355 0.845 ;
        RECT -26.685 -0.845 -26.355 -0.515 ;
        RECT -26.685 -2.205 -26.355 -1.875 ;
        RECT -26.685 -7.645 -26.355 -7.315 ;
        RECT -26.685 -9.005 -26.355 -8.675 ;
        RECT -26.685 -10.73 -26.355 -10.4 ;
        RECT -26.685 -15.805 -26.355 -15.475 ;
        RECT -26.685 -16.77 -26.355 -16.44 ;
        RECT -26.685 -18.525 -26.355 -18.195 ;
        RECT -26.685 -21.245 -26.355 -20.915 ;
        RECT -26.685 -32.125 -26.355 -31.795 ;
        RECT -26.685 -33.71 -26.355 -33.38 ;
        RECT -26.685 -34.845 -26.355 -34.515 ;
        RECT -26.685 -36.205 -26.355 -35.875 ;
        RECT -26.685 -38.925 -26.355 -38.595 ;
        RECT -26.685 -39.75 -26.355 -39.42 ;
        RECT -26.685 -41.645 -26.355 -41.315 ;
        RECT -26.685 -44.365 -26.355 -44.035 ;
        RECT -26.685 -49.805 -26.355 -49.475 ;
        RECT -26.685 -51.165 -26.355 -50.835 ;
        RECT -26.685 -53.885 -26.355 -53.555 ;
        RECT -26.685 -55.245 -26.355 -54.915 ;
        RECT -26.685 -59.325 -26.355 -58.995 ;
        RECT -26.685 -60.685 -26.355 -60.355 ;
        RECT -26.685 -67.485 -26.355 -67.155 ;
        RECT -26.685 -68.845 -26.355 -68.515 ;
        RECT -26.685 -70.205 -26.355 -69.875 ;
        RECT -26.685 -71.565 -26.355 -71.235 ;
        RECT -26.685 -72.925 -26.355 -72.595 ;
        RECT -26.685 -74.285 -26.355 -73.955 ;
        RECT -26.685 -75.645 -26.355 -75.315 ;
        RECT -26.685 -77.005 -26.355 -76.675 ;
        RECT -26.685 -78.365 -26.355 -78.035 ;
        RECT -26.685 -79.725 -26.355 -79.395 ;
        RECT -26.685 -81.085 -26.355 -80.755 ;
        RECT -26.685 -82.445 -26.355 -82.115 ;
        RECT -26.685 -83.805 -26.355 -83.475 ;
        RECT -26.685 -85.165 -26.355 -84.835 ;
        RECT -26.685 -86.525 -26.355 -86.195 ;
        RECT -26.685 -87.885 -26.355 -87.555 ;
        RECT -26.685 -89.245 -26.355 -88.915 ;
        RECT -26.685 -91.965 -26.355 -91.635 ;
        RECT -26.685 -93.325 -26.355 -92.995 ;
        RECT -26.685 -94.685 -26.355 -94.355 ;
        RECT -26.685 -96.045 -26.355 -95.715 ;
        RECT -26.685 -97.405 -26.355 -97.075 ;
        RECT -26.685 -100.125 -26.355 -99.795 ;
        RECT -26.685 -102.845 -26.355 -102.515 ;
        RECT -26.685 -104.205 -26.355 -103.875 ;
        RECT -26.685 -105.565 -26.355 -105.235 ;
        RECT -26.685 -108.285 -26.355 -107.955 ;
        RECT -26.685 -109.645 -26.355 -109.315 ;
        RECT -26.685 -112.365 -26.355 -112.035 ;
        RECT -26.685 -113.725 -26.355 -113.395 ;
        RECT -26.685 -115.085 -26.355 -114.755 ;
        RECT -26.685 -116.445 -26.355 -116.115 ;
        RECT -26.685 -117.805 -26.355 -117.475 ;
        RECT -26.685 -119.165 -26.355 -118.835 ;
        RECT -26.685 -120.525 -26.355 -120.195 ;
        RECT -26.685 -121.885 -26.355 -121.555 ;
        RECT -26.685 -123.245 -26.355 -122.915 ;
        RECT -26.685 -125.965 -26.355 -125.635 ;
        RECT -26.685 -127.325 -26.355 -126.995 ;
        RECT -26.685 -128.685 -26.355 -128.355 ;
        RECT -26.685 -132.765 -26.355 -132.435 ;
        RECT -26.685 -134.125 -26.355 -133.795 ;
        RECT -26.685 -135.485 -26.355 -135.155 ;
        RECT -26.685 -136.845 -26.355 -136.515 ;
        RECT -26.685 -140.925 -26.355 -140.595 ;
        RECT -26.685 -142.285 -26.355 -141.955 ;
        RECT -26.685 -143.645 -26.355 -143.315 ;
        RECT -26.685 -145.005 -26.355 -144.675 ;
        RECT -26.685 -146.365 -26.355 -146.035 ;
        RECT -26.685 -147.725 -26.355 -147.395 ;
        RECT -26.685 -151.805 -26.355 -151.475 ;
        RECT -26.685 -155.885 -26.355 -155.555 ;
        RECT -26.685 -157.245 -26.355 -156.915 ;
        RECT -26.685 -158.605 -26.355 -158.275 ;
        RECT -26.685 -159.965 -26.355 -159.635 ;
        RECT -26.685 -161.325 -26.355 -160.995 ;
        RECT -26.685 -162.685 -26.355 -162.355 ;
        RECT -26.685 -164.045 -26.355 -163.715 ;
        RECT -26.685 -165.405 -26.355 -165.075 ;
        RECT -26.685 -166.765 -26.355 -166.435 ;
        RECT -26.685 -168.655 -26.355 -168.325 ;
        RECT -26.685 -169.485 -26.355 -169.155 ;
        RECT -26.685 -170.845 -26.355 -170.515 ;
        RECT -26.685 -173.565 -26.355 -173.235 ;
        RECT -26.685 -174.925 -26.355 -174.595 ;
        RECT -26.685 -177.645 -26.355 -177.315 ;
        RECT -26.685 -183.29 -26.355 -182.16 ;
        RECT -26.68 -183.405 -26.36 245.285 ;
        RECT -26.685 244.04 -26.355 245.17 ;
        RECT -26.685 239.875 -26.355 240.205 ;
        RECT -26.685 238.515 -26.355 238.845 ;
        RECT -26.685 237.155 -26.355 237.485 ;
        RECT -26.685 235.795 -26.355 236.125 ;
        RECT -26.685 234.435 -26.355 234.765 ;
        RECT -26.685 233.075 -26.355 233.405 ;
        RECT -26.685 231.715 -26.355 232.045 ;
        RECT -26.685 230.355 -26.355 230.685 ;
        RECT -26.685 228.995 -26.355 229.325 ;
        RECT -26.685 227.635 -26.355 227.965 ;
        RECT -26.685 226.275 -26.355 226.605 ;
        RECT -26.685 224.915 -26.355 225.245 ;
        RECT -26.685 223.555 -26.355 223.885 ;
        RECT -26.685 222.195 -26.355 222.525 ;
        RECT -26.685 220.835 -26.355 221.165 ;
        RECT -26.685 219.475 -26.355 219.805 ;
        RECT -26.685 218.115 -26.355 218.445 ;
        RECT -26.685 216.755 -26.355 217.085 ;
        RECT -26.685 215.395 -26.355 215.725 ;
        RECT -26.685 214.035 -26.355 214.365 ;
        RECT -26.685 212.675 -26.355 213.005 ;
        RECT -26.685 211.315 -26.355 211.645 ;
        RECT -26.685 209.955 -26.355 210.285 ;
        RECT -26.685 208.595 -26.355 208.925 ;
        RECT -26.685 207.235 -26.355 207.565 ;
        RECT -26.685 205.875 -26.355 206.205 ;
        RECT -26.685 204.515 -26.355 204.845 ;
        RECT -26.685 203.155 -26.355 203.485 ;
        RECT -26.685 201.795 -26.355 202.125 ;
        RECT -26.685 200.435 -26.355 200.765 ;
        RECT -26.685 199.075 -26.355 199.405 ;
        RECT -26.685 197.715 -26.355 198.045 ;
        RECT -26.685 196.355 -26.355 196.685 ;
        RECT -26.685 194.995 -26.355 195.325 ;
        RECT -26.685 193.635 -26.355 193.965 ;
        RECT -26.685 192.275 -26.355 192.605 ;
        RECT -26.685 190.915 -26.355 191.245 ;
        RECT -26.685 189.555 -26.355 189.885 ;
        RECT -26.685 188.195 -26.355 188.525 ;
        RECT -26.685 186.835 -26.355 187.165 ;
        RECT -26.685 185.475 -26.355 185.805 ;
        RECT -26.685 184.115 -26.355 184.445 ;
        RECT -26.685 182.755 -26.355 183.085 ;
        RECT -26.685 181.395 -26.355 181.725 ;
        RECT -26.685 180.035 -26.355 180.365 ;
        RECT -26.685 178.675 -26.355 179.005 ;
        RECT -26.685 177.315 -26.355 177.645 ;
        RECT -26.685 175.955 -26.355 176.285 ;
        RECT -26.685 174.595 -26.355 174.925 ;
        RECT -26.685 173.235 -26.355 173.565 ;
        RECT -26.685 171.875 -26.355 172.205 ;
        RECT -26.685 170.515 -26.355 170.845 ;
        RECT -26.685 169.155 -26.355 169.485 ;
        RECT -26.685 167.795 -26.355 168.125 ;
        RECT -26.685 166.435 -26.355 166.765 ;
        RECT -26.685 165.075 -26.355 165.405 ;
        RECT -26.685 163.715 -26.355 164.045 ;
        RECT -26.685 162.355 -26.355 162.685 ;
        RECT -26.685 160.995 -26.355 161.325 ;
        RECT -26.685 159.635 -26.355 159.965 ;
        RECT -26.685 158.275 -26.355 158.605 ;
        RECT -26.685 156.915 -26.355 157.245 ;
        RECT -26.685 155.555 -26.355 155.885 ;
        RECT -26.685 154.195 -26.355 154.525 ;
        RECT -26.685 152.835 -26.355 153.165 ;
        RECT -26.685 151.475 -26.355 151.805 ;
        RECT -26.685 150.115 -26.355 150.445 ;
        RECT -26.685 148.755 -26.355 149.085 ;
        RECT -26.685 147.395 -26.355 147.725 ;
        RECT -26.685 146.035 -26.355 146.365 ;
        RECT -26.685 144.675 -26.355 145.005 ;
        RECT -26.685 143.315 -26.355 143.645 ;
    END
    PORT
      LAYER met3 ;
        RECT -34.845 244.04 -34.515 245.17 ;
        RECT -34.845 239.875 -34.515 240.205 ;
        RECT -34.845 238.515 -34.515 238.845 ;
        RECT -34.845 237.155 -34.515 237.485 ;
        RECT -34.845 235.795 -34.515 236.125 ;
        RECT -34.845 234.435 -34.515 234.765 ;
        RECT -34.845 233.075 -34.515 233.405 ;
        RECT -34.845 231.715 -34.515 232.045 ;
        RECT -34.845 230.355 -34.515 230.685 ;
        RECT -34.845 228.995 -34.515 229.325 ;
        RECT -34.845 227.635 -34.515 227.965 ;
        RECT -34.845 226.275 -34.515 226.605 ;
        RECT -34.845 224.915 -34.515 225.245 ;
        RECT -34.845 223.555 -34.515 223.885 ;
        RECT -34.845 222.195 -34.515 222.525 ;
        RECT -34.845 220.835 -34.515 221.165 ;
        RECT -34.845 219.475 -34.515 219.805 ;
        RECT -34.845 218.115 -34.515 218.445 ;
        RECT -34.845 216.755 -34.515 217.085 ;
        RECT -34.845 215.395 -34.515 215.725 ;
        RECT -34.845 214.035 -34.515 214.365 ;
        RECT -34.845 212.675 -34.515 213.005 ;
        RECT -34.845 211.315 -34.515 211.645 ;
        RECT -34.845 209.955 -34.515 210.285 ;
        RECT -34.845 208.595 -34.515 208.925 ;
        RECT -34.845 207.235 -34.515 207.565 ;
        RECT -34.845 205.875 -34.515 206.205 ;
        RECT -34.845 204.515 -34.515 204.845 ;
        RECT -34.845 203.155 -34.515 203.485 ;
        RECT -34.845 201.795 -34.515 202.125 ;
        RECT -34.845 200.435 -34.515 200.765 ;
        RECT -34.845 199.075 -34.515 199.405 ;
        RECT -34.845 197.715 -34.515 198.045 ;
        RECT -34.845 196.355 -34.515 196.685 ;
        RECT -34.845 194.995 -34.515 195.325 ;
        RECT -34.845 193.635 -34.515 193.965 ;
        RECT -34.845 192.275 -34.515 192.605 ;
        RECT -34.845 190.915 -34.515 191.245 ;
        RECT -34.845 189.555 -34.515 189.885 ;
        RECT -34.845 188.195 -34.515 188.525 ;
        RECT -34.845 186.835 -34.515 187.165 ;
        RECT -34.845 185.475 -34.515 185.805 ;
        RECT -34.845 184.115 -34.515 184.445 ;
        RECT -34.845 182.755 -34.515 183.085 ;
        RECT -34.845 181.395 -34.515 181.725 ;
        RECT -34.845 180.035 -34.515 180.365 ;
        RECT -34.845 178.675 -34.515 179.005 ;
        RECT -34.845 177.315 -34.515 177.645 ;
        RECT -34.845 175.955 -34.515 176.285 ;
        RECT -34.845 174.595 -34.515 174.925 ;
        RECT -34.845 173.235 -34.515 173.565 ;
        RECT -34.845 171.875 -34.515 172.205 ;
        RECT -34.845 170.515 -34.515 170.845 ;
        RECT -34.845 169.155 -34.515 169.485 ;
        RECT -34.845 167.795 -34.515 168.125 ;
        RECT -34.845 166.435 -34.515 166.765 ;
        RECT -34.845 165.075 -34.515 165.405 ;
        RECT -34.845 163.715 -34.515 164.045 ;
        RECT -34.845 162.355 -34.515 162.685 ;
        RECT -34.845 160.995 -34.515 161.325 ;
        RECT -34.845 159.635 -34.515 159.965 ;
        RECT -34.845 158.275 -34.515 158.605 ;
        RECT -34.845 156.915 -34.515 157.245 ;
        RECT -34.845 155.555 -34.515 155.885 ;
        RECT -34.845 154.195 -34.515 154.525 ;
        RECT -34.845 152.835 -34.515 153.165 ;
        RECT -34.845 151.475 -34.515 151.805 ;
        RECT -34.845 150.115 -34.515 150.445 ;
        RECT -34.845 148.755 -34.515 149.085 ;
        RECT -34.845 147.395 -34.515 147.725 ;
        RECT -34.845 146.035 -34.515 146.365 ;
        RECT -34.845 144.675 -34.515 145.005 ;
        RECT -34.845 143.315 -34.515 143.645 ;
        RECT -34.845 141.955 -34.515 142.285 ;
        RECT -34.845 140.595 -34.515 140.925 ;
        RECT -34.845 139.235 -34.515 139.565 ;
        RECT -34.845 137.875 -34.515 138.205 ;
        RECT -34.845 136.515 -34.515 136.845 ;
        RECT -34.845 135.155 -34.515 135.485 ;
        RECT -34.845 133.795 -34.515 134.125 ;
        RECT -34.845 132.435 -34.515 132.765 ;
        RECT -34.845 131.075 -34.515 131.405 ;
        RECT -34.845 129.715 -34.515 130.045 ;
        RECT -34.845 128.355 -34.515 128.685 ;
        RECT -34.845 126.995 -34.515 127.325 ;
        RECT -34.845 125.635 -34.515 125.965 ;
        RECT -34.845 124.275 -34.515 124.605 ;
        RECT -34.845 122.915 -34.515 123.245 ;
        RECT -34.845 121.555 -34.515 121.885 ;
        RECT -34.845 120.195 -34.515 120.525 ;
        RECT -34.845 118.835 -34.515 119.165 ;
        RECT -34.845 117.475 -34.515 117.805 ;
        RECT -34.845 116.115 -34.515 116.445 ;
        RECT -34.845 114.755 -34.515 115.085 ;
        RECT -34.845 113.395 -34.515 113.725 ;
        RECT -34.845 112.035 -34.515 112.365 ;
        RECT -34.845 110.675 -34.515 111.005 ;
        RECT -34.845 109.315 -34.515 109.645 ;
        RECT -34.845 107.955 -34.515 108.285 ;
        RECT -34.845 106.595 -34.515 106.925 ;
        RECT -34.845 105.235 -34.515 105.565 ;
        RECT -34.845 103.875 -34.515 104.205 ;
        RECT -34.845 102.515 -34.515 102.845 ;
        RECT -34.845 101.155 -34.515 101.485 ;
        RECT -34.845 99.795 -34.515 100.125 ;
        RECT -34.845 98.435 -34.515 98.765 ;
        RECT -34.845 97.075 -34.515 97.405 ;
        RECT -34.845 95.715 -34.515 96.045 ;
        RECT -34.845 94.355 -34.515 94.685 ;
        RECT -34.845 92.995 -34.515 93.325 ;
        RECT -34.845 91.635 -34.515 91.965 ;
        RECT -34.845 90.275 -34.515 90.605 ;
        RECT -34.845 88.915 -34.515 89.245 ;
        RECT -34.845 87.555 -34.515 87.885 ;
        RECT -34.845 86.195 -34.515 86.525 ;
        RECT -34.845 84.835 -34.515 85.165 ;
        RECT -34.845 83.475 -34.515 83.805 ;
        RECT -34.845 82.115 -34.515 82.445 ;
        RECT -34.845 80.755 -34.515 81.085 ;
        RECT -34.845 79.395 -34.515 79.725 ;
        RECT -34.845 78.035 -34.515 78.365 ;
        RECT -34.845 76.675 -34.515 77.005 ;
        RECT -34.845 75.315 -34.515 75.645 ;
        RECT -34.845 73.955 -34.515 74.285 ;
        RECT -34.845 72.595 -34.515 72.925 ;
        RECT -34.845 71.235 -34.515 71.565 ;
        RECT -34.845 69.875 -34.515 70.205 ;
        RECT -34.845 68.515 -34.515 68.845 ;
        RECT -34.845 67.155 -34.515 67.485 ;
        RECT -34.845 65.795 -34.515 66.125 ;
        RECT -34.845 64.435 -34.515 64.765 ;
        RECT -34.845 63.075 -34.515 63.405 ;
        RECT -34.845 61.715 -34.515 62.045 ;
        RECT -34.845 60.355 -34.515 60.685 ;
        RECT -34.845 58.995 -34.515 59.325 ;
        RECT -34.845 57.635 -34.515 57.965 ;
        RECT -34.845 56.275 -34.515 56.605 ;
        RECT -34.845 54.915 -34.515 55.245 ;
        RECT -34.845 53.555 -34.515 53.885 ;
        RECT -34.845 52.195 -34.515 52.525 ;
        RECT -34.845 50.835 -34.515 51.165 ;
        RECT -34.845 49.475 -34.515 49.805 ;
        RECT -34.845 48.115 -34.515 48.445 ;
        RECT -34.845 46.755 -34.515 47.085 ;
        RECT -34.845 45.395 -34.515 45.725 ;
        RECT -34.845 44.035 -34.515 44.365 ;
        RECT -34.845 42.675 -34.515 43.005 ;
        RECT -34.845 41.315 -34.515 41.645 ;
        RECT -34.845 39.955 -34.515 40.285 ;
        RECT -34.845 38.595 -34.515 38.925 ;
        RECT -34.845 37.235 -34.515 37.565 ;
        RECT -34.845 35.875 -34.515 36.205 ;
        RECT -34.845 34.515 -34.515 34.845 ;
        RECT -34.845 33.155 -34.515 33.485 ;
        RECT -34.845 31.795 -34.515 32.125 ;
        RECT -34.845 30.435 -34.515 30.765 ;
        RECT -34.845 29.075 -34.515 29.405 ;
        RECT -34.845 27.715 -34.515 28.045 ;
        RECT -34.845 26.355 -34.515 26.685 ;
        RECT -34.845 24.995 -34.515 25.325 ;
        RECT -34.845 23.635 -34.515 23.965 ;
        RECT -34.845 22.275 -34.515 22.605 ;
        RECT -34.845 20.915 -34.515 21.245 ;
        RECT -34.845 19.555 -34.515 19.885 ;
        RECT -34.845 18.195 -34.515 18.525 ;
        RECT -34.845 16.835 -34.515 17.165 ;
        RECT -34.845 15.475 -34.515 15.805 ;
        RECT -34.845 14.115 -34.515 14.445 ;
        RECT -34.845 12.755 -34.515 13.085 ;
        RECT -34.845 11.395 -34.515 11.725 ;
        RECT -34.845 10.035 -34.515 10.365 ;
        RECT -34.845 8.675 -34.515 9.005 ;
        RECT -34.845 7.315 -34.515 7.645 ;
        RECT -34.845 5.955 -34.515 6.285 ;
        RECT -34.845 4.595 -34.515 4.925 ;
        RECT -34.845 3.235 -34.515 3.565 ;
        RECT -34.845 1.875 -34.515 2.205 ;
        RECT -34.845 0.515 -34.515 0.845 ;
        RECT -34.845 -0.845 -34.515 -0.515 ;
        RECT -34.845 -7.645 -34.515 -7.315 ;
        RECT -34.845 -10.365 -34.515 -10.035 ;
        RECT -34.845 -14.445 -34.515 -14.115 ;
        RECT -34.845 -15.805 -34.515 -15.475 ;
        RECT -34.845 -17.165 -34.515 -16.835 ;
        RECT -34.845 -18.525 -34.515 -18.195 ;
        RECT -34.845 -19.885 -34.515 -19.555 ;
        RECT -34.845 -21.245 -34.515 -20.915 ;
        RECT -34.845 -22.605 -34.515 -22.275 ;
        RECT -34.845 -23.965 -34.515 -23.635 ;
        RECT -34.845 -25.325 -34.515 -24.995 ;
        RECT -34.845 -32.125 -34.515 -31.795 ;
        RECT -34.845 -33.71 -34.515 -33.38 ;
        RECT -34.845 -34.845 -34.515 -34.515 ;
        RECT -34.845 -36.205 -34.515 -35.875 ;
        RECT -34.845 -38.925 -34.515 -38.595 ;
        RECT -34.845 -39.75 -34.515 -39.42 ;
        RECT -34.845 -41.645 -34.515 -41.315 ;
        RECT -34.845 -44.365 -34.515 -44.035 ;
        RECT -34.845 -49.805 -34.515 -49.475 ;
        RECT -34.845 -51.165 -34.515 -50.835 ;
        RECT -34.845 -53.885 -34.515 -53.555 ;
        RECT -34.845 -55.245 -34.515 -54.915 ;
        RECT -34.845 -59.325 -34.515 -58.995 ;
        RECT -34.845 -60.685 -34.515 -60.355 ;
        RECT -34.845 -67.485 -34.515 -67.155 ;
        RECT -34.845 -68.845 -34.515 -68.515 ;
        RECT -34.845 -70.205 -34.515 -69.875 ;
        RECT -34.845 -71.565 -34.515 -71.235 ;
        RECT -34.845 -72.925 -34.515 -72.595 ;
        RECT -34.845 -74.285 -34.515 -73.955 ;
        RECT -34.845 -75.645 -34.515 -75.315 ;
        RECT -34.845 -77.005 -34.515 -76.675 ;
        RECT -34.845 -78.365 -34.515 -78.035 ;
        RECT -34.845 -79.725 -34.515 -79.395 ;
        RECT -34.845 -81.085 -34.515 -80.755 ;
        RECT -34.845 -82.445 -34.515 -82.115 ;
        RECT -34.845 -83.805 -34.515 -83.475 ;
        RECT -34.845 -85.165 -34.515 -84.835 ;
        RECT -34.845 -86.525 -34.515 -86.195 ;
        RECT -34.845 -87.885 -34.515 -87.555 ;
        RECT -34.845 -89.245 -34.515 -88.915 ;
        RECT -34.845 -90.81 -34.515 -90.48 ;
        RECT -34.845 -91.965 -34.515 -91.635 ;
        RECT -34.845 -93.325 -34.515 -92.995 ;
        RECT -34.845 -94.685 -34.515 -94.355 ;
        RECT -34.845 -96.045 -34.515 -95.715 ;
        RECT -34.845 -97.405 -34.515 -97.075 ;
        RECT -34.845 -100.125 -34.515 -99.795 ;
        RECT -34.845 -101.35 -34.515 -101.02 ;
        RECT -34.845 -102.845 -34.515 -102.515 ;
        RECT -34.845 -104.205 -34.515 -103.875 ;
        RECT -34.845 -105.565 -34.515 -105.235 ;
        RECT -34.845 -108.285 -34.515 -107.955 ;
        RECT -34.845 -109.645 -34.515 -109.315 ;
        RECT -34.84 -112.36 -34.52 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -34.845 -174.925 -34.515 -174.595 ;
        RECT -34.845 -177.645 -34.515 -177.315 ;
        RECT -34.845 -183.29 -34.515 -182.16 ;
        RECT -34.84 -183.405 -34.52 -173.92 ;
    END
    PORT
      LAYER met3 ;
        RECT -33.485 244.04 -33.155 245.17 ;
        RECT -33.485 239.875 -33.155 240.205 ;
        RECT -33.485 238.515 -33.155 238.845 ;
        RECT -33.485 237.155 -33.155 237.485 ;
        RECT -33.485 235.795 -33.155 236.125 ;
        RECT -33.485 234.435 -33.155 234.765 ;
        RECT -33.485 233.075 -33.155 233.405 ;
        RECT -33.485 231.715 -33.155 232.045 ;
        RECT -33.485 230.355 -33.155 230.685 ;
        RECT -33.485 228.995 -33.155 229.325 ;
        RECT -33.485 227.635 -33.155 227.965 ;
        RECT -33.485 226.275 -33.155 226.605 ;
        RECT -33.485 224.915 -33.155 225.245 ;
        RECT -33.485 223.555 -33.155 223.885 ;
        RECT -33.485 222.195 -33.155 222.525 ;
        RECT -33.485 220.835 -33.155 221.165 ;
        RECT -33.485 219.475 -33.155 219.805 ;
        RECT -33.485 218.115 -33.155 218.445 ;
        RECT -33.485 216.755 -33.155 217.085 ;
        RECT -33.485 215.395 -33.155 215.725 ;
        RECT -33.485 214.035 -33.155 214.365 ;
        RECT -33.485 212.675 -33.155 213.005 ;
        RECT -33.485 211.315 -33.155 211.645 ;
        RECT -33.485 209.955 -33.155 210.285 ;
        RECT -33.485 208.595 -33.155 208.925 ;
        RECT -33.485 207.235 -33.155 207.565 ;
        RECT -33.485 205.875 -33.155 206.205 ;
        RECT -33.485 204.515 -33.155 204.845 ;
        RECT -33.485 203.155 -33.155 203.485 ;
        RECT -33.485 201.795 -33.155 202.125 ;
        RECT -33.485 200.435 -33.155 200.765 ;
        RECT -33.485 199.075 -33.155 199.405 ;
        RECT -33.485 197.715 -33.155 198.045 ;
        RECT -33.485 196.355 -33.155 196.685 ;
        RECT -33.485 194.995 -33.155 195.325 ;
        RECT -33.485 193.635 -33.155 193.965 ;
        RECT -33.485 192.275 -33.155 192.605 ;
        RECT -33.485 190.915 -33.155 191.245 ;
        RECT -33.485 189.555 -33.155 189.885 ;
        RECT -33.485 188.195 -33.155 188.525 ;
        RECT -33.485 186.835 -33.155 187.165 ;
        RECT -33.485 185.475 -33.155 185.805 ;
        RECT -33.485 184.115 -33.155 184.445 ;
        RECT -33.485 182.755 -33.155 183.085 ;
        RECT -33.485 181.395 -33.155 181.725 ;
        RECT -33.485 180.035 -33.155 180.365 ;
        RECT -33.485 178.675 -33.155 179.005 ;
        RECT -33.485 177.315 -33.155 177.645 ;
        RECT -33.485 175.955 -33.155 176.285 ;
        RECT -33.485 174.595 -33.155 174.925 ;
        RECT -33.485 173.235 -33.155 173.565 ;
        RECT -33.485 171.875 -33.155 172.205 ;
        RECT -33.485 170.515 -33.155 170.845 ;
        RECT -33.485 169.155 -33.155 169.485 ;
        RECT -33.485 167.795 -33.155 168.125 ;
        RECT -33.485 166.435 -33.155 166.765 ;
        RECT -33.485 165.075 -33.155 165.405 ;
        RECT -33.485 163.715 -33.155 164.045 ;
        RECT -33.485 162.355 -33.155 162.685 ;
        RECT -33.485 160.995 -33.155 161.325 ;
        RECT -33.485 159.635 -33.155 159.965 ;
        RECT -33.485 158.275 -33.155 158.605 ;
        RECT -33.485 156.915 -33.155 157.245 ;
        RECT -33.485 155.555 -33.155 155.885 ;
        RECT -33.485 154.195 -33.155 154.525 ;
        RECT -33.485 152.835 -33.155 153.165 ;
        RECT -33.485 151.475 -33.155 151.805 ;
        RECT -33.485 150.115 -33.155 150.445 ;
        RECT -33.485 148.755 -33.155 149.085 ;
        RECT -33.485 147.395 -33.155 147.725 ;
        RECT -33.485 146.035 -33.155 146.365 ;
        RECT -33.485 144.675 -33.155 145.005 ;
        RECT -33.485 143.315 -33.155 143.645 ;
        RECT -33.485 141.955 -33.155 142.285 ;
        RECT -33.485 140.595 -33.155 140.925 ;
        RECT -33.485 139.235 -33.155 139.565 ;
        RECT -33.485 137.875 -33.155 138.205 ;
        RECT -33.485 136.515 -33.155 136.845 ;
        RECT -33.485 135.155 -33.155 135.485 ;
        RECT -33.485 133.795 -33.155 134.125 ;
        RECT -33.485 132.435 -33.155 132.765 ;
        RECT -33.485 131.075 -33.155 131.405 ;
        RECT -33.485 129.715 -33.155 130.045 ;
        RECT -33.485 128.355 -33.155 128.685 ;
        RECT -33.485 126.995 -33.155 127.325 ;
        RECT -33.485 125.635 -33.155 125.965 ;
        RECT -33.485 124.275 -33.155 124.605 ;
        RECT -33.485 122.915 -33.155 123.245 ;
        RECT -33.485 121.555 -33.155 121.885 ;
        RECT -33.485 120.195 -33.155 120.525 ;
        RECT -33.485 118.835 -33.155 119.165 ;
        RECT -33.485 117.475 -33.155 117.805 ;
        RECT -33.485 116.115 -33.155 116.445 ;
        RECT -33.485 114.755 -33.155 115.085 ;
        RECT -33.485 113.395 -33.155 113.725 ;
        RECT -33.485 112.035 -33.155 112.365 ;
        RECT -33.485 110.675 -33.155 111.005 ;
        RECT -33.485 109.315 -33.155 109.645 ;
        RECT -33.485 107.955 -33.155 108.285 ;
        RECT -33.485 106.595 -33.155 106.925 ;
        RECT -33.485 105.235 -33.155 105.565 ;
        RECT -33.485 103.875 -33.155 104.205 ;
        RECT -33.485 102.515 -33.155 102.845 ;
        RECT -33.485 101.155 -33.155 101.485 ;
        RECT -33.485 99.795 -33.155 100.125 ;
        RECT -33.485 98.435 -33.155 98.765 ;
        RECT -33.485 97.075 -33.155 97.405 ;
        RECT -33.485 95.715 -33.155 96.045 ;
        RECT -33.485 94.355 -33.155 94.685 ;
        RECT -33.485 92.995 -33.155 93.325 ;
        RECT -33.485 91.635 -33.155 91.965 ;
        RECT -33.485 90.275 -33.155 90.605 ;
        RECT -33.485 88.915 -33.155 89.245 ;
        RECT -33.485 87.555 -33.155 87.885 ;
        RECT -33.485 86.195 -33.155 86.525 ;
        RECT -33.485 84.835 -33.155 85.165 ;
        RECT -33.485 83.475 -33.155 83.805 ;
        RECT -33.485 82.115 -33.155 82.445 ;
        RECT -33.485 80.755 -33.155 81.085 ;
        RECT -33.485 79.395 -33.155 79.725 ;
        RECT -33.485 78.035 -33.155 78.365 ;
        RECT -33.485 76.675 -33.155 77.005 ;
        RECT -33.485 75.315 -33.155 75.645 ;
        RECT -33.485 73.955 -33.155 74.285 ;
        RECT -33.485 72.595 -33.155 72.925 ;
        RECT -33.485 71.235 -33.155 71.565 ;
        RECT -33.485 69.875 -33.155 70.205 ;
        RECT -33.485 68.515 -33.155 68.845 ;
        RECT -33.485 67.155 -33.155 67.485 ;
        RECT -33.485 65.795 -33.155 66.125 ;
        RECT -33.485 64.435 -33.155 64.765 ;
        RECT -33.485 63.075 -33.155 63.405 ;
        RECT -33.485 61.715 -33.155 62.045 ;
        RECT -33.485 60.355 -33.155 60.685 ;
        RECT -33.485 58.995 -33.155 59.325 ;
        RECT -33.485 57.635 -33.155 57.965 ;
        RECT -33.485 56.275 -33.155 56.605 ;
        RECT -33.485 54.915 -33.155 55.245 ;
        RECT -33.485 53.555 -33.155 53.885 ;
        RECT -33.485 52.195 -33.155 52.525 ;
        RECT -33.485 50.835 -33.155 51.165 ;
        RECT -33.485 49.475 -33.155 49.805 ;
        RECT -33.485 48.115 -33.155 48.445 ;
        RECT -33.485 46.755 -33.155 47.085 ;
        RECT -33.485 45.395 -33.155 45.725 ;
        RECT -33.485 44.035 -33.155 44.365 ;
        RECT -33.485 42.675 -33.155 43.005 ;
        RECT -33.485 41.315 -33.155 41.645 ;
        RECT -33.485 39.955 -33.155 40.285 ;
        RECT -33.485 38.595 -33.155 38.925 ;
        RECT -33.485 37.235 -33.155 37.565 ;
        RECT -33.485 35.875 -33.155 36.205 ;
        RECT -33.485 34.515 -33.155 34.845 ;
        RECT -33.485 33.155 -33.155 33.485 ;
        RECT -33.485 31.795 -33.155 32.125 ;
        RECT -33.485 30.435 -33.155 30.765 ;
        RECT -33.485 29.075 -33.155 29.405 ;
        RECT -33.485 27.715 -33.155 28.045 ;
        RECT -33.485 26.355 -33.155 26.685 ;
        RECT -33.485 24.995 -33.155 25.325 ;
        RECT -33.485 23.635 -33.155 23.965 ;
        RECT -33.485 22.275 -33.155 22.605 ;
        RECT -33.485 20.915 -33.155 21.245 ;
        RECT -33.485 19.555 -33.155 19.885 ;
        RECT -33.485 18.195 -33.155 18.525 ;
        RECT -33.485 16.835 -33.155 17.165 ;
        RECT -33.485 15.475 -33.155 15.805 ;
        RECT -33.485 14.115 -33.155 14.445 ;
        RECT -33.485 12.755 -33.155 13.085 ;
        RECT -33.485 11.395 -33.155 11.725 ;
        RECT -33.485 10.035 -33.155 10.365 ;
        RECT -33.485 8.675 -33.155 9.005 ;
        RECT -33.485 7.315 -33.155 7.645 ;
        RECT -33.485 5.955 -33.155 6.285 ;
        RECT -33.485 4.595 -33.155 4.925 ;
        RECT -33.485 3.235 -33.155 3.565 ;
        RECT -33.485 1.875 -33.155 2.205 ;
        RECT -33.485 0.515 -33.155 0.845 ;
        RECT -33.485 -0.845 -33.155 -0.515 ;
        RECT -33.485 -7.645 -33.155 -7.315 ;
        RECT -33.485 -10.365 -33.155 -10.035 ;
        RECT -33.485 -14.445 -33.155 -14.115 ;
        RECT -33.485 -15.805 -33.155 -15.475 ;
        RECT -33.485 -17.165 -33.155 -16.835 ;
        RECT -33.485 -18.525 -33.155 -18.195 ;
        RECT -33.485 -19.885 -33.155 -19.555 ;
        RECT -33.485 -21.245 -33.155 -20.915 ;
        RECT -33.485 -22.605 -33.155 -22.275 ;
        RECT -33.485 -23.965 -33.155 -23.635 ;
        RECT -33.485 -25.325 -33.155 -24.995 ;
        RECT -33.485 -32.125 -33.155 -31.795 ;
        RECT -33.485 -33.71 -33.155 -33.38 ;
        RECT -33.485 -34.845 -33.155 -34.515 ;
        RECT -33.485 -36.205 -33.155 -35.875 ;
        RECT -33.485 -38.925 -33.155 -38.595 ;
        RECT -33.485 -39.75 -33.155 -39.42 ;
        RECT -33.485 -41.645 -33.155 -41.315 ;
        RECT -33.485 -44.365 -33.155 -44.035 ;
        RECT -33.485 -49.805 -33.155 -49.475 ;
        RECT -33.485 -51.165 -33.155 -50.835 ;
        RECT -33.485 -53.885 -33.155 -53.555 ;
        RECT -33.485 -55.245 -33.155 -54.915 ;
        RECT -33.485 -59.325 -33.155 -58.995 ;
        RECT -33.485 -60.685 -33.155 -60.355 ;
        RECT -33.485 -68.845 -33.155 -68.515 ;
        RECT -33.485 -70.205 -33.155 -69.875 ;
        RECT -33.485 -71.565 -33.155 -71.235 ;
        RECT -33.485 -72.925 -33.155 -72.595 ;
        RECT -33.485 -74.285 -33.155 -73.955 ;
        RECT -33.485 -75.645 -33.155 -75.315 ;
        RECT -33.485 -77.005 -33.155 -76.675 ;
        RECT -33.485 -78.365 -33.155 -78.035 ;
        RECT -33.485 -79.725 -33.155 -79.395 ;
        RECT -33.485 -81.085 -33.155 -80.755 ;
        RECT -33.485 -82.445 -33.155 -82.115 ;
        RECT -33.485 -83.805 -33.155 -83.475 ;
        RECT -33.485 -85.165 -33.155 -84.835 ;
        RECT -33.485 -86.525 -33.155 -86.195 ;
        RECT -33.485 -87.885 -33.155 -87.555 ;
        RECT -33.485 -89.245 -33.155 -88.915 ;
        RECT -33.485 -90.81 -33.155 -90.48 ;
        RECT -33.485 -91.965 -33.155 -91.635 ;
        RECT -33.485 -93.325 -33.155 -92.995 ;
        RECT -33.485 -94.685 -33.155 -94.355 ;
        RECT -33.485 -96.045 -33.155 -95.715 ;
        RECT -33.485 -97.405 -33.155 -97.075 ;
        RECT -33.485 -100.125 -33.155 -99.795 ;
        RECT -33.485 -101.35 -33.155 -101.02 ;
        RECT -33.485 -102.845 -33.155 -102.515 ;
        RECT -33.485 -104.205 -33.155 -103.875 ;
        RECT -33.485 -105.565 -33.155 -105.235 ;
        RECT -33.485 -108.285 -33.155 -107.955 ;
        RECT -33.485 -109.645 -33.155 -109.315 ;
        RECT -33.485 -112.365 -33.155 -112.035 ;
        RECT -33.485 -113.725 -33.155 -113.395 ;
        RECT -33.485 -115.085 -33.155 -114.755 ;
        RECT -33.485 -116.445 -33.155 -116.115 ;
        RECT -33.485 -117.805 -33.155 -117.475 ;
        RECT -33.485 -119.165 -33.155 -118.835 ;
        RECT -33.485 -120.525 -33.155 -120.195 ;
        RECT -33.485 -121.885 -33.155 -121.555 ;
        RECT -33.485 -123.245 -33.155 -122.915 ;
        RECT -33.485 -125.965 -33.155 -125.635 ;
        RECT -33.485 -127.325 -33.155 -126.995 ;
        RECT -33.485 -128.685 -33.155 -128.355 ;
        RECT -33.485 -132.765 -33.155 -132.435 ;
        RECT -33.485 -134.125 -33.155 -133.795 ;
        RECT -33.485 -135.485 -33.155 -135.155 ;
        RECT -33.485 -136.845 -33.155 -136.515 ;
        RECT -33.485 -138.205 -33.155 -137.875 ;
        RECT -33.485 -140.925 -33.155 -140.595 ;
        RECT -33.485 -142.285 -33.155 -141.955 ;
        RECT -33.485 -143.645 -33.155 -143.315 ;
        RECT -33.485 -145.005 -33.155 -144.675 ;
        RECT -33.485 -146.365 -33.155 -146.035 ;
        RECT -33.485 -147.725 -33.155 -147.395 ;
        RECT -33.485 -150.445 -33.155 -150.115 ;
        RECT -33.485 -151.805 -33.155 -151.475 ;
        RECT -33.485 -155.885 -33.155 -155.555 ;
        RECT -33.485 -157.245 -33.155 -156.915 ;
        RECT -33.485 -158.605 -33.155 -158.275 ;
        RECT -33.485 -159.965 -33.155 -159.635 ;
        RECT -33.485 -161.325 -33.155 -160.995 ;
        RECT -33.485 -162.685 -33.155 -162.355 ;
        RECT -33.485 -164.045 -33.155 -163.715 ;
        RECT -33.485 -165.405 -33.155 -165.075 ;
        RECT -33.485 -166.765 -33.155 -166.435 ;
        RECT -33.485 -168.655 -33.155 -168.325 ;
        RECT -33.485 -169.485 -33.155 -169.155 ;
        RECT -33.485 -170.845 -33.155 -170.515 ;
        RECT -33.485 -172.205 -33.155 -171.875 ;
        RECT -33.485 -173.565 -33.155 -173.235 ;
        RECT -33.485 -174.925 -33.155 -174.595 ;
        RECT -33.485 -177.645 -33.155 -177.315 ;
        RECT -33.485 -183.29 -33.155 -182.16 ;
        RECT -33.48 -183.405 -33.16 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -32.125 205.875 -31.795 206.205 ;
        RECT -32.125 204.515 -31.795 204.845 ;
        RECT -32.125 203.155 -31.795 203.485 ;
        RECT -32.125 201.795 -31.795 202.125 ;
        RECT -32.125 200.435 -31.795 200.765 ;
        RECT -32.125 199.075 -31.795 199.405 ;
        RECT -32.125 197.715 -31.795 198.045 ;
        RECT -32.125 196.355 -31.795 196.685 ;
        RECT -32.125 194.995 -31.795 195.325 ;
        RECT -32.125 193.635 -31.795 193.965 ;
        RECT -32.125 192.275 -31.795 192.605 ;
        RECT -32.125 190.915 -31.795 191.245 ;
        RECT -32.125 189.555 -31.795 189.885 ;
        RECT -32.125 188.195 -31.795 188.525 ;
        RECT -32.125 186.835 -31.795 187.165 ;
        RECT -32.125 185.475 -31.795 185.805 ;
        RECT -32.125 184.115 -31.795 184.445 ;
        RECT -32.125 182.755 -31.795 183.085 ;
        RECT -32.125 181.395 -31.795 181.725 ;
        RECT -32.125 180.035 -31.795 180.365 ;
        RECT -32.125 178.675 -31.795 179.005 ;
        RECT -32.125 177.315 -31.795 177.645 ;
        RECT -32.125 175.955 -31.795 176.285 ;
        RECT -32.125 174.595 -31.795 174.925 ;
        RECT -32.125 173.235 -31.795 173.565 ;
        RECT -32.125 171.875 -31.795 172.205 ;
        RECT -32.125 170.515 -31.795 170.845 ;
        RECT -32.125 169.155 -31.795 169.485 ;
        RECT -32.125 167.795 -31.795 168.125 ;
        RECT -32.125 166.435 -31.795 166.765 ;
        RECT -32.125 165.075 -31.795 165.405 ;
        RECT -32.125 163.715 -31.795 164.045 ;
        RECT -32.125 162.355 -31.795 162.685 ;
        RECT -32.125 160.995 -31.795 161.325 ;
        RECT -32.125 159.635 -31.795 159.965 ;
        RECT -32.125 158.275 -31.795 158.605 ;
        RECT -32.125 156.915 -31.795 157.245 ;
        RECT -32.125 155.555 -31.795 155.885 ;
        RECT -32.125 154.195 -31.795 154.525 ;
        RECT -32.125 152.835 -31.795 153.165 ;
        RECT -32.125 151.475 -31.795 151.805 ;
        RECT -32.125 150.115 -31.795 150.445 ;
        RECT -32.125 148.755 -31.795 149.085 ;
        RECT -32.125 147.395 -31.795 147.725 ;
        RECT -32.125 146.035 -31.795 146.365 ;
        RECT -32.125 144.675 -31.795 145.005 ;
        RECT -32.125 143.315 -31.795 143.645 ;
        RECT -32.125 141.955 -31.795 142.285 ;
        RECT -32.125 140.595 -31.795 140.925 ;
        RECT -32.125 139.235 -31.795 139.565 ;
        RECT -32.125 137.875 -31.795 138.205 ;
        RECT -32.125 136.515 -31.795 136.845 ;
        RECT -32.125 135.155 -31.795 135.485 ;
        RECT -32.125 133.795 -31.795 134.125 ;
        RECT -32.125 132.435 -31.795 132.765 ;
        RECT -32.125 131.075 -31.795 131.405 ;
        RECT -32.125 129.715 -31.795 130.045 ;
        RECT -32.125 128.355 -31.795 128.685 ;
        RECT -32.125 126.995 -31.795 127.325 ;
        RECT -32.125 125.635 -31.795 125.965 ;
        RECT -32.125 124.275 -31.795 124.605 ;
        RECT -32.125 122.915 -31.795 123.245 ;
        RECT -32.125 121.555 -31.795 121.885 ;
        RECT -32.125 120.195 -31.795 120.525 ;
        RECT -32.125 118.835 -31.795 119.165 ;
        RECT -32.125 117.475 -31.795 117.805 ;
        RECT -32.125 116.115 -31.795 116.445 ;
        RECT -32.125 114.755 -31.795 115.085 ;
        RECT -32.125 113.395 -31.795 113.725 ;
        RECT -32.125 112.035 -31.795 112.365 ;
        RECT -32.125 110.675 -31.795 111.005 ;
        RECT -32.125 109.315 -31.795 109.645 ;
        RECT -32.125 107.955 -31.795 108.285 ;
        RECT -32.125 106.595 -31.795 106.925 ;
        RECT -32.125 105.235 -31.795 105.565 ;
        RECT -32.125 103.875 -31.795 104.205 ;
        RECT -32.125 102.515 -31.795 102.845 ;
        RECT -32.125 101.155 -31.795 101.485 ;
        RECT -32.125 99.795 -31.795 100.125 ;
        RECT -32.125 98.435 -31.795 98.765 ;
        RECT -32.125 97.075 -31.795 97.405 ;
        RECT -32.125 95.715 -31.795 96.045 ;
        RECT -32.125 94.355 -31.795 94.685 ;
        RECT -32.125 92.995 -31.795 93.325 ;
        RECT -32.125 91.635 -31.795 91.965 ;
        RECT -32.125 90.275 -31.795 90.605 ;
        RECT -32.125 88.915 -31.795 89.245 ;
        RECT -32.125 87.555 -31.795 87.885 ;
        RECT -32.125 86.195 -31.795 86.525 ;
        RECT -32.125 84.835 -31.795 85.165 ;
        RECT -32.125 83.475 -31.795 83.805 ;
        RECT -32.125 82.115 -31.795 82.445 ;
        RECT -32.125 80.755 -31.795 81.085 ;
        RECT -32.125 79.395 -31.795 79.725 ;
        RECT -32.125 78.035 -31.795 78.365 ;
        RECT -32.125 76.675 -31.795 77.005 ;
        RECT -32.125 75.315 -31.795 75.645 ;
        RECT -32.125 73.955 -31.795 74.285 ;
        RECT -32.125 72.595 -31.795 72.925 ;
        RECT -32.125 71.235 -31.795 71.565 ;
        RECT -32.125 69.875 -31.795 70.205 ;
        RECT -32.125 68.515 -31.795 68.845 ;
        RECT -32.125 67.155 -31.795 67.485 ;
        RECT -32.125 65.795 -31.795 66.125 ;
        RECT -32.125 64.435 -31.795 64.765 ;
        RECT -32.125 63.075 -31.795 63.405 ;
        RECT -32.125 61.715 -31.795 62.045 ;
        RECT -32.125 60.355 -31.795 60.685 ;
        RECT -32.125 58.995 -31.795 59.325 ;
        RECT -32.125 57.635 -31.795 57.965 ;
        RECT -32.125 56.275 -31.795 56.605 ;
        RECT -32.125 54.915 -31.795 55.245 ;
        RECT -32.125 53.555 -31.795 53.885 ;
        RECT -32.125 52.195 -31.795 52.525 ;
        RECT -32.125 50.835 -31.795 51.165 ;
        RECT -32.125 49.475 -31.795 49.805 ;
        RECT -32.125 48.115 -31.795 48.445 ;
        RECT -32.125 46.755 -31.795 47.085 ;
        RECT -32.125 45.395 -31.795 45.725 ;
        RECT -32.125 44.035 -31.795 44.365 ;
        RECT -32.125 42.675 -31.795 43.005 ;
        RECT -32.125 41.315 -31.795 41.645 ;
        RECT -32.125 39.955 -31.795 40.285 ;
        RECT -32.125 38.595 -31.795 38.925 ;
        RECT -32.125 37.235 -31.795 37.565 ;
        RECT -32.125 35.875 -31.795 36.205 ;
        RECT -32.125 34.515 -31.795 34.845 ;
        RECT -32.125 33.155 -31.795 33.485 ;
        RECT -32.125 31.795 -31.795 32.125 ;
        RECT -32.125 30.435 -31.795 30.765 ;
        RECT -32.125 29.075 -31.795 29.405 ;
        RECT -32.125 27.715 -31.795 28.045 ;
        RECT -32.125 26.355 -31.795 26.685 ;
        RECT -32.125 24.995 -31.795 25.325 ;
        RECT -32.125 23.635 -31.795 23.965 ;
        RECT -32.125 22.275 -31.795 22.605 ;
        RECT -32.125 20.915 -31.795 21.245 ;
        RECT -32.125 19.555 -31.795 19.885 ;
        RECT -32.125 18.195 -31.795 18.525 ;
        RECT -32.125 16.835 -31.795 17.165 ;
        RECT -32.125 15.475 -31.795 15.805 ;
        RECT -32.125 14.115 -31.795 14.445 ;
        RECT -32.125 12.755 -31.795 13.085 ;
        RECT -32.125 11.395 -31.795 11.725 ;
        RECT -32.125 10.035 -31.795 10.365 ;
        RECT -32.125 8.675 -31.795 9.005 ;
        RECT -32.125 7.315 -31.795 7.645 ;
        RECT -32.125 5.955 -31.795 6.285 ;
        RECT -32.125 4.595 -31.795 4.925 ;
        RECT -32.125 3.235 -31.795 3.565 ;
        RECT -32.125 1.875 -31.795 2.205 ;
        RECT -32.125 0.515 -31.795 0.845 ;
        RECT -32.125 -0.845 -31.795 -0.515 ;
        RECT -32.125 -7.645 -31.795 -7.315 ;
        RECT -32.125 -9.005 -31.795 -8.675 ;
        RECT -32.125 -10.365 -31.795 -10.035 ;
        RECT -32.125 -14.445 -31.795 -14.115 ;
        RECT -32.125 -15.805 -31.795 -15.475 ;
        RECT -32.125 -17.165 -31.795 -16.835 ;
        RECT -32.125 -18.525 -31.795 -18.195 ;
        RECT -32.125 -19.885 -31.795 -19.555 ;
        RECT -32.125 -21.245 -31.795 -20.915 ;
        RECT -32.125 -22.605 -31.795 -22.275 ;
        RECT -32.125 -23.965 -31.795 -23.635 ;
        RECT -32.125 -25.325 -31.795 -24.995 ;
        RECT -32.125 -32.125 -31.795 -31.795 ;
        RECT -32.125 -33.71 -31.795 -33.38 ;
        RECT -32.125 -34.845 -31.795 -34.515 ;
        RECT -32.125 -36.205 -31.795 -35.875 ;
        RECT -32.125 -38.925 -31.795 -38.595 ;
        RECT -32.125 -39.75 -31.795 -39.42 ;
        RECT -32.125 -41.645 -31.795 -41.315 ;
        RECT -32.125 -44.365 -31.795 -44.035 ;
        RECT -32.125 -49.805 -31.795 -49.475 ;
        RECT -32.125 -51.165 -31.795 -50.835 ;
        RECT -32.125 -53.885 -31.795 -53.555 ;
        RECT -32.125 -55.245 -31.795 -54.915 ;
        RECT -32.125 -59.325 -31.795 -58.995 ;
        RECT -32.125 -60.685 -31.795 -60.355 ;
        RECT -32.125 -68.845 -31.795 -68.515 ;
        RECT -32.125 -70.205 -31.795 -69.875 ;
        RECT -32.125 -71.565 -31.795 -71.235 ;
        RECT -32.125 -72.925 -31.795 -72.595 ;
        RECT -32.125 -74.285 -31.795 -73.955 ;
        RECT -32.125 -75.645 -31.795 -75.315 ;
        RECT -32.125 -77.005 -31.795 -76.675 ;
        RECT -32.125 -78.365 -31.795 -78.035 ;
        RECT -32.125 -79.725 -31.795 -79.395 ;
        RECT -32.125 -81.085 -31.795 -80.755 ;
        RECT -32.125 -82.445 -31.795 -82.115 ;
        RECT -32.125 -83.805 -31.795 -83.475 ;
        RECT -32.125 -85.165 -31.795 -84.835 ;
        RECT -32.125 -86.525 -31.795 -86.195 ;
        RECT -32.125 -87.885 -31.795 -87.555 ;
        RECT -32.125 -89.245 -31.795 -88.915 ;
        RECT -32.125 -90.81 -31.795 -90.48 ;
        RECT -32.125 -91.965 -31.795 -91.635 ;
        RECT -32.125 -93.325 -31.795 -92.995 ;
        RECT -32.125 -94.685 -31.795 -94.355 ;
        RECT -32.125 -96.045 -31.795 -95.715 ;
        RECT -32.125 -97.405 -31.795 -97.075 ;
        RECT -32.125 -100.125 -31.795 -99.795 ;
        RECT -32.125 -101.35 -31.795 -101.02 ;
        RECT -32.125 -102.845 -31.795 -102.515 ;
        RECT -32.125 -104.205 -31.795 -103.875 ;
        RECT -32.125 -105.565 -31.795 -105.235 ;
        RECT -32.125 -108.285 -31.795 -107.955 ;
        RECT -32.125 -109.645 -31.795 -109.315 ;
        RECT -32.125 -112.365 -31.795 -112.035 ;
        RECT -32.125 -113.725 -31.795 -113.395 ;
        RECT -32.125 -115.085 -31.795 -114.755 ;
        RECT -32.125 -116.445 -31.795 -116.115 ;
        RECT -32.125 -117.805 -31.795 -117.475 ;
        RECT -32.125 -119.165 -31.795 -118.835 ;
        RECT -32.125 -120.525 -31.795 -120.195 ;
        RECT -32.125 -121.885 -31.795 -121.555 ;
        RECT -32.125 -123.245 -31.795 -122.915 ;
        RECT -32.125 -125.965 -31.795 -125.635 ;
        RECT -32.125 -127.325 -31.795 -126.995 ;
        RECT -32.125 -128.685 -31.795 -128.355 ;
        RECT -32.125 -132.765 -31.795 -132.435 ;
        RECT -32.125 -134.125 -31.795 -133.795 ;
        RECT -32.125 -135.485 -31.795 -135.155 ;
        RECT -32.125 -136.845 -31.795 -136.515 ;
        RECT -32.125 -140.925 -31.795 -140.595 ;
        RECT -32.125 -142.285 -31.795 -141.955 ;
        RECT -32.125 -143.645 -31.795 -143.315 ;
        RECT -32.125 -145.005 -31.795 -144.675 ;
        RECT -32.125 -146.365 -31.795 -146.035 ;
        RECT -32.125 -147.725 -31.795 -147.395 ;
        RECT -32.125 -150.445 -31.795 -150.115 ;
        RECT -32.125 -151.805 -31.795 -151.475 ;
        RECT -32.125 -155.885 -31.795 -155.555 ;
        RECT -32.125 -157.245 -31.795 -156.915 ;
        RECT -32.125 -158.605 -31.795 -158.275 ;
        RECT -32.125 -159.965 -31.795 -159.635 ;
        RECT -32.125 -161.325 -31.795 -160.995 ;
        RECT -32.125 -162.685 -31.795 -162.355 ;
        RECT -32.125 -164.045 -31.795 -163.715 ;
        RECT -32.125 -165.405 -31.795 -165.075 ;
        RECT -32.125 -166.765 -31.795 -166.435 ;
        RECT -32.125 -168.655 -31.795 -168.325 ;
        RECT -32.125 -169.485 -31.795 -169.155 ;
        RECT -32.125 -170.845 -31.795 -170.515 ;
        RECT -32.125 -172.205 -31.795 -171.875 ;
        RECT -32.125 -173.565 -31.795 -173.235 ;
        RECT -32.125 -174.925 -31.795 -174.595 ;
        RECT -32.125 -177.645 -31.795 -177.315 ;
        RECT -32.125 -183.29 -31.795 -182.16 ;
        RECT -32.12 -183.405 -31.8 245.285 ;
        RECT -32.125 244.04 -31.795 245.17 ;
        RECT -32.125 239.875 -31.795 240.205 ;
        RECT -32.125 238.515 -31.795 238.845 ;
        RECT -32.125 237.155 -31.795 237.485 ;
        RECT -32.125 235.795 -31.795 236.125 ;
        RECT -32.125 234.435 -31.795 234.765 ;
        RECT -32.125 233.075 -31.795 233.405 ;
        RECT -32.125 231.715 -31.795 232.045 ;
        RECT -32.125 230.355 -31.795 230.685 ;
        RECT -32.125 228.995 -31.795 229.325 ;
        RECT -32.125 227.635 -31.795 227.965 ;
        RECT -32.125 226.275 -31.795 226.605 ;
        RECT -32.125 224.915 -31.795 225.245 ;
        RECT -32.125 223.555 -31.795 223.885 ;
        RECT -32.125 222.195 -31.795 222.525 ;
        RECT -32.125 220.835 -31.795 221.165 ;
        RECT -32.125 219.475 -31.795 219.805 ;
        RECT -32.125 218.115 -31.795 218.445 ;
        RECT -32.125 216.755 -31.795 217.085 ;
        RECT -32.125 215.395 -31.795 215.725 ;
        RECT -32.125 214.035 -31.795 214.365 ;
        RECT -32.125 212.675 -31.795 213.005 ;
        RECT -32.125 211.315 -31.795 211.645 ;
        RECT -32.125 209.955 -31.795 210.285 ;
        RECT -32.125 208.595 -31.795 208.925 ;
        RECT -32.125 207.235 -31.795 207.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -41.645 -174.925 -41.315 -174.595 ;
        RECT -41.645 -177.645 -41.315 -177.315 ;
        RECT -41.645 -183.29 -41.315 -182.16 ;
        RECT -41.64 -183.405 -41.32 -172.56 ;
    END
    PORT
      LAYER met3 ;
        RECT -40.285 244.04 -39.955 245.17 ;
        RECT -40.285 239.875 -39.955 240.205 ;
        RECT -40.285 238.515 -39.955 238.845 ;
        RECT -40.285 237.155 -39.955 237.485 ;
        RECT -40.285 235.795 -39.955 236.125 ;
        RECT -40.285 234.435 -39.955 234.765 ;
        RECT -40.285 233.075 -39.955 233.405 ;
        RECT -40.285 231.715 -39.955 232.045 ;
        RECT -40.285 230.355 -39.955 230.685 ;
        RECT -40.285 228.995 -39.955 229.325 ;
        RECT -40.285 227.635 -39.955 227.965 ;
        RECT -40.285 226.275 -39.955 226.605 ;
        RECT -40.285 224.915 -39.955 225.245 ;
        RECT -40.285 223.555 -39.955 223.885 ;
        RECT -40.285 222.195 -39.955 222.525 ;
        RECT -40.285 220.835 -39.955 221.165 ;
        RECT -40.285 219.475 -39.955 219.805 ;
        RECT -40.285 218.115 -39.955 218.445 ;
        RECT -40.285 216.755 -39.955 217.085 ;
        RECT -40.285 215.395 -39.955 215.725 ;
        RECT -40.285 214.035 -39.955 214.365 ;
        RECT -40.285 212.675 -39.955 213.005 ;
        RECT -40.285 211.315 -39.955 211.645 ;
        RECT -40.285 209.955 -39.955 210.285 ;
        RECT -40.285 208.595 -39.955 208.925 ;
        RECT -40.285 207.235 -39.955 207.565 ;
        RECT -40.285 205.875 -39.955 206.205 ;
        RECT -40.285 204.515 -39.955 204.845 ;
        RECT -40.285 203.155 -39.955 203.485 ;
        RECT -40.285 201.795 -39.955 202.125 ;
        RECT -40.285 200.435 -39.955 200.765 ;
        RECT -40.285 199.075 -39.955 199.405 ;
        RECT -40.285 197.715 -39.955 198.045 ;
        RECT -40.285 196.355 -39.955 196.685 ;
        RECT -40.285 194.995 -39.955 195.325 ;
        RECT -40.285 193.635 -39.955 193.965 ;
        RECT -40.285 192.275 -39.955 192.605 ;
        RECT -40.285 190.915 -39.955 191.245 ;
        RECT -40.285 189.555 -39.955 189.885 ;
        RECT -40.285 188.195 -39.955 188.525 ;
        RECT -40.285 186.835 -39.955 187.165 ;
        RECT -40.285 185.475 -39.955 185.805 ;
        RECT -40.285 184.115 -39.955 184.445 ;
        RECT -40.285 182.755 -39.955 183.085 ;
        RECT -40.285 181.395 -39.955 181.725 ;
        RECT -40.285 180.035 -39.955 180.365 ;
        RECT -40.285 178.675 -39.955 179.005 ;
        RECT -40.285 177.315 -39.955 177.645 ;
        RECT -40.285 175.955 -39.955 176.285 ;
        RECT -40.285 174.595 -39.955 174.925 ;
        RECT -40.285 173.235 -39.955 173.565 ;
        RECT -40.285 171.875 -39.955 172.205 ;
        RECT -40.285 170.515 -39.955 170.845 ;
        RECT -40.285 169.155 -39.955 169.485 ;
        RECT -40.285 167.795 -39.955 168.125 ;
        RECT -40.285 166.435 -39.955 166.765 ;
        RECT -40.285 165.075 -39.955 165.405 ;
        RECT -40.285 163.715 -39.955 164.045 ;
        RECT -40.285 162.355 -39.955 162.685 ;
        RECT -40.285 160.995 -39.955 161.325 ;
        RECT -40.285 159.635 -39.955 159.965 ;
        RECT -40.285 158.275 -39.955 158.605 ;
        RECT -40.285 156.915 -39.955 157.245 ;
        RECT -40.285 155.555 -39.955 155.885 ;
        RECT -40.285 154.195 -39.955 154.525 ;
        RECT -40.285 152.835 -39.955 153.165 ;
        RECT -40.285 151.475 -39.955 151.805 ;
        RECT -40.285 150.115 -39.955 150.445 ;
        RECT -40.285 148.755 -39.955 149.085 ;
        RECT -40.285 147.395 -39.955 147.725 ;
        RECT -40.285 146.035 -39.955 146.365 ;
        RECT -40.285 144.675 -39.955 145.005 ;
        RECT -40.285 143.315 -39.955 143.645 ;
        RECT -40.285 141.955 -39.955 142.285 ;
        RECT -40.285 140.595 -39.955 140.925 ;
        RECT -40.285 139.235 -39.955 139.565 ;
        RECT -40.285 137.875 -39.955 138.205 ;
        RECT -40.285 136.515 -39.955 136.845 ;
        RECT -40.285 135.155 -39.955 135.485 ;
        RECT -40.285 133.795 -39.955 134.125 ;
        RECT -40.285 132.435 -39.955 132.765 ;
        RECT -40.285 131.075 -39.955 131.405 ;
        RECT -40.285 129.715 -39.955 130.045 ;
        RECT -40.285 128.355 -39.955 128.685 ;
        RECT -40.285 126.995 -39.955 127.325 ;
        RECT -40.285 125.635 -39.955 125.965 ;
        RECT -40.285 124.275 -39.955 124.605 ;
        RECT -40.285 122.915 -39.955 123.245 ;
        RECT -40.285 121.555 -39.955 121.885 ;
        RECT -40.285 120.195 -39.955 120.525 ;
        RECT -40.285 118.835 -39.955 119.165 ;
        RECT -40.285 117.475 -39.955 117.805 ;
        RECT -40.285 116.115 -39.955 116.445 ;
        RECT -40.285 114.755 -39.955 115.085 ;
        RECT -40.285 113.395 -39.955 113.725 ;
        RECT -40.285 112.035 -39.955 112.365 ;
        RECT -40.285 110.675 -39.955 111.005 ;
        RECT -40.285 109.315 -39.955 109.645 ;
        RECT -40.285 107.955 -39.955 108.285 ;
        RECT -40.285 106.595 -39.955 106.925 ;
        RECT -40.285 105.235 -39.955 105.565 ;
        RECT -40.285 103.875 -39.955 104.205 ;
        RECT -40.285 102.515 -39.955 102.845 ;
        RECT -40.285 101.155 -39.955 101.485 ;
        RECT -40.285 99.795 -39.955 100.125 ;
        RECT -40.285 98.435 -39.955 98.765 ;
        RECT -40.285 97.075 -39.955 97.405 ;
        RECT -40.285 95.715 -39.955 96.045 ;
        RECT -40.285 94.355 -39.955 94.685 ;
        RECT -40.285 92.995 -39.955 93.325 ;
        RECT -40.285 91.635 -39.955 91.965 ;
        RECT -40.285 90.275 -39.955 90.605 ;
        RECT -40.285 88.915 -39.955 89.245 ;
        RECT -40.285 87.555 -39.955 87.885 ;
        RECT -40.285 86.195 -39.955 86.525 ;
        RECT -40.285 84.835 -39.955 85.165 ;
        RECT -40.285 83.475 -39.955 83.805 ;
        RECT -40.285 82.115 -39.955 82.445 ;
        RECT -40.285 80.755 -39.955 81.085 ;
        RECT -40.285 79.395 -39.955 79.725 ;
        RECT -40.285 78.035 -39.955 78.365 ;
        RECT -40.285 76.675 -39.955 77.005 ;
        RECT -40.285 75.315 -39.955 75.645 ;
        RECT -40.285 73.955 -39.955 74.285 ;
        RECT -40.285 72.595 -39.955 72.925 ;
        RECT -40.285 71.235 -39.955 71.565 ;
        RECT -40.285 69.875 -39.955 70.205 ;
        RECT -40.285 68.515 -39.955 68.845 ;
        RECT -40.285 67.155 -39.955 67.485 ;
        RECT -40.285 65.795 -39.955 66.125 ;
        RECT -40.285 64.435 -39.955 64.765 ;
        RECT -40.285 63.075 -39.955 63.405 ;
        RECT -40.285 61.715 -39.955 62.045 ;
        RECT -40.285 60.355 -39.955 60.685 ;
        RECT -40.285 58.995 -39.955 59.325 ;
        RECT -40.285 57.635 -39.955 57.965 ;
        RECT -40.285 56.275 -39.955 56.605 ;
        RECT -40.285 54.915 -39.955 55.245 ;
        RECT -40.285 53.555 -39.955 53.885 ;
        RECT -40.285 52.195 -39.955 52.525 ;
        RECT -40.285 50.835 -39.955 51.165 ;
        RECT -40.285 49.475 -39.955 49.805 ;
        RECT -40.285 48.115 -39.955 48.445 ;
        RECT -40.285 46.755 -39.955 47.085 ;
        RECT -40.285 45.395 -39.955 45.725 ;
        RECT -40.285 44.035 -39.955 44.365 ;
        RECT -40.285 42.675 -39.955 43.005 ;
        RECT -40.285 41.315 -39.955 41.645 ;
        RECT -40.285 39.955 -39.955 40.285 ;
        RECT -40.285 38.595 -39.955 38.925 ;
        RECT -40.285 37.235 -39.955 37.565 ;
        RECT -40.285 35.875 -39.955 36.205 ;
        RECT -40.285 34.515 -39.955 34.845 ;
        RECT -40.285 33.155 -39.955 33.485 ;
        RECT -40.285 31.795 -39.955 32.125 ;
        RECT -40.285 30.435 -39.955 30.765 ;
        RECT -40.285 29.075 -39.955 29.405 ;
        RECT -40.285 27.715 -39.955 28.045 ;
        RECT -40.285 26.355 -39.955 26.685 ;
        RECT -40.285 24.995 -39.955 25.325 ;
        RECT -40.285 23.635 -39.955 23.965 ;
        RECT -40.285 22.275 -39.955 22.605 ;
        RECT -40.285 20.915 -39.955 21.245 ;
        RECT -40.285 19.555 -39.955 19.885 ;
        RECT -40.285 18.195 -39.955 18.525 ;
        RECT -40.285 16.835 -39.955 17.165 ;
        RECT -40.285 15.475 -39.955 15.805 ;
        RECT -40.285 14.115 -39.955 14.445 ;
        RECT -40.285 12.755 -39.955 13.085 ;
        RECT -40.285 11.395 -39.955 11.725 ;
        RECT -40.285 10.035 -39.955 10.365 ;
        RECT -40.285 8.675 -39.955 9.005 ;
        RECT -40.285 7.315 -39.955 7.645 ;
        RECT -40.285 5.955 -39.955 6.285 ;
        RECT -40.285 4.595 -39.955 4.925 ;
        RECT -40.285 3.235 -39.955 3.565 ;
        RECT -40.285 1.875 -39.955 2.205 ;
        RECT -40.285 0.515 -39.955 0.845 ;
        RECT -40.285 -0.845 -39.955 -0.515 ;
        RECT -40.285 -2.205 -39.955 -1.875 ;
        RECT -40.285 -3.565 -39.955 -3.235 ;
        RECT -40.285 -4.925 -39.955 -4.595 ;
        RECT -40.285 -6.285 -39.955 -5.955 ;
        RECT -40.285 -10.365 -39.955 -10.035 ;
        RECT -40.285 -14.445 -39.955 -14.115 ;
        RECT -40.285 -15.805 -39.955 -15.475 ;
        RECT -40.285 -17.165 -39.955 -16.835 ;
        RECT -40.285 -18.525 -39.955 -18.195 ;
        RECT -40.285 -19.885 -39.955 -19.555 ;
        RECT -40.285 -21.245 -39.955 -20.915 ;
        RECT -40.285 -22.605 -39.955 -22.275 ;
        RECT -40.285 -23.965 -39.955 -23.635 ;
        RECT -40.285 -25.325 -39.955 -24.995 ;
        RECT -40.285 -32.125 -39.955 -31.795 ;
        RECT -40.285 -33.71 -39.955 -33.38 ;
        RECT -40.285 -34.845 -39.955 -34.515 ;
        RECT -40.285 -36.205 -39.955 -35.875 ;
        RECT -40.285 -38.925 -39.955 -38.595 ;
        RECT -40.285 -39.75 -39.955 -39.42 ;
        RECT -40.285 -41.645 -39.955 -41.315 ;
        RECT -40.285 -44.365 -39.955 -44.035 ;
        RECT -40.285 -49.805 -39.955 -49.475 ;
        RECT -40.285 -51.165 -39.955 -50.835 ;
        RECT -40.285 -53.885 -39.955 -53.555 ;
        RECT -40.285 -55.245 -39.955 -54.915 ;
        RECT -40.285 -59.325 -39.955 -58.995 ;
        RECT -40.285 -60.685 -39.955 -60.355 ;
        RECT -40.285 -67.485 -39.955 -67.155 ;
        RECT -40.285 -70.205 -39.955 -69.875 ;
        RECT -40.285 -71.565 -39.955 -71.235 ;
        RECT -40.285 -72.925 -39.955 -72.595 ;
        RECT -40.285 -74.285 -39.955 -73.955 ;
        RECT -40.285 -75.645 -39.955 -75.315 ;
        RECT -40.285 -77.005 -39.955 -76.675 ;
        RECT -40.285 -78.365 -39.955 -78.035 ;
        RECT -40.285 -79.725 -39.955 -79.395 ;
        RECT -40.285 -81.085 -39.955 -80.755 ;
        RECT -40.285 -82.445 -39.955 -82.115 ;
        RECT -40.285 -83.805 -39.955 -83.475 ;
        RECT -40.285 -85.165 -39.955 -84.835 ;
        RECT -40.285 -86.525 -39.955 -86.195 ;
        RECT -40.285 -87.885 -39.955 -87.555 ;
        RECT -40.285 -89.245 -39.955 -88.915 ;
        RECT -40.285 -90.81 -39.955 -90.48 ;
        RECT -40.285 -91.965 -39.955 -91.635 ;
        RECT -40.285 -93.325 -39.955 -92.995 ;
        RECT -40.285 -94.685 -39.955 -94.355 ;
        RECT -40.285 -96.045 -39.955 -95.715 ;
        RECT -40.285 -97.405 -39.955 -97.075 ;
        RECT -40.285 -100.125 -39.955 -99.795 ;
        RECT -40.285 -101.35 -39.955 -101.02 ;
        RECT -40.285 -102.845 -39.955 -102.515 ;
        RECT -40.285 -104.205 -39.955 -103.875 ;
        RECT -40.285 -105.565 -39.955 -105.235 ;
        RECT -40.285 -108.285 -39.955 -107.955 ;
        RECT -40.285 -109.645 -39.955 -109.315 ;
        RECT -40.285 -113.725 -39.955 -113.395 ;
        RECT -40.285 -115.085 -39.955 -114.755 ;
        RECT -40.285 -116.445 -39.955 -116.115 ;
        RECT -40.285 -117.805 -39.955 -117.475 ;
        RECT -40.285 -119.165 -39.955 -118.835 ;
        RECT -40.285 -120.525 -39.955 -120.195 ;
        RECT -40.285 -121.885 -39.955 -121.555 ;
        RECT -40.285 -123.245 -39.955 -122.915 ;
        RECT -40.285 -124.605 -39.955 -124.275 ;
        RECT -40.285 -125.965 -39.955 -125.635 ;
        RECT -40.285 -127.325 -39.955 -126.995 ;
        RECT -40.285 -128.685 -39.955 -128.355 ;
        RECT -40.285 -130.045 -39.955 -129.715 ;
        RECT -40.285 -132.765 -39.955 -132.435 ;
        RECT -40.285 -134.125 -39.955 -133.795 ;
        RECT -40.285 -135.485 -39.955 -135.155 ;
        RECT -40.285 -136.845 -39.955 -136.515 ;
        RECT -40.285 -138.205 -39.955 -137.875 ;
        RECT -40.285 -139.565 -39.955 -139.235 ;
        RECT -40.285 -140.925 -39.955 -140.595 ;
        RECT -40.285 -142.285 -39.955 -141.955 ;
        RECT -40.285 -143.645 -39.955 -143.315 ;
        RECT -40.285 -145.005 -39.955 -144.675 ;
        RECT -40.285 -146.365 -39.955 -146.035 ;
        RECT -40.285 -147.725 -39.955 -147.395 ;
        RECT -40.285 -150.445 -39.955 -150.115 ;
        RECT -40.285 -151.805 -39.955 -151.475 ;
        RECT -40.285 -154.525 -39.955 -154.195 ;
        RECT -40.285 -157.245 -39.955 -156.915 ;
        RECT -40.285 -158.605 -39.955 -158.275 ;
        RECT -40.285 -159.965 -39.955 -159.635 ;
        RECT -40.285 -161.325 -39.955 -160.995 ;
        RECT -40.285 -162.685 -39.955 -162.355 ;
        RECT -40.285 -164.045 -39.955 -163.715 ;
        RECT -40.285 -165.405 -39.955 -165.075 ;
        RECT -40.285 -166.765 -39.955 -166.435 ;
        RECT -40.285 -168.655 -39.955 -168.325 ;
        RECT -40.285 -169.485 -39.955 -169.155 ;
        RECT -40.285 -170.845 -39.955 -170.515 ;
        RECT -40.28 -172.2 -39.96 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -38.925 244.04 -38.595 245.17 ;
        RECT -38.925 239.875 -38.595 240.205 ;
        RECT -38.925 238.515 -38.595 238.845 ;
        RECT -38.925 237.155 -38.595 237.485 ;
        RECT -38.925 235.795 -38.595 236.125 ;
        RECT -38.925 234.435 -38.595 234.765 ;
        RECT -38.925 233.075 -38.595 233.405 ;
        RECT -38.925 231.715 -38.595 232.045 ;
        RECT -38.925 230.355 -38.595 230.685 ;
        RECT -38.925 228.995 -38.595 229.325 ;
        RECT -38.925 227.635 -38.595 227.965 ;
        RECT -38.925 226.275 -38.595 226.605 ;
        RECT -38.925 224.915 -38.595 225.245 ;
        RECT -38.925 223.555 -38.595 223.885 ;
        RECT -38.925 222.195 -38.595 222.525 ;
        RECT -38.925 220.835 -38.595 221.165 ;
        RECT -38.925 219.475 -38.595 219.805 ;
        RECT -38.925 218.115 -38.595 218.445 ;
        RECT -38.925 216.755 -38.595 217.085 ;
        RECT -38.925 215.395 -38.595 215.725 ;
        RECT -38.925 214.035 -38.595 214.365 ;
        RECT -38.925 212.675 -38.595 213.005 ;
        RECT -38.925 211.315 -38.595 211.645 ;
        RECT -38.925 209.955 -38.595 210.285 ;
        RECT -38.925 208.595 -38.595 208.925 ;
        RECT -38.925 207.235 -38.595 207.565 ;
        RECT -38.925 205.875 -38.595 206.205 ;
        RECT -38.925 204.515 -38.595 204.845 ;
        RECT -38.925 203.155 -38.595 203.485 ;
        RECT -38.925 201.795 -38.595 202.125 ;
        RECT -38.925 200.435 -38.595 200.765 ;
        RECT -38.925 199.075 -38.595 199.405 ;
        RECT -38.925 197.715 -38.595 198.045 ;
        RECT -38.925 196.355 -38.595 196.685 ;
        RECT -38.925 194.995 -38.595 195.325 ;
        RECT -38.925 193.635 -38.595 193.965 ;
        RECT -38.925 192.275 -38.595 192.605 ;
        RECT -38.925 190.915 -38.595 191.245 ;
        RECT -38.925 189.555 -38.595 189.885 ;
        RECT -38.925 188.195 -38.595 188.525 ;
        RECT -38.925 186.835 -38.595 187.165 ;
        RECT -38.925 185.475 -38.595 185.805 ;
        RECT -38.925 184.115 -38.595 184.445 ;
        RECT -38.925 182.755 -38.595 183.085 ;
        RECT -38.925 181.395 -38.595 181.725 ;
        RECT -38.925 180.035 -38.595 180.365 ;
        RECT -38.925 178.675 -38.595 179.005 ;
        RECT -38.925 177.315 -38.595 177.645 ;
        RECT -38.925 175.955 -38.595 176.285 ;
        RECT -38.925 174.595 -38.595 174.925 ;
        RECT -38.925 173.235 -38.595 173.565 ;
        RECT -38.925 171.875 -38.595 172.205 ;
        RECT -38.925 170.515 -38.595 170.845 ;
        RECT -38.925 169.155 -38.595 169.485 ;
        RECT -38.925 167.795 -38.595 168.125 ;
        RECT -38.925 166.435 -38.595 166.765 ;
        RECT -38.925 165.075 -38.595 165.405 ;
        RECT -38.925 163.715 -38.595 164.045 ;
        RECT -38.925 162.355 -38.595 162.685 ;
        RECT -38.925 160.995 -38.595 161.325 ;
        RECT -38.925 159.635 -38.595 159.965 ;
        RECT -38.925 158.275 -38.595 158.605 ;
        RECT -38.925 156.915 -38.595 157.245 ;
        RECT -38.925 155.555 -38.595 155.885 ;
        RECT -38.925 154.195 -38.595 154.525 ;
        RECT -38.925 152.835 -38.595 153.165 ;
        RECT -38.925 151.475 -38.595 151.805 ;
        RECT -38.925 150.115 -38.595 150.445 ;
        RECT -38.925 148.755 -38.595 149.085 ;
        RECT -38.925 147.395 -38.595 147.725 ;
        RECT -38.925 146.035 -38.595 146.365 ;
        RECT -38.925 144.675 -38.595 145.005 ;
        RECT -38.925 143.315 -38.595 143.645 ;
        RECT -38.925 141.955 -38.595 142.285 ;
        RECT -38.925 140.595 -38.595 140.925 ;
        RECT -38.925 139.235 -38.595 139.565 ;
        RECT -38.925 137.875 -38.595 138.205 ;
        RECT -38.925 136.515 -38.595 136.845 ;
        RECT -38.925 135.155 -38.595 135.485 ;
        RECT -38.925 133.795 -38.595 134.125 ;
        RECT -38.925 132.435 -38.595 132.765 ;
        RECT -38.925 131.075 -38.595 131.405 ;
        RECT -38.925 129.715 -38.595 130.045 ;
        RECT -38.925 128.355 -38.595 128.685 ;
        RECT -38.925 126.995 -38.595 127.325 ;
        RECT -38.925 125.635 -38.595 125.965 ;
        RECT -38.925 124.275 -38.595 124.605 ;
        RECT -38.925 122.915 -38.595 123.245 ;
        RECT -38.925 121.555 -38.595 121.885 ;
        RECT -38.925 120.195 -38.595 120.525 ;
        RECT -38.925 118.835 -38.595 119.165 ;
        RECT -38.925 117.475 -38.595 117.805 ;
        RECT -38.925 116.115 -38.595 116.445 ;
        RECT -38.925 114.755 -38.595 115.085 ;
        RECT -38.925 113.395 -38.595 113.725 ;
        RECT -38.925 112.035 -38.595 112.365 ;
        RECT -38.925 110.675 -38.595 111.005 ;
        RECT -38.925 109.315 -38.595 109.645 ;
        RECT -38.925 107.955 -38.595 108.285 ;
        RECT -38.925 106.595 -38.595 106.925 ;
        RECT -38.925 105.235 -38.595 105.565 ;
        RECT -38.925 103.875 -38.595 104.205 ;
        RECT -38.925 102.515 -38.595 102.845 ;
        RECT -38.925 101.155 -38.595 101.485 ;
        RECT -38.925 99.795 -38.595 100.125 ;
        RECT -38.925 98.435 -38.595 98.765 ;
        RECT -38.925 97.075 -38.595 97.405 ;
        RECT -38.925 95.715 -38.595 96.045 ;
        RECT -38.925 94.355 -38.595 94.685 ;
        RECT -38.925 92.995 -38.595 93.325 ;
        RECT -38.925 91.635 -38.595 91.965 ;
        RECT -38.925 90.275 -38.595 90.605 ;
        RECT -38.925 88.915 -38.595 89.245 ;
        RECT -38.925 87.555 -38.595 87.885 ;
        RECT -38.925 86.195 -38.595 86.525 ;
        RECT -38.925 84.835 -38.595 85.165 ;
        RECT -38.925 83.475 -38.595 83.805 ;
        RECT -38.925 82.115 -38.595 82.445 ;
        RECT -38.925 80.755 -38.595 81.085 ;
        RECT -38.925 79.395 -38.595 79.725 ;
        RECT -38.925 78.035 -38.595 78.365 ;
        RECT -38.925 76.675 -38.595 77.005 ;
        RECT -38.925 75.315 -38.595 75.645 ;
        RECT -38.925 73.955 -38.595 74.285 ;
        RECT -38.925 72.595 -38.595 72.925 ;
        RECT -38.925 71.235 -38.595 71.565 ;
        RECT -38.925 69.875 -38.595 70.205 ;
        RECT -38.925 68.515 -38.595 68.845 ;
        RECT -38.925 67.155 -38.595 67.485 ;
        RECT -38.925 65.795 -38.595 66.125 ;
        RECT -38.925 64.435 -38.595 64.765 ;
        RECT -38.925 63.075 -38.595 63.405 ;
        RECT -38.925 61.715 -38.595 62.045 ;
        RECT -38.925 60.355 -38.595 60.685 ;
        RECT -38.925 58.995 -38.595 59.325 ;
        RECT -38.925 57.635 -38.595 57.965 ;
        RECT -38.925 56.275 -38.595 56.605 ;
        RECT -38.925 54.915 -38.595 55.245 ;
        RECT -38.925 53.555 -38.595 53.885 ;
        RECT -38.925 52.195 -38.595 52.525 ;
        RECT -38.925 50.835 -38.595 51.165 ;
        RECT -38.925 49.475 -38.595 49.805 ;
        RECT -38.925 48.115 -38.595 48.445 ;
        RECT -38.925 46.755 -38.595 47.085 ;
        RECT -38.925 45.395 -38.595 45.725 ;
        RECT -38.925 44.035 -38.595 44.365 ;
        RECT -38.925 42.675 -38.595 43.005 ;
        RECT -38.925 41.315 -38.595 41.645 ;
        RECT -38.925 39.955 -38.595 40.285 ;
        RECT -38.925 38.595 -38.595 38.925 ;
        RECT -38.925 37.235 -38.595 37.565 ;
        RECT -38.925 35.875 -38.595 36.205 ;
        RECT -38.925 34.515 -38.595 34.845 ;
        RECT -38.925 33.155 -38.595 33.485 ;
        RECT -38.925 31.795 -38.595 32.125 ;
        RECT -38.925 30.435 -38.595 30.765 ;
        RECT -38.925 29.075 -38.595 29.405 ;
        RECT -38.925 27.715 -38.595 28.045 ;
        RECT -38.925 26.355 -38.595 26.685 ;
        RECT -38.925 24.995 -38.595 25.325 ;
        RECT -38.925 23.635 -38.595 23.965 ;
        RECT -38.925 22.275 -38.595 22.605 ;
        RECT -38.925 20.915 -38.595 21.245 ;
        RECT -38.925 19.555 -38.595 19.885 ;
        RECT -38.925 18.195 -38.595 18.525 ;
        RECT -38.925 16.835 -38.595 17.165 ;
        RECT -38.925 15.475 -38.595 15.805 ;
        RECT -38.925 14.115 -38.595 14.445 ;
        RECT -38.925 12.755 -38.595 13.085 ;
        RECT -38.925 11.395 -38.595 11.725 ;
        RECT -38.925 10.035 -38.595 10.365 ;
        RECT -38.925 8.675 -38.595 9.005 ;
        RECT -38.925 7.315 -38.595 7.645 ;
        RECT -38.925 5.955 -38.595 6.285 ;
        RECT -38.925 4.595 -38.595 4.925 ;
        RECT -38.925 3.235 -38.595 3.565 ;
        RECT -38.925 1.875 -38.595 2.205 ;
        RECT -38.925 0.515 -38.595 0.845 ;
        RECT -38.925 -0.845 -38.595 -0.515 ;
        RECT -38.925 -2.205 -38.595 -1.875 ;
        RECT -38.925 -3.565 -38.595 -3.235 ;
        RECT -38.925 -4.925 -38.595 -4.595 ;
        RECT -38.925 -10.365 -38.595 -10.035 ;
        RECT -38.925 -14.445 -38.595 -14.115 ;
        RECT -38.925 -15.805 -38.595 -15.475 ;
        RECT -38.925 -17.165 -38.595 -16.835 ;
        RECT -38.925 -18.525 -38.595 -18.195 ;
        RECT -38.925 -19.885 -38.595 -19.555 ;
        RECT -38.925 -21.245 -38.595 -20.915 ;
        RECT -38.925 -22.605 -38.595 -22.275 ;
        RECT -38.925 -23.965 -38.595 -23.635 ;
        RECT -38.925 -25.325 -38.595 -24.995 ;
        RECT -38.925 -32.125 -38.595 -31.795 ;
        RECT -38.925 -33.71 -38.595 -33.38 ;
        RECT -38.925 -34.845 -38.595 -34.515 ;
        RECT -38.925 -36.205 -38.595 -35.875 ;
        RECT -38.925 -38.925 -38.595 -38.595 ;
        RECT -38.925 -39.75 -38.595 -39.42 ;
        RECT -38.925 -41.645 -38.595 -41.315 ;
        RECT -38.925 -44.365 -38.595 -44.035 ;
        RECT -38.925 -49.805 -38.595 -49.475 ;
        RECT -38.925 -51.165 -38.595 -50.835 ;
        RECT -38.925 -53.885 -38.595 -53.555 ;
        RECT -38.925 -55.245 -38.595 -54.915 ;
        RECT -38.925 -59.325 -38.595 -58.995 ;
        RECT -38.925 -60.685 -38.595 -60.355 ;
        RECT -38.925 -67.485 -38.595 -67.155 ;
        RECT -38.925 -70.205 -38.595 -69.875 ;
        RECT -38.925 -71.565 -38.595 -71.235 ;
        RECT -38.925 -72.925 -38.595 -72.595 ;
        RECT -38.925 -74.285 -38.595 -73.955 ;
        RECT -38.925 -75.645 -38.595 -75.315 ;
        RECT -38.925 -77.005 -38.595 -76.675 ;
        RECT -38.925 -78.365 -38.595 -78.035 ;
        RECT -38.925 -79.725 -38.595 -79.395 ;
        RECT -38.925 -81.085 -38.595 -80.755 ;
        RECT -38.925 -82.445 -38.595 -82.115 ;
        RECT -38.925 -83.805 -38.595 -83.475 ;
        RECT -38.925 -85.165 -38.595 -84.835 ;
        RECT -38.925 -86.525 -38.595 -86.195 ;
        RECT -38.925 -87.885 -38.595 -87.555 ;
        RECT -38.925 -89.245 -38.595 -88.915 ;
        RECT -38.925 -90.81 -38.595 -90.48 ;
        RECT -38.925 -91.965 -38.595 -91.635 ;
        RECT -38.925 -93.325 -38.595 -92.995 ;
        RECT -38.925 -94.685 -38.595 -94.355 ;
        RECT -38.925 -96.045 -38.595 -95.715 ;
        RECT -38.925 -97.405 -38.595 -97.075 ;
        RECT -38.925 -100.125 -38.595 -99.795 ;
        RECT -38.925 -101.35 -38.595 -101.02 ;
        RECT -38.925 -102.845 -38.595 -102.515 ;
        RECT -38.925 -104.205 -38.595 -103.875 ;
        RECT -38.925 -105.565 -38.595 -105.235 ;
        RECT -38.925 -108.285 -38.595 -107.955 ;
        RECT -38.925 -109.645 -38.595 -109.315 ;
        RECT -38.925 -112.365 -38.595 -112.035 ;
        RECT -38.925 -113.725 -38.595 -113.395 ;
        RECT -38.925 -115.085 -38.595 -114.755 ;
        RECT -38.925 -116.445 -38.595 -116.115 ;
        RECT -38.925 -117.805 -38.595 -117.475 ;
        RECT -38.925 -119.165 -38.595 -118.835 ;
        RECT -38.925 -120.525 -38.595 -120.195 ;
        RECT -38.925 -121.885 -38.595 -121.555 ;
        RECT -38.925 -123.245 -38.595 -122.915 ;
        RECT -38.925 -124.605 -38.595 -124.275 ;
        RECT -38.925 -125.965 -38.595 -125.635 ;
        RECT -38.925 -127.325 -38.595 -126.995 ;
        RECT -38.925 -128.685 -38.595 -128.355 ;
        RECT -38.925 -130.045 -38.595 -129.715 ;
        RECT -38.925 -132.765 -38.595 -132.435 ;
        RECT -38.925 -134.125 -38.595 -133.795 ;
        RECT -38.925 -135.485 -38.595 -135.155 ;
        RECT -38.925 -136.845 -38.595 -136.515 ;
        RECT -38.925 -138.205 -38.595 -137.875 ;
        RECT -38.925 -139.565 -38.595 -139.235 ;
        RECT -38.925 -140.925 -38.595 -140.595 ;
        RECT -38.925 -142.285 -38.595 -141.955 ;
        RECT -38.925 -143.645 -38.595 -143.315 ;
        RECT -38.925 -145.005 -38.595 -144.675 ;
        RECT -38.925 -146.365 -38.595 -146.035 ;
        RECT -38.925 -147.725 -38.595 -147.395 ;
        RECT -38.925 -150.445 -38.595 -150.115 ;
        RECT -38.925 -151.805 -38.595 -151.475 ;
        RECT -38.925 -154.525 -38.595 -154.195 ;
        RECT -38.925 -155.885 -38.595 -155.555 ;
        RECT -38.925 -157.245 -38.595 -156.915 ;
        RECT -38.925 -158.605 -38.595 -158.275 ;
        RECT -38.925 -159.965 -38.595 -159.635 ;
        RECT -38.925 -161.325 -38.595 -160.995 ;
        RECT -38.925 -162.685 -38.595 -162.355 ;
        RECT -38.925 -164.045 -38.595 -163.715 ;
        RECT -38.925 -165.405 -38.595 -165.075 ;
        RECT -38.925 -166.765 -38.595 -166.435 ;
        RECT -38.925 -168.655 -38.595 -168.325 ;
        RECT -38.925 -169.485 -38.595 -169.155 ;
        RECT -38.925 -170.845 -38.595 -170.515 ;
        RECT -38.925 -173.565 -38.595 -173.235 ;
        RECT -38.925 -174.925 -38.595 -174.595 ;
        RECT -38.925 -177.645 -38.595 -177.315 ;
        RECT -38.925 -183.29 -38.595 -182.16 ;
        RECT -38.92 -183.405 -38.6 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -37.565 244.04 -37.235 245.17 ;
        RECT -37.565 239.875 -37.235 240.205 ;
        RECT -37.565 238.515 -37.235 238.845 ;
        RECT -37.565 237.155 -37.235 237.485 ;
        RECT -37.565 235.795 -37.235 236.125 ;
        RECT -37.565 234.435 -37.235 234.765 ;
        RECT -37.565 233.075 -37.235 233.405 ;
        RECT -37.565 231.715 -37.235 232.045 ;
        RECT -37.565 230.355 -37.235 230.685 ;
        RECT -37.565 228.995 -37.235 229.325 ;
        RECT -37.565 227.635 -37.235 227.965 ;
        RECT -37.565 226.275 -37.235 226.605 ;
        RECT -37.565 224.915 -37.235 225.245 ;
        RECT -37.565 223.555 -37.235 223.885 ;
        RECT -37.565 222.195 -37.235 222.525 ;
        RECT -37.565 220.835 -37.235 221.165 ;
        RECT -37.565 219.475 -37.235 219.805 ;
        RECT -37.565 218.115 -37.235 218.445 ;
        RECT -37.565 216.755 -37.235 217.085 ;
        RECT -37.565 215.395 -37.235 215.725 ;
        RECT -37.565 214.035 -37.235 214.365 ;
        RECT -37.565 212.675 -37.235 213.005 ;
        RECT -37.565 211.315 -37.235 211.645 ;
        RECT -37.565 209.955 -37.235 210.285 ;
        RECT -37.565 208.595 -37.235 208.925 ;
        RECT -37.565 207.235 -37.235 207.565 ;
        RECT -37.565 205.875 -37.235 206.205 ;
        RECT -37.565 204.515 -37.235 204.845 ;
        RECT -37.565 203.155 -37.235 203.485 ;
        RECT -37.565 201.795 -37.235 202.125 ;
        RECT -37.565 200.435 -37.235 200.765 ;
        RECT -37.565 199.075 -37.235 199.405 ;
        RECT -37.565 197.715 -37.235 198.045 ;
        RECT -37.565 196.355 -37.235 196.685 ;
        RECT -37.565 194.995 -37.235 195.325 ;
        RECT -37.565 193.635 -37.235 193.965 ;
        RECT -37.565 192.275 -37.235 192.605 ;
        RECT -37.565 190.915 -37.235 191.245 ;
        RECT -37.565 189.555 -37.235 189.885 ;
        RECT -37.565 188.195 -37.235 188.525 ;
        RECT -37.565 186.835 -37.235 187.165 ;
        RECT -37.565 185.475 -37.235 185.805 ;
        RECT -37.565 184.115 -37.235 184.445 ;
        RECT -37.565 182.755 -37.235 183.085 ;
        RECT -37.565 181.395 -37.235 181.725 ;
        RECT -37.565 180.035 -37.235 180.365 ;
        RECT -37.565 178.675 -37.235 179.005 ;
        RECT -37.565 177.315 -37.235 177.645 ;
        RECT -37.565 175.955 -37.235 176.285 ;
        RECT -37.565 174.595 -37.235 174.925 ;
        RECT -37.565 173.235 -37.235 173.565 ;
        RECT -37.565 171.875 -37.235 172.205 ;
        RECT -37.565 170.515 -37.235 170.845 ;
        RECT -37.565 169.155 -37.235 169.485 ;
        RECT -37.565 167.795 -37.235 168.125 ;
        RECT -37.565 166.435 -37.235 166.765 ;
        RECT -37.565 165.075 -37.235 165.405 ;
        RECT -37.565 163.715 -37.235 164.045 ;
        RECT -37.565 162.355 -37.235 162.685 ;
        RECT -37.565 160.995 -37.235 161.325 ;
        RECT -37.565 159.635 -37.235 159.965 ;
        RECT -37.565 158.275 -37.235 158.605 ;
        RECT -37.565 156.915 -37.235 157.245 ;
        RECT -37.565 155.555 -37.235 155.885 ;
        RECT -37.565 154.195 -37.235 154.525 ;
        RECT -37.565 152.835 -37.235 153.165 ;
        RECT -37.565 151.475 -37.235 151.805 ;
        RECT -37.565 150.115 -37.235 150.445 ;
        RECT -37.565 148.755 -37.235 149.085 ;
        RECT -37.565 147.395 -37.235 147.725 ;
        RECT -37.565 146.035 -37.235 146.365 ;
        RECT -37.565 144.675 -37.235 145.005 ;
        RECT -37.565 143.315 -37.235 143.645 ;
        RECT -37.565 141.955 -37.235 142.285 ;
        RECT -37.565 140.595 -37.235 140.925 ;
        RECT -37.565 139.235 -37.235 139.565 ;
        RECT -37.565 137.875 -37.235 138.205 ;
        RECT -37.565 136.515 -37.235 136.845 ;
        RECT -37.565 135.155 -37.235 135.485 ;
        RECT -37.565 133.795 -37.235 134.125 ;
        RECT -37.565 132.435 -37.235 132.765 ;
        RECT -37.565 131.075 -37.235 131.405 ;
        RECT -37.565 129.715 -37.235 130.045 ;
        RECT -37.565 128.355 -37.235 128.685 ;
        RECT -37.565 126.995 -37.235 127.325 ;
        RECT -37.565 125.635 -37.235 125.965 ;
        RECT -37.565 124.275 -37.235 124.605 ;
        RECT -37.565 122.915 -37.235 123.245 ;
        RECT -37.565 121.555 -37.235 121.885 ;
        RECT -37.565 120.195 -37.235 120.525 ;
        RECT -37.565 118.835 -37.235 119.165 ;
        RECT -37.565 117.475 -37.235 117.805 ;
        RECT -37.565 116.115 -37.235 116.445 ;
        RECT -37.565 114.755 -37.235 115.085 ;
        RECT -37.565 113.395 -37.235 113.725 ;
        RECT -37.565 112.035 -37.235 112.365 ;
        RECT -37.565 110.675 -37.235 111.005 ;
        RECT -37.565 109.315 -37.235 109.645 ;
        RECT -37.565 107.955 -37.235 108.285 ;
        RECT -37.565 106.595 -37.235 106.925 ;
        RECT -37.565 105.235 -37.235 105.565 ;
        RECT -37.565 103.875 -37.235 104.205 ;
        RECT -37.565 102.515 -37.235 102.845 ;
        RECT -37.565 101.155 -37.235 101.485 ;
        RECT -37.565 99.795 -37.235 100.125 ;
        RECT -37.565 98.435 -37.235 98.765 ;
        RECT -37.565 97.075 -37.235 97.405 ;
        RECT -37.565 95.715 -37.235 96.045 ;
        RECT -37.565 94.355 -37.235 94.685 ;
        RECT -37.565 92.995 -37.235 93.325 ;
        RECT -37.565 91.635 -37.235 91.965 ;
        RECT -37.565 90.275 -37.235 90.605 ;
        RECT -37.565 88.915 -37.235 89.245 ;
        RECT -37.565 87.555 -37.235 87.885 ;
        RECT -37.565 86.195 -37.235 86.525 ;
        RECT -37.565 84.835 -37.235 85.165 ;
        RECT -37.565 83.475 -37.235 83.805 ;
        RECT -37.565 82.115 -37.235 82.445 ;
        RECT -37.565 80.755 -37.235 81.085 ;
        RECT -37.565 79.395 -37.235 79.725 ;
        RECT -37.565 78.035 -37.235 78.365 ;
        RECT -37.565 76.675 -37.235 77.005 ;
        RECT -37.565 75.315 -37.235 75.645 ;
        RECT -37.565 73.955 -37.235 74.285 ;
        RECT -37.565 72.595 -37.235 72.925 ;
        RECT -37.565 71.235 -37.235 71.565 ;
        RECT -37.565 69.875 -37.235 70.205 ;
        RECT -37.565 68.515 -37.235 68.845 ;
        RECT -37.565 67.155 -37.235 67.485 ;
        RECT -37.565 65.795 -37.235 66.125 ;
        RECT -37.565 64.435 -37.235 64.765 ;
        RECT -37.565 63.075 -37.235 63.405 ;
        RECT -37.565 61.715 -37.235 62.045 ;
        RECT -37.565 60.355 -37.235 60.685 ;
        RECT -37.565 58.995 -37.235 59.325 ;
        RECT -37.565 57.635 -37.235 57.965 ;
        RECT -37.565 56.275 -37.235 56.605 ;
        RECT -37.565 54.915 -37.235 55.245 ;
        RECT -37.565 53.555 -37.235 53.885 ;
        RECT -37.565 52.195 -37.235 52.525 ;
        RECT -37.565 50.835 -37.235 51.165 ;
        RECT -37.565 49.475 -37.235 49.805 ;
        RECT -37.565 48.115 -37.235 48.445 ;
        RECT -37.565 46.755 -37.235 47.085 ;
        RECT -37.565 45.395 -37.235 45.725 ;
        RECT -37.565 44.035 -37.235 44.365 ;
        RECT -37.565 42.675 -37.235 43.005 ;
        RECT -37.565 41.315 -37.235 41.645 ;
        RECT -37.565 39.955 -37.235 40.285 ;
        RECT -37.565 38.595 -37.235 38.925 ;
        RECT -37.565 37.235 -37.235 37.565 ;
        RECT -37.565 35.875 -37.235 36.205 ;
        RECT -37.565 34.515 -37.235 34.845 ;
        RECT -37.565 33.155 -37.235 33.485 ;
        RECT -37.565 31.795 -37.235 32.125 ;
        RECT -37.565 30.435 -37.235 30.765 ;
        RECT -37.565 29.075 -37.235 29.405 ;
        RECT -37.565 27.715 -37.235 28.045 ;
        RECT -37.565 26.355 -37.235 26.685 ;
        RECT -37.565 24.995 -37.235 25.325 ;
        RECT -37.565 23.635 -37.235 23.965 ;
        RECT -37.565 22.275 -37.235 22.605 ;
        RECT -37.565 20.915 -37.235 21.245 ;
        RECT -37.565 19.555 -37.235 19.885 ;
        RECT -37.565 18.195 -37.235 18.525 ;
        RECT -37.565 16.835 -37.235 17.165 ;
        RECT -37.565 15.475 -37.235 15.805 ;
        RECT -37.565 14.115 -37.235 14.445 ;
        RECT -37.565 12.755 -37.235 13.085 ;
        RECT -37.565 11.395 -37.235 11.725 ;
        RECT -37.565 10.035 -37.235 10.365 ;
        RECT -37.565 8.675 -37.235 9.005 ;
        RECT -37.565 7.315 -37.235 7.645 ;
        RECT -37.565 5.955 -37.235 6.285 ;
        RECT -37.565 4.595 -37.235 4.925 ;
        RECT -37.565 3.235 -37.235 3.565 ;
        RECT -37.565 1.875 -37.235 2.205 ;
        RECT -37.565 0.515 -37.235 0.845 ;
        RECT -37.565 -0.845 -37.235 -0.515 ;
        RECT -37.565 -2.205 -37.235 -1.875 ;
        RECT -37.565 -3.565 -37.235 -3.235 ;
        RECT -37.565 -10.365 -37.235 -10.035 ;
        RECT -37.565 -14.445 -37.235 -14.115 ;
        RECT -37.565 -15.805 -37.235 -15.475 ;
        RECT -37.565 -17.165 -37.235 -16.835 ;
        RECT -37.565 -18.525 -37.235 -18.195 ;
        RECT -37.565 -19.885 -37.235 -19.555 ;
        RECT -37.565 -21.245 -37.235 -20.915 ;
        RECT -37.565 -22.605 -37.235 -22.275 ;
        RECT -37.565 -23.965 -37.235 -23.635 ;
        RECT -37.565 -25.325 -37.235 -24.995 ;
        RECT -37.565 -32.125 -37.235 -31.795 ;
        RECT -37.565 -33.71 -37.235 -33.38 ;
        RECT -37.565 -34.845 -37.235 -34.515 ;
        RECT -37.565 -36.205 -37.235 -35.875 ;
        RECT -37.565 -38.925 -37.235 -38.595 ;
        RECT -37.565 -39.75 -37.235 -39.42 ;
        RECT -37.565 -41.645 -37.235 -41.315 ;
        RECT -37.565 -44.365 -37.235 -44.035 ;
        RECT -37.565 -49.805 -37.235 -49.475 ;
        RECT -37.565 -51.165 -37.235 -50.835 ;
        RECT -37.565 -52.525 -37.235 -52.195 ;
        RECT -37.565 -53.885 -37.235 -53.555 ;
        RECT -37.565 -55.245 -37.235 -54.915 ;
        RECT -37.565 -56.605 -37.235 -56.275 ;
        RECT -37.565 -57.965 -37.235 -57.635 ;
        RECT -37.565 -59.325 -37.235 -58.995 ;
        RECT -37.565 -60.685 -37.235 -60.355 ;
        RECT -37.565 -62.045 -37.235 -61.715 ;
        RECT -37.565 -64.765 -37.235 -64.435 ;
        RECT -37.565 -66.125 -37.235 -65.795 ;
        RECT -37.565 -67.485 -37.235 -67.155 ;
        RECT -37.565 -68.845 -37.235 -68.515 ;
        RECT -37.565 -70.205 -37.235 -69.875 ;
        RECT -37.565 -71.565 -37.235 -71.235 ;
        RECT -37.565 -72.925 -37.235 -72.595 ;
        RECT -37.565 -74.285 -37.235 -73.955 ;
        RECT -37.565 -75.645 -37.235 -75.315 ;
        RECT -37.565 -77.005 -37.235 -76.675 ;
        RECT -37.565 -78.365 -37.235 -78.035 ;
        RECT -37.565 -79.725 -37.235 -79.395 ;
        RECT -37.565 -81.085 -37.235 -80.755 ;
        RECT -37.565 -82.445 -37.235 -82.115 ;
        RECT -37.565 -83.805 -37.235 -83.475 ;
        RECT -37.565 -85.165 -37.235 -84.835 ;
        RECT -37.565 -86.525 -37.235 -86.195 ;
        RECT -37.565 -87.885 -37.235 -87.555 ;
        RECT -37.565 -89.245 -37.235 -88.915 ;
        RECT -37.565 -90.81 -37.235 -90.48 ;
        RECT -37.565 -91.965 -37.235 -91.635 ;
        RECT -37.565 -93.325 -37.235 -92.995 ;
        RECT -37.565 -94.685 -37.235 -94.355 ;
        RECT -37.565 -96.045 -37.235 -95.715 ;
        RECT -37.565 -97.405 -37.235 -97.075 ;
        RECT -37.565 -100.125 -37.235 -99.795 ;
        RECT -37.565 -101.35 -37.235 -101.02 ;
        RECT -37.565 -102.845 -37.235 -102.515 ;
        RECT -37.565 -104.205 -37.235 -103.875 ;
        RECT -37.565 -105.565 -37.235 -105.235 ;
        RECT -37.565 -108.285 -37.235 -107.955 ;
        RECT -37.565 -109.645 -37.235 -109.315 ;
        RECT -37.565 -112.365 -37.235 -112.035 ;
        RECT -37.565 -113.725 -37.235 -113.395 ;
        RECT -37.565 -115.085 -37.235 -114.755 ;
        RECT -37.565 -116.445 -37.235 -116.115 ;
        RECT -37.565 -117.805 -37.235 -117.475 ;
        RECT -37.565 -119.165 -37.235 -118.835 ;
        RECT -37.565 -120.525 -37.235 -120.195 ;
        RECT -37.565 -121.885 -37.235 -121.555 ;
        RECT -37.565 -123.245 -37.235 -122.915 ;
        RECT -37.565 -124.605 -37.235 -124.275 ;
        RECT -37.565 -125.965 -37.235 -125.635 ;
        RECT -37.565 -127.325 -37.235 -126.995 ;
        RECT -37.565 -128.685 -37.235 -128.355 ;
        RECT -37.565 -132.765 -37.235 -132.435 ;
        RECT -37.565 -134.125 -37.235 -133.795 ;
        RECT -37.565 -135.485 -37.235 -135.155 ;
        RECT -37.565 -136.845 -37.235 -136.515 ;
        RECT -37.565 -138.205 -37.235 -137.875 ;
        RECT -37.565 -139.565 -37.235 -139.235 ;
        RECT -37.565 -140.925 -37.235 -140.595 ;
        RECT -37.565 -142.285 -37.235 -141.955 ;
        RECT -37.565 -143.645 -37.235 -143.315 ;
        RECT -37.565 -145.005 -37.235 -144.675 ;
        RECT -37.565 -146.365 -37.235 -146.035 ;
        RECT -37.565 -147.725 -37.235 -147.395 ;
        RECT -37.565 -150.445 -37.235 -150.115 ;
        RECT -37.565 -151.805 -37.235 -151.475 ;
        RECT -37.565 -155.885 -37.235 -155.555 ;
        RECT -37.565 -157.245 -37.235 -156.915 ;
        RECT -37.565 -158.605 -37.235 -158.275 ;
        RECT -37.565 -159.965 -37.235 -159.635 ;
        RECT -37.565 -161.325 -37.235 -160.995 ;
        RECT -37.565 -162.685 -37.235 -162.355 ;
        RECT -37.565 -164.045 -37.235 -163.715 ;
        RECT -37.565 -165.405 -37.235 -165.075 ;
        RECT -37.565 -166.765 -37.235 -166.435 ;
        RECT -37.565 -168.655 -37.235 -168.325 ;
        RECT -37.565 -169.485 -37.235 -169.155 ;
        RECT -37.565 -170.845 -37.235 -170.515 ;
        RECT -37.565 -172.205 -37.235 -171.875 ;
        RECT -37.565 -173.565 -37.235 -173.235 ;
        RECT -37.565 -174.925 -37.235 -174.595 ;
        RECT -37.565 -177.645 -37.235 -177.315 ;
        RECT -37.565 -183.29 -37.235 -182.16 ;
        RECT -37.56 -183.405 -37.24 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -36.205 -101.35 -35.875 -101.02 ;
        RECT -36.205 -102.845 -35.875 -102.515 ;
        RECT -36.205 -104.205 -35.875 -103.875 ;
        RECT -36.205 -105.565 -35.875 -105.235 ;
        RECT -36.205 -108.285 -35.875 -107.955 ;
        RECT -36.205 -109.645 -35.875 -109.315 ;
        RECT -36.205 -112.365 -35.875 -112.035 ;
        RECT -36.205 -113.725 -35.875 -113.395 ;
        RECT -36.205 -115.085 -35.875 -114.755 ;
        RECT -36.205 -116.445 -35.875 -116.115 ;
        RECT -36.205 -117.805 -35.875 -117.475 ;
        RECT -36.205 -119.165 -35.875 -118.835 ;
        RECT -36.205 -120.525 -35.875 -120.195 ;
        RECT -36.205 -121.885 -35.875 -121.555 ;
        RECT -36.205 -123.245 -35.875 -122.915 ;
        RECT -36.205 -124.605 -35.875 -124.275 ;
        RECT -36.205 -125.965 -35.875 -125.635 ;
        RECT -36.205 -127.325 -35.875 -126.995 ;
        RECT -36.205 -128.685 -35.875 -128.355 ;
        RECT -36.205 -132.765 -35.875 -132.435 ;
        RECT -36.205 -134.125 -35.875 -133.795 ;
        RECT -36.205 -135.485 -35.875 -135.155 ;
        RECT -36.205 -136.845 -35.875 -136.515 ;
        RECT -36.205 -138.205 -35.875 -137.875 ;
        RECT -36.205 -139.565 -35.875 -139.235 ;
        RECT -36.205 -140.925 -35.875 -140.595 ;
        RECT -36.205 -142.285 -35.875 -141.955 ;
        RECT -36.205 -143.645 -35.875 -143.315 ;
        RECT -36.205 -145.005 -35.875 -144.675 ;
        RECT -36.205 -146.365 -35.875 -146.035 ;
        RECT -36.205 -147.725 -35.875 -147.395 ;
        RECT -36.205 -150.445 -35.875 -150.115 ;
        RECT -36.205 -151.805 -35.875 -151.475 ;
        RECT -36.205 -155.885 -35.875 -155.555 ;
        RECT -36.205 -157.245 -35.875 -156.915 ;
        RECT -36.205 -158.605 -35.875 -158.275 ;
        RECT -36.205 -159.965 -35.875 -159.635 ;
        RECT -36.205 -161.325 -35.875 -160.995 ;
        RECT -36.205 -162.685 -35.875 -162.355 ;
        RECT -36.205 -164.045 -35.875 -163.715 ;
        RECT -36.205 -165.405 -35.875 -165.075 ;
        RECT -36.205 -166.765 -35.875 -166.435 ;
        RECT -36.205 -168.655 -35.875 -168.325 ;
        RECT -36.205 -169.485 -35.875 -169.155 ;
        RECT -36.205 -170.845 -35.875 -170.515 ;
        RECT -36.205 -172.205 -35.875 -171.875 ;
        RECT -36.205 -174.925 -35.875 -174.595 ;
        RECT -36.205 -177.645 -35.875 -177.315 ;
        RECT -36.205 -183.29 -35.875 -182.16 ;
        RECT -36.2 -183.405 -35.88 245.285 ;
        RECT -36.205 244.04 -35.875 245.17 ;
        RECT -36.205 239.875 -35.875 240.205 ;
        RECT -36.205 238.515 -35.875 238.845 ;
        RECT -36.205 237.155 -35.875 237.485 ;
        RECT -36.205 235.795 -35.875 236.125 ;
        RECT -36.205 234.435 -35.875 234.765 ;
        RECT -36.205 233.075 -35.875 233.405 ;
        RECT -36.205 231.715 -35.875 232.045 ;
        RECT -36.205 230.355 -35.875 230.685 ;
        RECT -36.205 228.995 -35.875 229.325 ;
        RECT -36.205 227.635 -35.875 227.965 ;
        RECT -36.205 226.275 -35.875 226.605 ;
        RECT -36.205 224.915 -35.875 225.245 ;
        RECT -36.205 223.555 -35.875 223.885 ;
        RECT -36.205 222.195 -35.875 222.525 ;
        RECT -36.205 220.835 -35.875 221.165 ;
        RECT -36.205 219.475 -35.875 219.805 ;
        RECT -36.205 218.115 -35.875 218.445 ;
        RECT -36.205 216.755 -35.875 217.085 ;
        RECT -36.205 215.395 -35.875 215.725 ;
        RECT -36.205 214.035 -35.875 214.365 ;
        RECT -36.205 212.675 -35.875 213.005 ;
        RECT -36.205 211.315 -35.875 211.645 ;
        RECT -36.205 209.955 -35.875 210.285 ;
        RECT -36.205 208.595 -35.875 208.925 ;
        RECT -36.205 207.235 -35.875 207.565 ;
        RECT -36.205 205.875 -35.875 206.205 ;
        RECT -36.205 204.515 -35.875 204.845 ;
        RECT -36.205 203.155 -35.875 203.485 ;
        RECT -36.205 201.795 -35.875 202.125 ;
        RECT -36.205 200.435 -35.875 200.765 ;
        RECT -36.205 199.075 -35.875 199.405 ;
        RECT -36.205 197.715 -35.875 198.045 ;
        RECT -36.205 196.355 -35.875 196.685 ;
        RECT -36.205 194.995 -35.875 195.325 ;
        RECT -36.205 193.635 -35.875 193.965 ;
        RECT -36.205 192.275 -35.875 192.605 ;
        RECT -36.205 190.915 -35.875 191.245 ;
        RECT -36.205 189.555 -35.875 189.885 ;
        RECT -36.205 188.195 -35.875 188.525 ;
        RECT -36.205 186.835 -35.875 187.165 ;
        RECT -36.205 185.475 -35.875 185.805 ;
        RECT -36.205 184.115 -35.875 184.445 ;
        RECT -36.205 182.755 -35.875 183.085 ;
        RECT -36.205 181.395 -35.875 181.725 ;
        RECT -36.205 180.035 -35.875 180.365 ;
        RECT -36.205 178.675 -35.875 179.005 ;
        RECT -36.205 177.315 -35.875 177.645 ;
        RECT -36.205 175.955 -35.875 176.285 ;
        RECT -36.205 174.595 -35.875 174.925 ;
        RECT -36.205 173.235 -35.875 173.565 ;
        RECT -36.205 171.875 -35.875 172.205 ;
        RECT -36.205 170.515 -35.875 170.845 ;
        RECT -36.205 169.155 -35.875 169.485 ;
        RECT -36.205 167.795 -35.875 168.125 ;
        RECT -36.205 166.435 -35.875 166.765 ;
        RECT -36.205 165.075 -35.875 165.405 ;
        RECT -36.205 163.715 -35.875 164.045 ;
        RECT -36.205 162.355 -35.875 162.685 ;
        RECT -36.205 160.995 -35.875 161.325 ;
        RECT -36.205 159.635 -35.875 159.965 ;
        RECT -36.205 158.275 -35.875 158.605 ;
        RECT -36.205 156.915 -35.875 157.245 ;
        RECT -36.205 155.555 -35.875 155.885 ;
        RECT -36.205 154.195 -35.875 154.525 ;
        RECT -36.205 152.835 -35.875 153.165 ;
        RECT -36.205 151.475 -35.875 151.805 ;
        RECT -36.205 150.115 -35.875 150.445 ;
        RECT -36.205 148.755 -35.875 149.085 ;
        RECT -36.205 147.395 -35.875 147.725 ;
        RECT -36.205 146.035 -35.875 146.365 ;
        RECT -36.205 144.675 -35.875 145.005 ;
        RECT -36.205 143.315 -35.875 143.645 ;
        RECT -36.205 141.955 -35.875 142.285 ;
        RECT -36.205 140.595 -35.875 140.925 ;
        RECT -36.205 139.235 -35.875 139.565 ;
        RECT -36.205 137.875 -35.875 138.205 ;
        RECT -36.205 136.515 -35.875 136.845 ;
        RECT -36.205 135.155 -35.875 135.485 ;
        RECT -36.205 133.795 -35.875 134.125 ;
        RECT -36.205 132.435 -35.875 132.765 ;
        RECT -36.205 131.075 -35.875 131.405 ;
        RECT -36.205 129.715 -35.875 130.045 ;
        RECT -36.205 128.355 -35.875 128.685 ;
        RECT -36.205 126.995 -35.875 127.325 ;
        RECT -36.205 125.635 -35.875 125.965 ;
        RECT -36.205 124.275 -35.875 124.605 ;
        RECT -36.205 122.915 -35.875 123.245 ;
        RECT -36.205 121.555 -35.875 121.885 ;
        RECT -36.205 120.195 -35.875 120.525 ;
        RECT -36.205 118.835 -35.875 119.165 ;
        RECT -36.205 117.475 -35.875 117.805 ;
        RECT -36.205 116.115 -35.875 116.445 ;
        RECT -36.205 114.755 -35.875 115.085 ;
        RECT -36.205 113.395 -35.875 113.725 ;
        RECT -36.205 112.035 -35.875 112.365 ;
        RECT -36.205 110.675 -35.875 111.005 ;
        RECT -36.205 109.315 -35.875 109.645 ;
        RECT -36.205 107.955 -35.875 108.285 ;
        RECT -36.205 106.595 -35.875 106.925 ;
        RECT -36.205 105.235 -35.875 105.565 ;
        RECT -36.205 103.875 -35.875 104.205 ;
        RECT -36.205 102.515 -35.875 102.845 ;
        RECT -36.205 101.155 -35.875 101.485 ;
        RECT -36.205 99.795 -35.875 100.125 ;
        RECT -36.205 98.435 -35.875 98.765 ;
        RECT -36.205 97.075 -35.875 97.405 ;
        RECT -36.205 95.715 -35.875 96.045 ;
        RECT -36.205 94.355 -35.875 94.685 ;
        RECT -36.205 92.995 -35.875 93.325 ;
        RECT -36.205 91.635 -35.875 91.965 ;
        RECT -36.205 90.275 -35.875 90.605 ;
        RECT -36.205 88.915 -35.875 89.245 ;
        RECT -36.205 87.555 -35.875 87.885 ;
        RECT -36.205 86.195 -35.875 86.525 ;
        RECT -36.205 84.835 -35.875 85.165 ;
        RECT -36.205 83.475 -35.875 83.805 ;
        RECT -36.205 82.115 -35.875 82.445 ;
        RECT -36.205 80.755 -35.875 81.085 ;
        RECT -36.205 79.395 -35.875 79.725 ;
        RECT -36.205 78.035 -35.875 78.365 ;
        RECT -36.205 76.675 -35.875 77.005 ;
        RECT -36.205 75.315 -35.875 75.645 ;
        RECT -36.205 73.955 -35.875 74.285 ;
        RECT -36.205 72.595 -35.875 72.925 ;
        RECT -36.205 71.235 -35.875 71.565 ;
        RECT -36.205 69.875 -35.875 70.205 ;
        RECT -36.205 68.515 -35.875 68.845 ;
        RECT -36.205 67.155 -35.875 67.485 ;
        RECT -36.205 65.795 -35.875 66.125 ;
        RECT -36.205 64.435 -35.875 64.765 ;
        RECT -36.205 63.075 -35.875 63.405 ;
        RECT -36.205 61.715 -35.875 62.045 ;
        RECT -36.205 60.355 -35.875 60.685 ;
        RECT -36.205 58.995 -35.875 59.325 ;
        RECT -36.205 57.635 -35.875 57.965 ;
        RECT -36.205 56.275 -35.875 56.605 ;
        RECT -36.205 54.915 -35.875 55.245 ;
        RECT -36.205 53.555 -35.875 53.885 ;
        RECT -36.205 52.195 -35.875 52.525 ;
        RECT -36.205 50.835 -35.875 51.165 ;
        RECT -36.205 49.475 -35.875 49.805 ;
        RECT -36.205 48.115 -35.875 48.445 ;
        RECT -36.205 46.755 -35.875 47.085 ;
        RECT -36.205 45.395 -35.875 45.725 ;
        RECT -36.205 44.035 -35.875 44.365 ;
        RECT -36.205 42.675 -35.875 43.005 ;
        RECT -36.205 41.315 -35.875 41.645 ;
        RECT -36.205 39.955 -35.875 40.285 ;
        RECT -36.205 38.595 -35.875 38.925 ;
        RECT -36.205 37.235 -35.875 37.565 ;
        RECT -36.205 35.875 -35.875 36.205 ;
        RECT -36.205 34.515 -35.875 34.845 ;
        RECT -36.205 33.155 -35.875 33.485 ;
        RECT -36.205 31.795 -35.875 32.125 ;
        RECT -36.205 30.435 -35.875 30.765 ;
        RECT -36.205 29.075 -35.875 29.405 ;
        RECT -36.205 27.715 -35.875 28.045 ;
        RECT -36.205 26.355 -35.875 26.685 ;
        RECT -36.205 24.995 -35.875 25.325 ;
        RECT -36.205 23.635 -35.875 23.965 ;
        RECT -36.205 22.275 -35.875 22.605 ;
        RECT -36.205 20.915 -35.875 21.245 ;
        RECT -36.205 19.555 -35.875 19.885 ;
        RECT -36.205 18.195 -35.875 18.525 ;
        RECT -36.205 16.835 -35.875 17.165 ;
        RECT -36.205 15.475 -35.875 15.805 ;
        RECT -36.205 14.115 -35.875 14.445 ;
        RECT -36.205 12.755 -35.875 13.085 ;
        RECT -36.205 11.395 -35.875 11.725 ;
        RECT -36.205 10.035 -35.875 10.365 ;
        RECT -36.205 8.675 -35.875 9.005 ;
        RECT -36.205 7.315 -35.875 7.645 ;
        RECT -36.205 5.955 -35.875 6.285 ;
        RECT -36.205 4.595 -35.875 4.925 ;
        RECT -36.205 3.235 -35.875 3.565 ;
        RECT -36.205 1.875 -35.875 2.205 ;
        RECT -36.205 0.515 -35.875 0.845 ;
        RECT -36.205 -0.845 -35.875 -0.515 ;
        RECT -36.205 -2.205 -35.875 -1.875 ;
        RECT -36.205 -7.645 -35.875 -7.315 ;
        RECT -36.205 -10.365 -35.875 -10.035 ;
        RECT -36.205 -14.445 -35.875 -14.115 ;
        RECT -36.205 -15.805 -35.875 -15.475 ;
        RECT -36.205 -17.165 -35.875 -16.835 ;
        RECT -36.205 -18.525 -35.875 -18.195 ;
        RECT -36.205 -19.885 -35.875 -19.555 ;
        RECT -36.205 -21.245 -35.875 -20.915 ;
        RECT -36.205 -22.605 -35.875 -22.275 ;
        RECT -36.205 -23.965 -35.875 -23.635 ;
        RECT -36.205 -25.325 -35.875 -24.995 ;
        RECT -36.205 -32.125 -35.875 -31.795 ;
        RECT -36.205 -33.71 -35.875 -33.38 ;
        RECT -36.205 -34.845 -35.875 -34.515 ;
        RECT -36.205 -36.205 -35.875 -35.875 ;
        RECT -36.205 -38.925 -35.875 -38.595 ;
        RECT -36.205 -39.75 -35.875 -39.42 ;
        RECT -36.205 -41.645 -35.875 -41.315 ;
        RECT -36.205 -44.365 -35.875 -44.035 ;
        RECT -36.205 -49.805 -35.875 -49.475 ;
        RECT -36.205 -51.165 -35.875 -50.835 ;
        RECT -36.205 -52.525 -35.875 -52.195 ;
        RECT -36.205 -53.885 -35.875 -53.555 ;
        RECT -36.205 -55.245 -35.875 -54.915 ;
        RECT -36.205 -56.605 -35.875 -56.275 ;
        RECT -36.205 -57.965 -35.875 -57.635 ;
        RECT -36.205 -59.325 -35.875 -58.995 ;
        RECT -36.205 -60.685 -35.875 -60.355 ;
        RECT -36.205 -62.045 -35.875 -61.715 ;
        RECT -36.205 -64.765 -35.875 -64.435 ;
        RECT -36.205 -66.125 -35.875 -65.795 ;
        RECT -36.205 -67.485 -35.875 -67.155 ;
        RECT -36.205 -68.845 -35.875 -68.515 ;
        RECT -36.205 -70.205 -35.875 -69.875 ;
        RECT -36.205 -71.565 -35.875 -71.235 ;
        RECT -36.205 -72.925 -35.875 -72.595 ;
        RECT -36.205 -74.285 -35.875 -73.955 ;
        RECT -36.205 -75.645 -35.875 -75.315 ;
        RECT -36.205 -77.005 -35.875 -76.675 ;
        RECT -36.205 -78.365 -35.875 -78.035 ;
        RECT -36.205 -79.725 -35.875 -79.395 ;
        RECT -36.205 -81.085 -35.875 -80.755 ;
        RECT -36.205 -82.445 -35.875 -82.115 ;
        RECT -36.205 -83.805 -35.875 -83.475 ;
        RECT -36.205 -85.165 -35.875 -84.835 ;
        RECT -36.205 -86.525 -35.875 -86.195 ;
        RECT -36.205 -87.885 -35.875 -87.555 ;
        RECT -36.205 -89.245 -35.875 -88.915 ;
        RECT -36.205 -90.81 -35.875 -90.48 ;
        RECT -36.205 -91.965 -35.875 -91.635 ;
        RECT -36.205 -93.325 -35.875 -92.995 ;
        RECT -36.205 -94.685 -35.875 -94.355 ;
        RECT -36.205 -96.045 -35.875 -95.715 ;
        RECT -36.205 -97.405 -35.875 -97.075 ;
        RECT -36.205 -100.125 -35.875 -99.795 ;
    END
    PORT
      LAYER met3 ;
        RECT -45.725 244.04 -45.395 245.17 ;
        RECT -45.725 239.875 -45.395 240.205 ;
        RECT -45.725 238.515 -45.395 238.845 ;
        RECT -45.725 237.155 -45.395 237.485 ;
        RECT -45.725 235.795 -45.395 236.125 ;
        RECT -45.725 234.435 -45.395 234.765 ;
        RECT -45.725 233.075 -45.395 233.405 ;
        RECT -45.725 231.715 -45.395 232.045 ;
        RECT -45.725 230.355 -45.395 230.685 ;
        RECT -45.725 228.995 -45.395 229.325 ;
        RECT -45.725 227.635 -45.395 227.965 ;
        RECT -45.725 226.275 -45.395 226.605 ;
        RECT -45.725 224.915 -45.395 225.245 ;
        RECT -45.725 223.555 -45.395 223.885 ;
        RECT -45.725 222.195 -45.395 222.525 ;
        RECT -45.725 220.835 -45.395 221.165 ;
        RECT -45.725 219.475 -45.395 219.805 ;
        RECT -45.725 218.115 -45.395 218.445 ;
        RECT -45.725 216.755 -45.395 217.085 ;
        RECT -45.725 215.395 -45.395 215.725 ;
        RECT -45.725 214.035 -45.395 214.365 ;
        RECT -45.725 212.675 -45.395 213.005 ;
        RECT -45.725 211.315 -45.395 211.645 ;
        RECT -45.725 209.955 -45.395 210.285 ;
        RECT -45.725 208.595 -45.395 208.925 ;
        RECT -45.725 207.235 -45.395 207.565 ;
        RECT -45.725 205.875 -45.395 206.205 ;
        RECT -45.725 204.515 -45.395 204.845 ;
        RECT -45.725 203.155 -45.395 203.485 ;
        RECT -45.725 201.795 -45.395 202.125 ;
        RECT -45.725 200.435 -45.395 200.765 ;
        RECT -45.725 199.075 -45.395 199.405 ;
        RECT -45.725 197.715 -45.395 198.045 ;
        RECT -45.725 196.355 -45.395 196.685 ;
        RECT -45.725 194.995 -45.395 195.325 ;
        RECT -45.725 193.635 -45.395 193.965 ;
        RECT -45.725 192.275 -45.395 192.605 ;
        RECT -45.725 190.915 -45.395 191.245 ;
        RECT -45.725 189.555 -45.395 189.885 ;
        RECT -45.725 188.195 -45.395 188.525 ;
        RECT -45.725 186.835 -45.395 187.165 ;
        RECT -45.725 185.475 -45.395 185.805 ;
        RECT -45.725 184.115 -45.395 184.445 ;
        RECT -45.725 182.755 -45.395 183.085 ;
        RECT -45.725 181.395 -45.395 181.725 ;
        RECT -45.725 180.035 -45.395 180.365 ;
        RECT -45.725 178.675 -45.395 179.005 ;
        RECT -45.725 177.315 -45.395 177.645 ;
        RECT -45.725 175.955 -45.395 176.285 ;
        RECT -45.725 174.595 -45.395 174.925 ;
        RECT -45.725 173.235 -45.395 173.565 ;
        RECT -45.725 171.875 -45.395 172.205 ;
        RECT -45.725 170.515 -45.395 170.845 ;
        RECT -45.725 169.155 -45.395 169.485 ;
        RECT -45.725 167.795 -45.395 168.125 ;
        RECT -45.725 166.435 -45.395 166.765 ;
        RECT -45.725 165.075 -45.395 165.405 ;
        RECT -45.725 163.715 -45.395 164.045 ;
        RECT -45.725 162.355 -45.395 162.685 ;
        RECT -45.725 160.995 -45.395 161.325 ;
        RECT -45.725 159.635 -45.395 159.965 ;
        RECT -45.725 158.275 -45.395 158.605 ;
        RECT -45.725 156.915 -45.395 157.245 ;
        RECT -45.725 155.555 -45.395 155.885 ;
        RECT -45.725 154.195 -45.395 154.525 ;
        RECT -45.725 152.835 -45.395 153.165 ;
        RECT -45.725 151.475 -45.395 151.805 ;
        RECT -45.725 150.115 -45.395 150.445 ;
        RECT -45.725 148.755 -45.395 149.085 ;
        RECT -45.725 147.395 -45.395 147.725 ;
        RECT -45.725 146.035 -45.395 146.365 ;
        RECT -45.725 144.675 -45.395 145.005 ;
        RECT -45.725 143.315 -45.395 143.645 ;
        RECT -45.725 141.955 -45.395 142.285 ;
        RECT -45.725 140.595 -45.395 140.925 ;
        RECT -45.725 139.235 -45.395 139.565 ;
        RECT -45.725 137.875 -45.395 138.205 ;
        RECT -45.725 136.515 -45.395 136.845 ;
        RECT -45.725 135.155 -45.395 135.485 ;
        RECT -45.725 133.795 -45.395 134.125 ;
        RECT -45.725 132.435 -45.395 132.765 ;
        RECT -45.725 131.075 -45.395 131.405 ;
        RECT -45.725 129.715 -45.395 130.045 ;
        RECT -45.725 128.355 -45.395 128.685 ;
        RECT -45.725 126.995 -45.395 127.325 ;
        RECT -45.725 125.635 -45.395 125.965 ;
        RECT -45.725 124.275 -45.395 124.605 ;
        RECT -45.725 122.915 -45.395 123.245 ;
        RECT -45.725 121.555 -45.395 121.885 ;
        RECT -45.725 120.195 -45.395 120.525 ;
        RECT -45.725 118.835 -45.395 119.165 ;
        RECT -45.725 117.475 -45.395 117.805 ;
        RECT -45.725 116.115 -45.395 116.445 ;
        RECT -45.725 114.755 -45.395 115.085 ;
        RECT -45.725 113.395 -45.395 113.725 ;
        RECT -45.725 112.035 -45.395 112.365 ;
        RECT -45.725 110.675 -45.395 111.005 ;
        RECT -45.725 109.315 -45.395 109.645 ;
        RECT -45.725 107.955 -45.395 108.285 ;
        RECT -45.725 106.595 -45.395 106.925 ;
        RECT -45.725 105.235 -45.395 105.565 ;
        RECT -45.725 103.875 -45.395 104.205 ;
        RECT -45.725 102.515 -45.395 102.845 ;
        RECT -45.725 101.155 -45.395 101.485 ;
        RECT -45.725 99.795 -45.395 100.125 ;
        RECT -45.725 98.435 -45.395 98.765 ;
        RECT -45.725 97.075 -45.395 97.405 ;
        RECT -45.725 95.715 -45.395 96.045 ;
        RECT -45.725 94.355 -45.395 94.685 ;
        RECT -45.725 92.995 -45.395 93.325 ;
        RECT -45.725 91.635 -45.395 91.965 ;
        RECT -45.725 90.275 -45.395 90.605 ;
        RECT -45.725 88.915 -45.395 89.245 ;
        RECT -45.725 87.555 -45.395 87.885 ;
        RECT -45.725 86.195 -45.395 86.525 ;
        RECT -45.725 84.835 -45.395 85.165 ;
        RECT -45.725 83.475 -45.395 83.805 ;
        RECT -45.725 82.115 -45.395 82.445 ;
        RECT -45.725 80.755 -45.395 81.085 ;
        RECT -45.725 79.395 -45.395 79.725 ;
        RECT -45.725 78.035 -45.395 78.365 ;
        RECT -45.725 76.675 -45.395 77.005 ;
        RECT -45.725 75.315 -45.395 75.645 ;
        RECT -45.725 73.955 -45.395 74.285 ;
        RECT -45.725 72.595 -45.395 72.925 ;
        RECT -45.725 71.235 -45.395 71.565 ;
        RECT -45.725 69.875 -45.395 70.205 ;
        RECT -45.725 68.515 -45.395 68.845 ;
        RECT -45.725 67.155 -45.395 67.485 ;
        RECT -45.725 65.795 -45.395 66.125 ;
        RECT -45.725 64.435 -45.395 64.765 ;
        RECT -45.725 63.075 -45.395 63.405 ;
        RECT -45.725 61.715 -45.395 62.045 ;
        RECT -45.725 60.355 -45.395 60.685 ;
        RECT -45.725 58.995 -45.395 59.325 ;
        RECT -45.725 57.635 -45.395 57.965 ;
        RECT -45.725 56.275 -45.395 56.605 ;
        RECT -45.725 54.915 -45.395 55.245 ;
        RECT -45.725 53.555 -45.395 53.885 ;
        RECT -45.725 52.195 -45.395 52.525 ;
        RECT -45.725 50.835 -45.395 51.165 ;
        RECT -45.725 49.475 -45.395 49.805 ;
        RECT -45.725 48.115 -45.395 48.445 ;
        RECT -45.725 46.755 -45.395 47.085 ;
        RECT -45.725 45.395 -45.395 45.725 ;
        RECT -45.725 44.035 -45.395 44.365 ;
        RECT -45.725 42.675 -45.395 43.005 ;
        RECT -45.725 41.315 -45.395 41.645 ;
        RECT -45.725 39.955 -45.395 40.285 ;
        RECT -45.725 38.595 -45.395 38.925 ;
        RECT -45.725 37.235 -45.395 37.565 ;
        RECT -45.725 35.875 -45.395 36.205 ;
        RECT -45.725 34.515 -45.395 34.845 ;
        RECT -45.725 33.155 -45.395 33.485 ;
        RECT -45.725 31.795 -45.395 32.125 ;
        RECT -45.725 30.435 -45.395 30.765 ;
        RECT -45.725 29.075 -45.395 29.405 ;
        RECT -45.725 27.715 -45.395 28.045 ;
        RECT -45.725 26.355 -45.395 26.685 ;
        RECT -45.725 24.995 -45.395 25.325 ;
        RECT -45.725 23.635 -45.395 23.965 ;
        RECT -45.725 22.275 -45.395 22.605 ;
        RECT -45.725 20.915 -45.395 21.245 ;
        RECT -45.725 19.555 -45.395 19.885 ;
        RECT -45.725 18.195 -45.395 18.525 ;
        RECT -45.725 16.835 -45.395 17.165 ;
        RECT -45.725 15.475 -45.395 15.805 ;
        RECT -45.725 14.115 -45.395 14.445 ;
        RECT -45.725 12.755 -45.395 13.085 ;
        RECT -45.725 11.395 -45.395 11.725 ;
        RECT -45.725 10.035 -45.395 10.365 ;
        RECT -45.725 8.675 -45.395 9.005 ;
        RECT -45.725 7.315 -45.395 7.645 ;
        RECT -45.725 5.955 -45.395 6.285 ;
        RECT -45.725 4.595 -45.395 4.925 ;
        RECT -45.725 3.235 -45.395 3.565 ;
        RECT -45.725 1.875 -45.395 2.205 ;
        RECT -45.725 0.515 -45.395 0.845 ;
        RECT -45.725 -0.845 -45.395 -0.515 ;
        RECT -45.725 -2.205 -45.395 -1.875 ;
        RECT -45.725 -4.925 -45.395 -4.595 ;
        RECT -45.725 -6.285 -45.395 -5.955 ;
        RECT -45.725 -7.645 -45.395 -7.315 ;
        RECT -45.725 -9.005 -45.395 -8.675 ;
        RECT -45.725 -10.365 -45.395 -10.035 ;
        RECT -45.725 -14.445 -45.395 -14.115 ;
        RECT -45.725 -15.805 -45.395 -15.475 ;
        RECT -45.725 -17.165 -45.395 -16.835 ;
        RECT -45.725 -18.525 -45.395 -18.195 ;
        RECT -45.725 -19.885 -45.395 -19.555 ;
        RECT -45.725 -21.245 -45.395 -20.915 ;
        RECT -45.725 -22.605 -45.395 -22.275 ;
        RECT -45.725 -23.965 -45.395 -23.635 ;
        RECT -45.725 -25.325 -45.395 -24.995 ;
        RECT -45.725 -32.125 -45.395 -31.795 ;
        RECT -45.725 -33.71 -45.395 -33.38 ;
        RECT -45.725 -34.845 -45.395 -34.515 ;
        RECT -45.725 -36.205 -45.395 -35.875 ;
        RECT -45.725 -38.925 -45.395 -38.595 ;
        RECT -45.725 -39.75 -45.395 -39.42 ;
        RECT -45.725 -41.645 -45.395 -41.315 ;
        RECT -45.725 -44.365 -45.395 -44.035 ;
        RECT -45.725 -49.805 -45.395 -49.475 ;
        RECT -45.725 -51.165 -45.395 -50.835 ;
        RECT -45.725 -53.885 -45.395 -53.555 ;
        RECT -45.725 -55.245 -45.395 -54.915 ;
        RECT -45.725 -59.325 -45.395 -58.995 ;
        RECT -45.725 -60.685 -45.395 -60.355 ;
        RECT -45.725 -67.485 -45.395 -67.155 ;
        RECT -45.725 -68.845 -45.395 -68.515 ;
        RECT -45.725 -70.205 -45.395 -69.875 ;
        RECT -45.725 -71.565 -45.395 -71.235 ;
        RECT -45.725 -72.925 -45.395 -72.595 ;
        RECT -45.725 -74.285 -45.395 -73.955 ;
        RECT -45.725 -75.645 -45.395 -75.315 ;
        RECT -45.725 -77.005 -45.395 -76.675 ;
        RECT -45.725 -78.365 -45.395 -78.035 ;
        RECT -45.725 -79.725 -45.395 -79.395 ;
        RECT -45.725 -81.085 -45.395 -80.755 ;
        RECT -45.725 -82.445 -45.395 -82.115 ;
        RECT -45.725 -83.805 -45.395 -83.475 ;
        RECT -45.725 -85.165 -45.395 -84.835 ;
        RECT -45.725 -86.525 -45.395 -86.195 ;
        RECT -45.725 -87.885 -45.395 -87.555 ;
        RECT -45.725 -89.245 -45.395 -88.915 ;
        RECT -45.725 -90.81 -45.395 -90.48 ;
        RECT -45.725 -91.965 -45.395 -91.635 ;
        RECT -45.725 -93.325 -45.395 -92.995 ;
        RECT -45.725 -94.685 -45.395 -94.355 ;
        RECT -45.725 -96.045 -45.395 -95.715 ;
        RECT -45.725 -97.405 -45.395 -97.075 ;
        RECT -45.725 -100.125 -45.395 -99.795 ;
        RECT -45.725 -101.35 -45.395 -101.02 ;
        RECT -45.725 -102.845 -45.395 -102.515 ;
        RECT -45.725 -104.205 -45.395 -103.875 ;
        RECT -45.725 -105.565 -45.395 -105.235 ;
        RECT -45.725 -108.285 -45.395 -107.955 ;
        RECT -45.725 -109.645 -45.395 -109.315 ;
        RECT -45.725 -115.085 -45.395 -114.755 ;
        RECT -45.725 -116.445 -45.395 -116.115 ;
        RECT -45.725 -117.805 -45.395 -117.475 ;
        RECT -45.725 -119.165 -45.395 -118.835 ;
        RECT -45.725 -120.525 -45.395 -120.195 ;
        RECT -45.725 -121.885 -45.395 -121.555 ;
        RECT -45.725 -123.245 -45.395 -122.915 ;
        RECT -45.725 -124.605 -45.395 -124.275 ;
        RECT -45.725 -125.965 -45.395 -125.635 ;
        RECT -45.725 -127.325 -45.395 -126.995 ;
        RECT -45.725 -128.685 -45.395 -128.355 ;
        RECT -45.725 -130.045 -45.395 -129.715 ;
        RECT -45.725 -131.405 -45.395 -131.075 ;
        RECT -45.725 -132.765 -45.395 -132.435 ;
        RECT -45.725 -134.125 -45.395 -133.795 ;
        RECT -45.725 -135.485 -45.395 -135.155 ;
        RECT -45.725 -136.845 -45.395 -136.515 ;
        RECT -45.725 -138.205 -45.395 -137.875 ;
        RECT -45.725 -139.565 -45.395 -139.235 ;
        RECT -45.725 -140.925 -45.395 -140.595 ;
        RECT -45.725 -142.285 -45.395 -141.955 ;
        RECT -45.725 -143.645 -45.395 -143.315 ;
        RECT -45.725 -145.005 -45.395 -144.675 ;
        RECT -45.725 -146.365 -45.395 -146.035 ;
        RECT -45.725 -147.725 -45.395 -147.395 ;
        RECT -45.725 -149.085 -45.395 -148.755 ;
        RECT -45.725 -150.445 -45.395 -150.115 ;
        RECT -45.725 -151.805 -45.395 -151.475 ;
        RECT -45.725 -153.165 -45.395 -152.835 ;
        RECT -45.725 -154.525 -45.395 -154.195 ;
        RECT -45.725 -155.885 -45.395 -155.555 ;
        RECT -45.725 -157.245 -45.395 -156.915 ;
        RECT -45.725 -158.605 -45.395 -158.275 ;
        RECT -45.725 -159.965 -45.395 -159.635 ;
        RECT -45.725 -161.325 -45.395 -160.995 ;
        RECT -45.725 -162.685 -45.395 -162.355 ;
        RECT -45.725 -164.045 -45.395 -163.715 ;
        RECT -45.725 -165.405 -45.395 -165.075 ;
        RECT -45.725 -166.765 -45.395 -166.435 ;
        RECT -45.725 -168.655 -45.395 -168.325 ;
        RECT -45.725 -169.485 -45.395 -169.155 ;
        RECT -45.725 -170.845 -45.395 -170.515 ;
        RECT -45.725 -173.565 -45.395 -173.235 ;
        RECT -45.725 -174.925 -45.395 -174.595 ;
        RECT -45.725 -177.645 -45.395 -177.315 ;
        RECT -45.725 -183.29 -45.395 -182.16 ;
        RECT -45.72 -183.405 -45.4 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -44.365 244.04 -44.035 245.17 ;
        RECT -44.365 239.875 -44.035 240.205 ;
        RECT -44.365 238.515 -44.035 238.845 ;
        RECT -44.365 237.155 -44.035 237.485 ;
        RECT -44.365 235.795 -44.035 236.125 ;
        RECT -44.365 234.435 -44.035 234.765 ;
        RECT -44.365 233.075 -44.035 233.405 ;
        RECT -44.365 231.715 -44.035 232.045 ;
        RECT -44.365 230.355 -44.035 230.685 ;
        RECT -44.365 228.995 -44.035 229.325 ;
        RECT -44.365 227.635 -44.035 227.965 ;
        RECT -44.365 226.275 -44.035 226.605 ;
        RECT -44.365 224.915 -44.035 225.245 ;
        RECT -44.365 223.555 -44.035 223.885 ;
        RECT -44.365 222.195 -44.035 222.525 ;
        RECT -44.365 220.835 -44.035 221.165 ;
        RECT -44.365 219.475 -44.035 219.805 ;
        RECT -44.365 218.115 -44.035 218.445 ;
        RECT -44.365 216.755 -44.035 217.085 ;
        RECT -44.365 215.395 -44.035 215.725 ;
        RECT -44.365 214.035 -44.035 214.365 ;
        RECT -44.365 212.675 -44.035 213.005 ;
        RECT -44.365 211.315 -44.035 211.645 ;
        RECT -44.365 209.955 -44.035 210.285 ;
        RECT -44.365 208.595 -44.035 208.925 ;
        RECT -44.365 207.235 -44.035 207.565 ;
        RECT -44.365 205.875 -44.035 206.205 ;
        RECT -44.365 204.515 -44.035 204.845 ;
        RECT -44.365 203.155 -44.035 203.485 ;
        RECT -44.365 201.795 -44.035 202.125 ;
        RECT -44.365 200.435 -44.035 200.765 ;
        RECT -44.365 199.075 -44.035 199.405 ;
        RECT -44.365 197.715 -44.035 198.045 ;
        RECT -44.365 196.355 -44.035 196.685 ;
        RECT -44.365 194.995 -44.035 195.325 ;
        RECT -44.365 193.635 -44.035 193.965 ;
        RECT -44.365 192.275 -44.035 192.605 ;
        RECT -44.365 190.915 -44.035 191.245 ;
        RECT -44.365 189.555 -44.035 189.885 ;
        RECT -44.365 188.195 -44.035 188.525 ;
        RECT -44.365 186.835 -44.035 187.165 ;
        RECT -44.365 185.475 -44.035 185.805 ;
        RECT -44.365 184.115 -44.035 184.445 ;
        RECT -44.365 182.755 -44.035 183.085 ;
        RECT -44.365 181.395 -44.035 181.725 ;
        RECT -44.365 180.035 -44.035 180.365 ;
        RECT -44.365 178.675 -44.035 179.005 ;
        RECT -44.365 177.315 -44.035 177.645 ;
        RECT -44.365 175.955 -44.035 176.285 ;
        RECT -44.365 174.595 -44.035 174.925 ;
        RECT -44.365 173.235 -44.035 173.565 ;
        RECT -44.365 171.875 -44.035 172.205 ;
        RECT -44.365 170.515 -44.035 170.845 ;
        RECT -44.365 169.155 -44.035 169.485 ;
        RECT -44.365 167.795 -44.035 168.125 ;
        RECT -44.365 166.435 -44.035 166.765 ;
        RECT -44.365 165.075 -44.035 165.405 ;
        RECT -44.365 163.715 -44.035 164.045 ;
        RECT -44.365 162.355 -44.035 162.685 ;
        RECT -44.365 160.995 -44.035 161.325 ;
        RECT -44.365 159.635 -44.035 159.965 ;
        RECT -44.365 158.275 -44.035 158.605 ;
        RECT -44.365 156.915 -44.035 157.245 ;
        RECT -44.365 155.555 -44.035 155.885 ;
        RECT -44.365 154.195 -44.035 154.525 ;
        RECT -44.365 152.835 -44.035 153.165 ;
        RECT -44.365 151.475 -44.035 151.805 ;
        RECT -44.365 150.115 -44.035 150.445 ;
        RECT -44.365 148.755 -44.035 149.085 ;
        RECT -44.365 147.395 -44.035 147.725 ;
        RECT -44.365 146.035 -44.035 146.365 ;
        RECT -44.365 144.675 -44.035 145.005 ;
        RECT -44.365 143.315 -44.035 143.645 ;
        RECT -44.365 141.955 -44.035 142.285 ;
        RECT -44.365 140.595 -44.035 140.925 ;
        RECT -44.365 139.235 -44.035 139.565 ;
        RECT -44.365 137.875 -44.035 138.205 ;
        RECT -44.365 136.515 -44.035 136.845 ;
        RECT -44.365 135.155 -44.035 135.485 ;
        RECT -44.365 133.795 -44.035 134.125 ;
        RECT -44.365 132.435 -44.035 132.765 ;
        RECT -44.365 131.075 -44.035 131.405 ;
        RECT -44.365 129.715 -44.035 130.045 ;
        RECT -44.365 128.355 -44.035 128.685 ;
        RECT -44.365 126.995 -44.035 127.325 ;
        RECT -44.365 125.635 -44.035 125.965 ;
        RECT -44.365 124.275 -44.035 124.605 ;
        RECT -44.365 122.915 -44.035 123.245 ;
        RECT -44.365 121.555 -44.035 121.885 ;
        RECT -44.365 120.195 -44.035 120.525 ;
        RECT -44.365 118.835 -44.035 119.165 ;
        RECT -44.365 117.475 -44.035 117.805 ;
        RECT -44.365 116.115 -44.035 116.445 ;
        RECT -44.365 114.755 -44.035 115.085 ;
        RECT -44.365 113.395 -44.035 113.725 ;
        RECT -44.365 112.035 -44.035 112.365 ;
        RECT -44.365 110.675 -44.035 111.005 ;
        RECT -44.365 109.315 -44.035 109.645 ;
        RECT -44.365 107.955 -44.035 108.285 ;
        RECT -44.365 106.595 -44.035 106.925 ;
        RECT -44.365 105.235 -44.035 105.565 ;
        RECT -44.365 103.875 -44.035 104.205 ;
        RECT -44.365 102.515 -44.035 102.845 ;
        RECT -44.365 101.155 -44.035 101.485 ;
        RECT -44.365 99.795 -44.035 100.125 ;
        RECT -44.365 98.435 -44.035 98.765 ;
        RECT -44.365 97.075 -44.035 97.405 ;
        RECT -44.365 95.715 -44.035 96.045 ;
        RECT -44.365 94.355 -44.035 94.685 ;
        RECT -44.365 92.995 -44.035 93.325 ;
        RECT -44.365 91.635 -44.035 91.965 ;
        RECT -44.365 90.275 -44.035 90.605 ;
        RECT -44.365 88.915 -44.035 89.245 ;
        RECT -44.365 87.555 -44.035 87.885 ;
        RECT -44.365 86.195 -44.035 86.525 ;
        RECT -44.365 84.835 -44.035 85.165 ;
        RECT -44.365 83.475 -44.035 83.805 ;
        RECT -44.365 82.115 -44.035 82.445 ;
        RECT -44.365 80.755 -44.035 81.085 ;
        RECT -44.365 79.395 -44.035 79.725 ;
        RECT -44.365 78.035 -44.035 78.365 ;
        RECT -44.365 76.675 -44.035 77.005 ;
        RECT -44.365 75.315 -44.035 75.645 ;
        RECT -44.365 73.955 -44.035 74.285 ;
        RECT -44.365 72.595 -44.035 72.925 ;
        RECT -44.365 71.235 -44.035 71.565 ;
        RECT -44.365 69.875 -44.035 70.205 ;
        RECT -44.365 68.515 -44.035 68.845 ;
        RECT -44.365 67.155 -44.035 67.485 ;
        RECT -44.365 65.795 -44.035 66.125 ;
        RECT -44.365 64.435 -44.035 64.765 ;
        RECT -44.365 63.075 -44.035 63.405 ;
        RECT -44.365 61.715 -44.035 62.045 ;
        RECT -44.365 60.355 -44.035 60.685 ;
        RECT -44.365 58.995 -44.035 59.325 ;
        RECT -44.365 57.635 -44.035 57.965 ;
        RECT -44.365 56.275 -44.035 56.605 ;
        RECT -44.365 54.915 -44.035 55.245 ;
        RECT -44.365 53.555 -44.035 53.885 ;
        RECT -44.365 52.195 -44.035 52.525 ;
        RECT -44.365 50.835 -44.035 51.165 ;
        RECT -44.365 49.475 -44.035 49.805 ;
        RECT -44.365 48.115 -44.035 48.445 ;
        RECT -44.365 46.755 -44.035 47.085 ;
        RECT -44.365 45.395 -44.035 45.725 ;
        RECT -44.365 44.035 -44.035 44.365 ;
        RECT -44.365 42.675 -44.035 43.005 ;
        RECT -44.365 41.315 -44.035 41.645 ;
        RECT -44.365 39.955 -44.035 40.285 ;
        RECT -44.365 38.595 -44.035 38.925 ;
        RECT -44.365 37.235 -44.035 37.565 ;
        RECT -44.365 35.875 -44.035 36.205 ;
        RECT -44.365 34.515 -44.035 34.845 ;
        RECT -44.365 33.155 -44.035 33.485 ;
        RECT -44.365 31.795 -44.035 32.125 ;
        RECT -44.365 30.435 -44.035 30.765 ;
        RECT -44.365 29.075 -44.035 29.405 ;
        RECT -44.365 27.715 -44.035 28.045 ;
        RECT -44.365 26.355 -44.035 26.685 ;
        RECT -44.365 24.995 -44.035 25.325 ;
        RECT -44.365 23.635 -44.035 23.965 ;
        RECT -44.365 22.275 -44.035 22.605 ;
        RECT -44.365 20.915 -44.035 21.245 ;
        RECT -44.365 19.555 -44.035 19.885 ;
        RECT -44.365 18.195 -44.035 18.525 ;
        RECT -44.365 16.835 -44.035 17.165 ;
        RECT -44.365 15.475 -44.035 15.805 ;
        RECT -44.365 14.115 -44.035 14.445 ;
        RECT -44.365 12.755 -44.035 13.085 ;
        RECT -44.365 11.395 -44.035 11.725 ;
        RECT -44.365 10.035 -44.035 10.365 ;
        RECT -44.365 8.675 -44.035 9.005 ;
        RECT -44.365 7.315 -44.035 7.645 ;
        RECT -44.365 5.955 -44.035 6.285 ;
        RECT -44.365 4.595 -44.035 4.925 ;
        RECT -44.365 3.235 -44.035 3.565 ;
        RECT -44.365 1.875 -44.035 2.205 ;
        RECT -44.365 0.515 -44.035 0.845 ;
        RECT -44.365 -0.845 -44.035 -0.515 ;
        RECT -44.365 -2.205 -44.035 -1.875 ;
        RECT -44.365 -4.925 -44.035 -4.595 ;
        RECT -44.365 -6.285 -44.035 -5.955 ;
        RECT -44.365 -7.645 -44.035 -7.315 ;
        RECT -44.365 -10.365 -44.035 -10.035 ;
        RECT -44.365 -14.445 -44.035 -14.115 ;
        RECT -44.365 -15.805 -44.035 -15.475 ;
        RECT -44.365 -17.165 -44.035 -16.835 ;
        RECT -44.365 -18.525 -44.035 -18.195 ;
        RECT -44.365 -19.885 -44.035 -19.555 ;
        RECT -44.365 -21.245 -44.035 -20.915 ;
        RECT -44.365 -22.605 -44.035 -22.275 ;
        RECT -44.365 -23.965 -44.035 -23.635 ;
        RECT -44.365 -25.325 -44.035 -24.995 ;
        RECT -44.365 -32.125 -44.035 -31.795 ;
        RECT -44.365 -33.71 -44.035 -33.38 ;
        RECT -44.365 -34.845 -44.035 -34.515 ;
        RECT -44.365 -36.205 -44.035 -35.875 ;
        RECT -44.365 -38.925 -44.035 -38.595 ;
        RECT -44.365 -39.75 -44.035 -39.42 ;
        RECT -44.365 -41.645 -44.035 -41.315 ;
        RECT -44.365 -44.365 -44.035 -44.035 ;
        RECT -44.365 -49.805 -44.035 -49.475 ;
        RECT -44.365 -51.165 -44.035 -50.835 ;
        RECT -44.365 -53.885 -44.035 -53.555 ;
        RECT -44.365 -55.245 -44.035 -54.915 ;
        RECT -44.365 -59.325 -44.035 -58.995 ;
        RECT -44.365 -60.685 -44.035 -60.355 ;
        RECT -44.36 -64.08 -44.04 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -44.365 -70.205 -44.035 -69.875 ;
        RECT -44.365 -71.565 -44.035 -71.235 ;
        RECT -44.365 -72.925 -44.035 -72.595 ;
        RECT -44.365 -74.285 -44.035 -73.955 ;
        RECT -44.365 -75.645 -44.035 -75.315 ;
        RECT -44.365 -77.005 -44.035 -76.675 ;
        RECT -44.365 -78.365 -44.035 -78.035 ;
        RECT -44.365 -79.725 -44.035 -79.395 ;
        RECT -44.365 -81.085 -44.035 -80.755 ;
        RECT -44.365 -82.445 -44.035 -82.115 ;
        RECT -44.365 -83.805 -44.035 -83.475 ;
        RECT -44.365 -85.165 -44.035 -84.835 ;
        RECT -44.365 -86.525 -44.035 -86.195 ;
        RECT -44.365 -87.885 -44.035 -87.555 ;
        RECT -44.365 -89.245 -44.035 -88.915 ;
        RECT -44.365 -90.81 -44.035 -90.48 ;
        RECT -44.365 -91.965 -44.035 -91.635 ;
        RECT -44.365 -93.325 -44.035 -92.995 ;
        RECT -44.365 -94.685 -44.035 -94.355 ;
        RECT -44.365 -96.045 -44.035 -95.715 ;
        RECT -44.365 -97.405 -44.035 -97.075 ;
        RECT -44.365 -100.125 -44.035 -99.795 ;
        RECT -44.365 -101.35 -44.035 -101.02 ;
        RECT -44.365 -102.845 -44.035 -102.515 ;
        RECT -44.365 -104.205 -44.035 -103.875 ;
        RECT -44.365 -105.565 -44.035 -105.235 ;
        RECT -44.365 -108.285 -44.035 -107.955 ;
        RECT -44.365 -109.645 -44.035 -109.315 ;
        RECT -44.365 -115.085 -44.035 -114.755 ;
        RECT -44.365 -116.445 -44.035 -116.115 ;
        RECT -44.365 -117.805 -44.035 -117.475 ;
        RECT -44.365 -119.165 -44.035 -118.835 ;
        RECT -44.365 -120.525 -44.035 -120.195 ;
        RECT -44.365 -121.885 -44.035 -121.555 ;
        RECT -44.365 -123.245 -44.035 -122.915 ;
        RECT -44.365 -124.605 -44.035 -124.275 ;
        RECT -44.365 -125.965 -44.035 -125.635 ;
        RECT -44.365 -127.325 -44.035 -126.995 ;
        RECT -44.365 -128.685 -44.035 -128.355 ;
        RECT -44.365 -130.045 -44.035 -129.715 ;
        RECT -44.365 -131.405 -44.035 -131.075 ;
        RECT -44.365 -132.765 -44.035 -132.435 ;
        RECT -44.365 -134.125 -44.035 -133.795 ;
        RECT -44.365 -135.485 -44.035 -135.155 ;
        RECT -44.365 -136.845 -44.035 -136.515 ;
        RECT -44.365 -138.205 -44.035 -137.875 ;
        RECT -44.365 -139.565 -44.035 -139.235 ;
        RECT -44.365 -140.925 -44.035 -140.595 ;
        RECT -44.365 -142.285 -44.035 -141.955 ;
        RECT -44.365 -143.645 -44.035 -143.315 ;
        RECT -44.365 -145.005 -44.035 -144.675 ;
        RECT -44.365 -146.365 -44.035 -146.035 ;
        RECT -44.365 -147.725 -44.035 -147.395 ;
        RECT -44.365 -149.085 -44.035 -148.755 ;
        RECT -44.365 -150.445 -44.035 -150.115 ;
        RECT -44.365 -151.805 -44.035 -151.475 ;
        RECT -44.365 -153.165 -44.035 -152.835 ;
        RECT -44.365 -154.525 -44.035 -154.195 ;
        RECT -44.365 -155.885 -44.035 -155.555 ;
        RECT -44.365 -157.245 -44.035 -156.915 ;
        RECT -44.365 -158.605 -44.035 -158.275 ;
        RECT -44.365 -159.965 -44.035 -159.635 ;
        RECT -44.365 -161.325 -44.035 -160.995 ;
        RECT -44.365 -162.685 -44.035 -162.355 ;
        RECT -44.365 -164.045 -44.035 -163.715 ;
        RECT -44.365 -165.405 -44.035 -165.075 ;
        RECT -44.365 -166.765 -44.035 -166.435 ;
        RECT -44.365 -168.655 -44.035 -168.325 ;
        RECT -44.365 -169.485 -44.035 -169.155 ;
        RECT -44.365 -170.845 -44.035 -170.515 ;
        RECT -44.365 -172.205 -44.035 -171.875 ;
        RECT -44.365 -173.565 -44.035 -173.235 ;
        RECT -44.365 -174.925 -44.035 -174.595 ;
        RECT -44.365 -177.645 -44.035 -177.315 ;
        RECT -44.365 -183.29 -44.035 -182.16 ;
        RECT -44.36 -183.405 -44.04 -68.52 ;
    END
    PORT
      LAYER met3 ;
        RECT -43.005 244.04 -42.675 245.17 ;
        RECT -43.005 239.875 -42.675 240.205 ;
        RECT -43.005 238.515 -42.675 238.845 ;
        RECT -43.005 237.155 -42.675 237.485 ;
        RECT -43.005 235.795 -42.675 236.125 ;
        RECT -43.005 234.435 -42.675 234.765 ;
        RECT -43.005 233.075 -42.675 233.405 ;
        RECT -43.005 231.715 -42.675 232.045 ;
        RECT -43.005 230.355 -42.675 230.685 ;
        RECT -43.005 228.995 -42.675 229.325 ;
        RECT -43.005 227.635 -42.675 227.965 ;
        RECT -43.005 226.275 -42.675 226.605 ;
        RECT -43.005 224.915 -42.675 225.245 ;
        RECT -43.005 223.555 -42.675 223.885 ;
        RECT -43.005 222.195 -42.675 222.525 ;
        RECT -43.005 220.835 -42.675 221.165 ;
        RECT -43.005 219.475 -42.675 219.805 ;
        RECT -43.005 218.115 -42.675 218.445 ;
        RECT -43.005 216.755 -42.675 217.085 ;
        RECT -43.005 215.395 -42.675 215.725 ;
        RECT -43.005 214.035 -42.675 214.365 ;
        RECT -43.005 212.675 -42.675 213.005 ;
        RECT -43.005 211.315 -42.675 211.645 ;
        RECT -43.005 209.955 -42.675 210.285 ;
        RECT -43.005 208.595 -42.675 208.925 ;
        RECT -43.005 207.235 -42.675 207.565 ;
        RECT -43.005 205.875 -42.675 206.205 ;
        RECT -43.005 204.515 -42.675 204.845 ;
        RECT -43.005 203.155 -42.675 203.485 ;
        RECT -43.005 201.795 -42.675 202.125 ;
        RECT -43.005 200.435 -42.675 200.765 ;
        RECT -43.005 199.075 -42.675 199.405 ;
        RECT -43.005 197.715 -42.675 198.045 ;
        RECT -43.005 196.355 -42.675 196.685 ;
        RECT -43.005 194.995 -42.675 195.325 ;
        RECT -43.005 193.635 -42.675 193.965 ;
        RECT -43.005 192.275 -42.675 192.605 ;
        RECT -43.005 190.915 -42.675 191.245 ;
        RECT -43.005 189.555 -42.675 189.885 ;
        RECT -43.005 188.195 -42.675 188.525 ;
        RECT -43.005 186.835 -42.675 187.165 ;
        RECT -43.005 185.475 -42.675 185.805 ;
        RECT -43.005 184.115 -42.675 184.445 ;
        RECT -43.005 182.755 -42.675 183.085 ;
        RECT -43.005 181.395 -42.675 181.725 ;
        RECT -43.005 180.035 -42.675 180.365 ;
        RECT -43.005 178.675 -42.675 179.005 ;
        RECT -43.005 177.315 -42.675 177.645 ;
        RECT -43.005 175.955 -42.675 176.285 ;
        RECT -43.005 174.595 -42.675 174.925 ;
        RECT -43.005 173.235 -42.675 173.565 ;
        RECT -43.005 171.875 -42.675 172.205 ;
        RECT -43.005 170.515 -42.675 170.845 ;
        RECT -43.005 169.155 -42.675 169.485 ;
        RECT -43.005 167.795 -42.675 168.125 ;
        RECT -43.005 166.435 -42.675 166.765 ;
        RECT -43.005 165.075 -42.675 165.405 ;
        RECT -43.005 163.715 -42.675 164.045 ;
        RECT -43.005 162.355 -42.675 162.685 ;
        RECT -43.005 160.995 -42.675 161.325 ;
        RECT -43.005 159.635 -42.675 159.965 ;
        RECT -43.005 158.275 -42.675 158.605 ;
        RECT -43.005 156.915 -42.675 157.245 ;
        RECT -43.005 155.555 -42.675 155.885 ;
        RECT -43.005 154.195 -42.675 154.525 ;
        RECT -43.005 152.835 -42.675 153.165 ;
        RECT -43.005 151.475 -42.675 151.805 ;
        RECT -43.005 150.115 -42.675 150.445 ;
        RECT -43.005 148.755 -42.675 149.085 ;
        RECT -43.005 147.395 -42.675 147.725 ;
        RECT -43.005 146.035 -42.675 146.365 ;
        RECT -43.005 144.675 -42.675 145.005 ;
        RECT -43.005 143.315 -42.675 143.645 ;
        RECT -43.005 141.955 -42.675 142.285 ;
        RECT -43.005 140.595 -42.675 140.925 ;
        RECT -43.005 139.235 -42.675 139.565 ;
        RECT -43.005 137.875 -42.675 138.205 ;
        RECT -43.005 136.515 -42.675 136.845 ;
        RECT -43.005 135.155 -42.675 135.485 ;
        RECT -43.005 133.795 -42.675 134.125 ;
        RECT -43.005 132.435 -42.675 132.765 ;
        RECT -43.005 131.075 -42.675 131.405 ;
        RECT -43.005 129.715 -42.675 130.045 ;
        RECT -43.005 128.355 -42.675 128.685 ;
        RECT -43.005 126.995 -42.675 127.325 ;
        RECT -43.005 125.635 -42.675 125.965 ;
        RECT -43.005 124.275 -42.675 124.605 ;
        RECT -43.005 122.915 -42.675 123.245 ;
        RECT -43.005 121.555 -42.675 121.885 ;
        RECT -43.005 120.195 -42.675 120.525 ;
        RECT -43.005 118.835 -42.675 119.165 ;
        RECT -43.005 117.475 -42.675 117.805 ;
        RECT -43.005 116.115 -42.675 116.445 ;
        RECT -43.005 114.755 -42.675 115.085 ;
        RECT -43.005 113.395 -42.675 113.725 ;
        RECT -43.005 112.035 -42.675 112.365 ;
        RECT -43.005 110.675 -42.675 111.005 ;
        RECT -43.005 109.315 -42.675 109.645 ;
        RECT -43.005 107.955 -42.675 108.285 ;
        RECT -43.005 106.595 -42.675 106.925 ;
        RECT -43.005 105.235 -42.675 105.565 ;
        RECT -43.005 103.875 -42.675 104.205 ;
        RECT -43.005 102.515 -42.675 102.845 ;
        RECT -43.005 101.155 -42.675 101.485 ;
        RECT -43.005 99.795 -42.675 100.125 ;
        RECT -43.005 98.435 -42.675 98.765 ;
        RECT -43.005 97.075 -42.675 97.405 ;
        RECT -43.005 95.715 -42.675 96.045 ;
        RECT -43.005 94.355 -42.675 94.685 ;
        RECT -43.005 92.995 -42.675 93.325 ;
        RECT -43.005 91.635 -42.675 91.965 ;
        RECT -43.005 90.275 -42.675 90.605 ;
        RECT -43.005 88.915 -42.675 89.245 ;
        RECT -43.005 87.555 -42.675 87.885 ;
        RECT -43.005 86.195 -42.675 86.525 ;
        RECT -43.005 84.835 -42.675 85.165 ;
        RECT -43.005 83.475 -42.675 83.805 ;
        RECT -43.005 82.115 -42.675 82.445 ;
        RECT -43.005 80.755 -42.675 81.085 ;
        RECT -43.005 79.395 -42.675 79.725 ;
        RECT -43.005 78.035 -42.675 78.365 ;
        RECT -43.005 76.675 -42.675 77.005 ;
        RECT -43.005 75.315 -42.675 75.645 ;
        RECT -43.005 73.955 -42.675 74.285 ;
        RECT -43.005 72.595 -42.675 72.925 ;
        RECT -43.005 71.235 -42.675 71.565 ;
        RECT -43.005 69.875 -42.675 70.205 ;
        RECT -43.005 68.515 -42.675 68.845 ;
        RECT -43.005 67.155 -42.675 67.485 ;
        RECT -43.005 65.795 -42.675 66.125 ;
        RECT -43.005 64.435 -42.675 64.765 ;
        RECT -43.005 63.075 -42.675 63.405 ;
        RECT -43.005 61.715 -42.675 62.045 ;
        RECT -43.005 60.355 -42.675 60.685 ;
        RECT -43.005 58.995 -42.675 59.325 ;
        RECT -43.005 57.635 -42.675 57.965 ;
        RECT -43.005 56.275 -42.675 56.605 ;
        RECT -43.005 54.915 -42.675 55.245 ;
        RECT -43.005 53.555 -42.675 53.885 ;
        RECT -43.005 52.195 -42.675 52.525 ;
        RECT -43.005 50.835 -42.675 51.165 ;
        RECT -43.005 49.475 -42.675 49.805 ;
        RECT -43.005 48.115 -42.675 48.445 ;
        RECT -43.005 46.755 -42.675 47.085 ;
        RECT -43.005 45.395 -42.675 45.725 ;
        RECT -43.005 44.035 -42.675 44.365 ;
        RECT -43.005 42.675 -42.675 43.005 ;
        RECT -43.005 41.315 -42.675 41.645 ;
        RECT -43.005 39.955 -42.675 40.285 ;
        RECT -43.005 38.595 -42.675 38.925 ;
        RECT -43.005 37.235 -42.675 37.565 ;
        RECT -43.005 35.875 -42.675 36.205 ;
        RECT -43.005 34.515 -42.675 34.845 ;
        RECT -43.005 33.155 -42.675 33.485 ;
        RECT -43.005 31.795 -42.675 32.125 ;
        RECT -43.005 30.435 -42.675 30.765 ;
        RECT -43.005 29.075 -42.675 29.405 ;
        RECT -43.005 27.715 -42.675 28.045 ;
        RECT -43.005 26.355 -42.675 26.685 ;
        RECT -43.005 24.995 -42.675 25.325 ;
        RECT -43.005 23.635 -42.675 23.965 ;
        RECT -43.005 22.275 -42.675 22.605 ;
        RECT -43.005 20.915 -42.675 21.245 ;
        RECT -43.005 19.555 -42.675 19.885 ;
        RECT -43.005 18.195 -42.675 18.525 ;
        RECT -43.005 16.835 -42.675 17.165 ;
        RECT -43.005 15.475 -42.675 15.805 ;
        RECT -43.005 14.115 -42.675 14.445 ;
        RECT -43.005 12.755 -42.675 13.085 ;
        RECT -43.005 11.395 -42.675 11.725 ;
        RECT -43.005 10.035 -42.675 10.365 ;
        RECT -43.005 8.675 -42.675 9.005 ;
        RECT -43.005 7.315 -42.675 7.645 ;
        RECT -43.005 5.955 -42.675 6.285 ;
        RECT -43.005 4.595 -42.675 4.925 ;
        RECT -43.005 3.235 -42.675 3.565 ;
        RECT -43.005 1.875 -42.675 2.205 ;
        RECT -43.005 0.515 -42.675 0.845 ;
        RECT -43.005 -0.845 -42.675 -0.515 ;
        RECT -43.005 -2.205 -42.675 -1.875 ;
        RECT -43.005 -4.925 -42.675 -4.595 ;
        RECT -43.005 -6.285 -42.675 -5.955 ;
        RECT -43.005 -10.365 -42.675 -10.035 ;
        RECT -43.005 -14.445 -42.675 -14.115 ;
        RECT -43.005 -15.805 -42.675 -15.475 ;
        RECT -43.005 -17.165 -42.675 -16.835 ;
        RECT -43.005 -18.525 -42.675 -18.195 ;
        RECT -43.005 -19.885 -42.675 -19.555 ;
        RECT -43.005 -21.245 -42.675 -20.915 ;
        RECT -43.005 -22.605 -42.675 -22.275 ;
        RECT -43.005 -23.965 -42.675 -23.635 ;
        RECT -43.005 -25.325 -42.675 -24.995 ;
        RECT -43.005 -32.125 -42.675 -31.795 ;
        RECT -43.005 -33.71 -42.675 -33.38 ;
        RECT -43.005 -34.845 -42.675 -34.515 ;
        RECT -43.005 -36.205 -42.675 -35.875 ;
        RECT -43.005 -38.925 -42.675 -38.595 ;
        RECT -43.005 -39.75 -42.675 -39.42 ;
        RECT -43.005 -41.645 -42.675 -41.315 ;
        RECT -43.005 -44.365 -42.675 -44.035 ;
        RECT -43.005 -49.805 -42.675 -49.475 ;
        RECT -43.005 -51.165 -42.675 -50.835 ;
        RECT -43.005 -53.885 -42.675 -53.555 ;
        RECT -43.005 -55.245 -42.675 -54.915 ;
        RECT -43.005 -59.325 -42.675 -58.995 ;
        RECT -43.005 -60.685 -42.675 -60.355 ;
        RECT -43 -63.4 -42.68 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -43.005 -67.485 -42.675 -67.155 ;
        RECT -43.005 -70.205 -42.675 -69.875 ;
        RECT -43.005 -71.565 -42.675 -71.235 ;
        RECT -43.005 -72.925 -42.675 -72.595 ;
        RECT -43.005 -74.285 -42.675 -73.955 ;
        RECT -43.005 -75.645 -42.675 -75.315 ;
        RECT -43.005 -77.005 -42.675 -76.675 ;
        RECT -43.005 -78.365 -42.675 -78.035 ;
        RECT -43.005 -79.725 -42.675 -79.395 ;
        RECT -43.005 -81.085 -42.675 -80.755 ;
        RECT -43.005 -82.445 -42.675 -82.115 ;
        RECT -43.005 -83.805 -42.675 -83.475 ;
        RECT -43.005 -85.165 -42.675 -84.835 ;
        RECT -43.005 -86.525 -42.675 -86.195 ;
        RECT -43.005 -87.885 -42.675 -87.555 ;
        RECT -43.005 -89.245 -42.675 -88.915 ;
        RECT -43.005 -90.81 -42.675 -90.48 ;
        RECT -43.005 -91.965 -42.675 -91.635 ;
        RECT -43.005 -93.325 -42.675 -92.995 ;
        RECT -43.005 -94.685 -42.675 -94.355 ;
        RECT -43.005 -96.045 -42.675 -95.715 ;
        RECT -43.005 -97.405 -42.675 -97.075 ;
        RECT -43.005 -100.125 -42.675 -99.795 ;
        RECT -43.005 -101.35 -42.675 -101.02 ;
        RECT -43.005 -102.845 -42.675 -102.515 ;
        RECT -43.005 -104.205 -42.675 -103.875 ;
        RECT -43.005 -105.565 -42.675 -105.235 ;
        RECT -43.005 -108.285 -42.675 -107.955 ;
        RECT -43.005 -109.645 -42.675 -109.315 ;
        RECT -43.005 -112.365 -42.675 -112.035 ;
        RECT -43.005 -113.725 -42.675 -113.395 ;
        RECT -43.005 -115.085 -42.675 -114.755 ;
        RECT -43.005 -116.445 -42.675 -116.115 ;
        RECT -43.005 -117.805 -42.675 -117.475 ;
        RECT -43.005 -119.165 -42.675 -118.835 ;
        RECT -43.005 -120.525 -42.675 -120.195 ;
        RECT -43.005 -121.885 -42.675 -121.555 ;
        RECT -43.005 -123.245 -42.675 -122.915 ;
        RECT -43.005 -124.605 -42.675 -124.275 ;
        RECT -43.005 -125.965 -42.675 -125.635 ;
        RECT -43.005 -127.325 -42.675 -126.995 ;
        RECT -43.005 -128.685 -42.675 -128.355 ;
        RECT -43.005 -130.045 -42.675 -129.715 ;
        RECT -43.005 -131.405 -42.675 -131.075 ;
        RECT -43.005 -132.765 -42.675 -132.435 ;
        RECT -43.005 -134.125 -42.675 -133.795 ;
        RECT -43.005 -135.485 -42.675 -135.155 ;
        RECT -43.005 -136.845 -42.675 -136.515 ;
        RECT -43.005 -138.205 -42.675 -137.875 ;
        RECT -43.005 -139.565 -42.675 -139.235 ;
        RECT -43.005 -140.925 -42.675 -140.595 ;
        RECT -43.005 -142.285 -42.675 -141.955 ;
        RECT -43.005 -143.645 -42.675 -143.315 ;
        RECT -43.005 -145.005 -42.675 -144.675 ;
        RECT -43.005 -146.365 -42.675 -146.035 ;
        RECT -43.005 -147.725 -42.675 -147.395 ;
        RECT -43.005 -149.085 -42.675 -148.755 ;
        RECT -43.005 -150.445 -42.675 -150.115 ;
        RECT -43.005 -151.805 -42.675 -151.475 ;
        RECT -43.005 -153.165 -42.675 -152.835 ;
        RECT -43.005 -154.525 -42.675 -154.195 ;
        RECT -43.005 -155.885 -42.675 -155.555 ;
        RECT -43.005 -157.245 -42.675 -156.915 ;
        RECT -43.005 -158.605 -42.675 -158.275 ;
        RECT -43.005 -159.965 -42.675 -159.635 ;
        RECT -43.005 -161.325 -42.675 -160.995 ;
        RECT -43.005 -162.685 -42.675 -162.355 ;
        RECT -43.005 -164.045 -42.675 -163.715 ;
        RECT -43.005 -165.405 -42.675 -165.075 ;
        RECT -43.005 -166.765 -42.675 -166.435 ;
        RECT -43.005 -168.655 -42.675 -168.325 ;
        RECT -43.005 -169.485 -42.675 -169.155 ;
        RECT -43.005 -170.845 -42.675 -170.515 ;
        RECT -43.005 -172.205 -42.675 -171.875 ;
        RECT -43.005 -173.565 -42.675 -173.235 ;
        RECT -43.005 -174.925 -42.675 -174.595 ;
        RECT -43.005 -177.645 -42.675 -177.315 ;
        RECT -43.005 -183.29 -42.675 -182.16 ;
        RECT -43 -183.405 -42.68 -67.155 ;
    END
    PORT
      LAYER met3 ;
        RECT -41.645 101.155 -41.315 101.485 ;
        RECT -41.645 99.795 -41.315 100.125 ;
        RECT -41.645 98.435 -41.315 98.765 ;
        RECT -41.645 97.075 -41.315 97.405 ;
        RECT -41.645 95.715 -41.315 96.045 ;
        RECT -41.645 94.355 -41.315 94.685 ;
        RECT -41.645 92.995 -41.315 93.325 ;
        RECT -41.645 91.635 -41.315 91.965 ;
        RECT -41.645 90.275 -41.315 90.605 ;
        RECT -41.645 88.915 -41.315 89.245 ;
        RECT -41.645 87.555 -41.315 87.885 ;
        RECT -41.645 86.195 -41.315 86.525 ;
        RECT -41.645 84.835 -41.315 85.165 ;
        RECT -41.645 83.475 -41.315 83.805 ;
        RECT -41.645 82.115 -41.315 82.445 ;
        RECT -41.645 80.755 -41.315 81.085 ;
        RECT -41.645 79.395 -41.315 79.725 ;
        RECT -41.645 78.035 -41.315 78.365 ;
        RECT -41.645 76.675 -41.315 77.005 ;
        RECT -41.645 75.315 -41.315 75.645 ;
        RECT -41.645 73.955 -41.315 74.285 ;
        RECT -41.645 72.595 -41.315 72.925 ;
        RECT -41.645 71.235 -41.315 71.565 ;
        RECT -41.645 69.875 -41.315 70.205 ;
        RECT -41.645 68.515 -41.315 68.845 ;
        RECT -41.645 67.155 -41.315 67.485 ;
        RECT -41.645 65.795 -41.315 66.125 ;
        RECT -41.645 64.435 -41.315 64.765 ;
        RECT -41.645 63.075 -41.315 63.405 ;
        RECT -41.645 61.715 -41.315 62.045 ;
        RECT -41.645 60.355 -41.315 60.685 ;
        RECT -41.645 58.995 -41.315 59.325 ;
        RECT -41.645 57.635 -41.315 57.965 ;
        RECT -41.645 56.275 -41.315 56.605 ;
        RECT -41.645 54.915 -41.315 55.245 ;
        RECT -41.645 53.555 -41.315 53.885 ;
        RECT -41.645 52.195 -41.315 52.525 ;
        RECT -41.645 50.835 -41.315 51.165 ;
        RECT -41.645 49.475 -41.315 49.805 ;
        RECT -41.645 48.115 -41.315 48.445 ;
        RECT -41.645 46.755 -41.315 47.085 ;
        RECT -41.645 45.395 -41.315 45.725 ;
        RECT -41.645 44.035 -41.315 44.365 ;
        RECT -41.645 42.675 -41.315 43.005 ;
        RECT -41.645 41.315 -41.315 41.645 ;
        RECT -41.645 39.955 -41.315 40.285 ;
        RECT -41.645 38.595 -41.315 38.925 ;
        RECT -41.645 37.235 -41.315 37.565 ;
        RECT -41.645 35.875 -41.315 36.205 ;
        RECT -41.645 34.515 -41.315 34.845 ;
        RECT -41.645 33.155 -41.315 33.485 ;
        RECT -41.645 31.795 -41.315 32.125 ;
        RECT -41.645 30.435 -41.315 30.765 ;
        RECT -41.645 29.075 -41.315 29.405 ;
        RECT -41.645 27.715 -41.315 28.045 ;
        RECT -41.645 26.355 -41.315 26.685 ;
        RECT -41.645 24.995 -41.315 25.325 ;
        RECT -41.645 23.635 -41.315 23.965 ;
        RECT -41.645 22.275 -41.315 22.605 ;
        RECT -41.645 20.915 -41.315 21.245 ;
        RECT -41.645 19.555 -41.315 19.885 ;
        RECT -41.645 18.195 -41.315 18.525 ;
        RECT -41.645 16.835 -41.315 17.165 ;
        RECT -41.645 15.475 -41.315 15.805 ;
        RECT -41.645 14.115 -41.315 14.445 ;
        RECT -41.645 12.755 -41.315 13.085 ;
        RECT -41.645 11.395 -41.315 11.725 ;
        RECT -41.645 10.035 -41.315 10.365 ;
        RECT -41.645 8.675 -41.315 9.005 ;
        RECT -41.645 7.315 -41.315 7.645 ;
        RECT -41.645 5.955 -41.315 6.285 ;
        RECT -41.645 4.595 -41.315 4.925 ;
        RECT -41.645 3.235 -41.315 3.565 ;
        RECT -41.645 1.875 -41.315 2.205 ;
        RECT -41.645 0.515 -41.315 0.845 ;
        RECT -41.645 -0.845 -41.315 -0.515 ;
        RECT -41.645 -2.205 -41.315 -1.875 ;
        RECT -41.645 -4.925 -41.315 -4.595 ;
        RECT -41.645 -6.285 -41.315 -5.955 ;
        RECT -41.645 -10.365 -41.315 -10.035 ;
        RECT -41.645 -14.445 -41.315 -14.115 ;
        RECT -41.645 -15.805 -41.315 -15.475 ;
        RECT -41.645 -17.165 -41.315 -16.835 ;
        RECT -41.645 -18.525 -41.315 -18.195 ;
        RECT -41.645 -19.885 -41.315 -19.555 ;
        RECT -41.645 -21.245 -41.315 -20.915 ;
        RECT -41.645 -22.605 -41.315 -22.275 ;
        RECT -41.645 -23.965 -41.315 -23.635 ;
        RECT -41.645 -25.325 -41.315 -24.995 ;
        RECT -41.645 -32.125 -41.315 -31.795 ;
        RECT -41.645 -33.71 -41.315 -33.38 ;
        RECT -41.645 -34.845 -41.315 -34.515 ;
        RECT -41.645 -36.205 -41.315 -35.875 ;
        RECT -41.645 -38.925 -41.315 -38.595 ;
        RECT -41.645 -39.75 -41.315 -39.42 ;
        RECT -41.645 -41.645 -41.315 -41.315 ;
        RECT -41.645 -44.365 -41.315 -44.035 ;
        RECT -41.645 -49.805 -41.315 -49.475 ;
        RECT -41.645 -51.165 -41.315 -50.835 ;
        RECT -41.645 -53.885 -41.315 -53.555 ;
        RECT -41.645 -55.245 -41.315 -54.915 ;
        RECT -41.645 -59.325 -41.315 -58.995 ;
        RECT -41.645 -60.685 -41.315 -60.355 ;
        RECT -41.645 -67.485 -41.315 -67.155 ;
        RECT -41.645 -70.205 -41.315 -69.875 ;
        RECT -41.645 -71.565 -41.315 -71.235 ;
        RECT -41.645 -72.925 -41.315 -72.595 ;
        RECT -41.645 -74.285 -41.315 -73.955 ;
        RECT -41.645 -75.645 -41.315 -75.315 ;
        RECT -41.645 -77.005 -41.315 -76.675 ;
        RECT -41.645 -78.365 -41.315 -78.035 ;
        RECT -41.645 -79.725 -41.315 -79.395 ;
        RECT -41.645 -81.085 -41.315 -80.755 ;
        RECT -41.645 -82.445 -41.315 -82.115 ;
        RECT -41.645 -83.805 -41.315 -83.475 ;
        RECT -41.645 -85.165 -41.315 -84.835 ;
        RECT -41.645 -86.525 -41.315 -86.195 ;
        RECT -41.645 -87.885 -41.315 -87.555 ;
        RECT -41.645 -89.245 -41.315 -88.915 ;
        RECT -41.645 -90.81 -41.315 -90.48 ;
        RECT -41.645 -91.965 -41.315 -91.635 ;
        RECT -41.645 -93.325 -41.315 -92.995 ;
        RECT -41.645 -94.685 -41.315 -94.355 ;
        RECT -41.645 -96.045 -41.315 -95.715 ;
        RECT -41.645 -97.405 -41.315 -97.075 ;
        RECT -41.645 -100.125 -41.315 -99.795 ;
        RECT -41.645 -101.35 -41.315 -101.02 ;
        RECT -41.645 -102.845 -41.315 -102.515 ;
        RECT -41.645 -104.205 -41.315 -103.875 ;
        RECT -41.645 -105.565 -41.315 -105.235 ;
        RECT -41.645 -108.285 -41.315 -107.955 ;
        RECT -41.645 -109.645 -41.315 -109.315 ;
        RECT -41.64 -111.68 -41.32 245.285 ;
        RECT -41.645 244.04 -41.315 245.17 ;
        RECT -41.645 239.875 -41.315 240.205 ;
        RECT -41.645 238.515 -41.315 238.845 ;
        RECT -41.645 237.155 -41.315 237.485 ;
        RECT -41.645 235.795 -41.315 236.125 ;
        RECT -41.645 234.435 -41.315 234.765 ;
        RECT -41.645 233.075 -41.315 233.405 ;
        RECT -41.645 231.715 -41.315 232.045 ;
        RECT -41.645 230.355 -41.315 230.685 ;
        RECT -41.645 228.995 -41.315 229.325 ;
        RECT -41.645 227.635 -41.315 227.965 ;
        RECT -41.645 226.275 -41.315 226.605 ;
        RECT -41.645 224.915 -41.315 225.245 ;
        RECT -41.645 223.555 -41.315 223.885 ;
        RECT -41.645 222.195 -41.315 222.525 ;
        RECT -41.645 220.835 -41.315 221.165 ;
        RECT -41.645 219.475 -41.315 219.805 ;
        RECT -41.645 218.115 -41.315 218.445 ;
        RECT -41.645 216.755 -41.315 217.085 ;
        RECT -41.645 215.395 -41.315 215.725 ;
        RECT -41.645 214.035 -41.315 214.365 ;
        RECT -41.645 212.675 -41.315 213.005 ;
        RECT -41.645 211.315 -41.315 211.645 ;
        RECT -41.645 209.955 -41.315 210.285 ;
        RECT -41.645 208.595 -41.315 208.925 ;
        RECT -41.645 207.235 -41.315 207.565 ;
        RECT -41.645 205.875 -41.315 206.205 ;
        RECT -41.645 204.515 -41.315 204.845 ;
        RECT -41.645 203.155 -41.315 203.485 ;
        RECT -41.645 201.795 -41.315 202.125 ;
        RECT -41.645 200.435 -41.315 200.765 ;
        RECT -41.645 199.075 -41.315 199.405 ;
        RECT -41.645 197.715 -41.315 198.045 ;
        RECT -41.645 196.355 -41.315 196.685 ;
        RECT -41.645 194.995 -41.315 195.325 ;
        RECT -41.645 193.635 -41.315 193.965 ;
        RECT -41.645 192.275 -41.315 192.605 ;
        RECT -41.645 190.915 -41.315 191.245 ;
        RECT -41.645 189.555 -41.315 189.885 ;
        RECT -41.645 188.195 -41.315 188.525 ;
        RECT -41.645 186.835 -41.315 187.165 ;
        RECT -41.645 185.475 -41.315 185.805 ;
        RECT -41.645 184.115 -41.315 184.445 ;
        RECT -41.645 182.755 -41.315 183.085 ;
        RECT -41.645 181.395 -41.315 181.725 ;
        RECT -41.645 180.035 -41.315 180.365 ;
        RECT -41.645 178.675 -41.315 179.005 ;
        RECT -41.645 177.315 -41.315 177.645 ;
        RECT -41.645 175.955 -41.315 176.285 ;
        RECT -41.645 174.595 -41.315 174.925 ;
        RECT -41.645 173.235 -41.315 173.565 ;
        RECT -41.645 171.875 -41.315 172.205 ;
        RECT -41.645 170.515 -41.315 170.845 ;
        RECT -41.645 169.155 -41.315 169.485 ;
        RECT -41.645 167.795 -41.315 168.125 ;
        RECT -41.645 166.435 -41.315 166.765 ;
        RECT -41.645 165.075 -41.315 165.405 ;
        RECT -41.645 163.715 -41.315 164.045 ;
        RECT -41.645 162.355 -41.315 162.685 ;
        RECT -41.645 160.995 -41.315 161.325 ;
        RECT -41.645 159.635 -41.315 159.965 ;
        RECT -41.645 158.275 -41.315 158.605 ;
        RECT -41.645 156.915 -41.315 157.245 ;
        RECT -41.645 155.555 -41.315 155.885 ;
        RECT -41.645 154.195 -41.315 154.525 ;
        RECT -41.645 152.835 -41.315 153.165 ;
        RECT -41.645 151.475 -41.315 151.805 ;
        RECT -41.645 150.115 -41.315 150.445 ;
        RECT -41.645 148.755 -41.315 149.085 ;
        RECT -41.645 147.395 -41.315 147.725 ;
        RECT -41.645 146.035 -41.315 146.365 ;
        RECT -41.645 144.675 -41.315 145.005 ;
        RECT -41.645 143.315 -41.315 143.645 ;
        RECT -41.645 141.955 -41.315 142.285 ;
        RECT -41.645 140.595 -41.315 140.925 ;
        RECT -41.645 139.235 -41.315 139.565 ;
        RECT -41.645 137.875 -41.315 138.205 ;
        RECT -41.645 136.515 -41.315 136.845 ;
        RECT -41.645 135.155 -41.315 135.485 ;
        RECT -41.645 133.795 -41.315 134.125 ;
        RECT -41.645 132.435 -41.315 132.765 ;
        RECT -41.645 131.075 -41.315 131.405 ;
        RECT -41.645 129.715 -41.315 130.045 ;
        RECT -41.645 128.355 -41.315 128.685 ;
        RECT -41.645 126.995 -41.315 127.325 ;
        RECT -41.645 125.635 -41.315 125.965 ;
        RECT -41.645 124.275 -41.315 124.605 ;
        RECT -41.645 122.915 -41.315 123.245 ;
        RECT -41.645 121.555 -41.315 121.885 ;
        RECT -41.645 120.195 -41.315 120.525 ;
        RECT -41.645 118.835 -41.315 119.165 ;
        RECT -41.645 117.475 -41.315 117.805 ;
        RECT -41.645 116.115 -41.315 116.445 ;
        RECT -41.645 114.755 -41.315 115.085 ;
        RECT -41.645 113.395 -41.315 113.725 ;
        RECT -41.645 112.035 -41.315 112.365 ;
        RECT -41.645 110.675 -41.315 111.005 ;
        RECT -41.645 109.315 -41.315 109.645 ;
        RECT -41.645 107.955 -41.315 108.285 ;
        RECT -41.645 106.595 -41.315 106.925 ;
        RECT -41.645 105.235 -41.315 105.565 ;
        RECT -41.645 103.875 -41.315 104.205 ;
        RECT -41.645 102.515 -41.315 102.845 ;
    END
    PORT
      LAYER met3 ;
        RECT -49.805 244.04 -49.475 245.17 ;
        RECT -49.805 239.875 -49.475 240.205 ;
        RECT -49.805 238.515 -49.475 238.845 ;
        RECT -49.805 237.155 -49.475 237.485 ;
        RECT -49.805 235.795 -49.475 236.125 ;
        RECT -49.805 234.435 -49.475 234.765 ;
        RECT -49.805 233.075 -49.475 233.405 ;
        RECT -49.805 231.715 -49.475 232.045 ;
        RECT -49.805 230.355 -49.475 230.685 ;
        RECT -49.805 228.995 -49.475 229.325 ;
        RECT -49.805 227.635 -49.475 227.965 ;
        RECT -49.805 226.275 -49.475 226.605 ;
        RECT -49.805 224.915 -49.475 225.245 ;
        RECT -49.805 223.555 -49.475 223.885 ;
        RECT -49.805 222.195 -49.475 222.525 ;
        RECT -49.805 220.835 -49.475 221.165 ;
        RECT -49.805 219.475 -49.475 219.805 ;
        RECT -49.805 218.115 -49.475 218.445 ;
        RECT -49.805 216.755 -49.475 217.085 ;
        RECT -49.805 215.395 -49.475 215.725 ;
        RECT -49.805 214.035 -49.475 214.365 ;
        RECT -49.805 212.675 -49.475 213.005 ;
        RECT -49.805 211.315 -49.475 211.645 ;
        RECT -49.805 209.955 -49.475 210.285 ;
        RECT -49.805 208.595 -49.475 208.925 ;
        RECT -49.805 207.235 -49.475 207.565 ;
        RECT -49.805 205.875 -49.475 206.205 ;
        RECT -49.805 204.515 -49.475 204.845 ;
        RECT -49.805 203.155 -49.475 203.485 ;
        RECT -49.805 201.795 -49.475 202.125 ;
        RECT -49.805 200.435 -49.475 200.765 ;
        RECT -49.805 199.075 -49.475 199.405 ;
        RECT -49.805 197.715 -49.475 198.045 ;
        RECT -49.805 196.355 -49.475 196.685 ;
        RECT -49.805 194.995 -49.475 195.325 ;
        RECT -49.805 193.635 -49.475 193.965 ;
        RECT -49.805 192.275 -49.475 192.605 ;
        RECT -49.805 190.915 -49.475 191.245 ;
        RECT -49.805 189.555 -49.475 189.885 ;
        RECT -49.805 188.195 -49.475 188.525 ;
        RECT -49.805 186.835 -49.475 187.165 ;
        RECT -49.805 185.475 -49.475 185.805 ;
        RECT -49.805 184.115 -49.475 184.445 ;
        RECT -49.805 182.755 -49.475 183.085 ;
        RECT -49.805 181.395 -49.475 181.725 ;
        RECT -49.805 180.035 -49.475 180.365 ;
        RECT -49.805 178.675 -49.475 179.005 ;
        RECT -49.805 177.315 -49.475 177.645 ;
        RECT -49.805 175.955 -49.475 176.285 ;
        RECT -49.805 174.595 -49.475 174.925 ;
        RECT -49.805 173.235 -49.475 173.565 ;
        RECT -49.805 171.875 -49.475 172.205 ;
        RECT -49.805 170.515 -49.475 170.845 ;
        RECT -49.805 169.155 -49.475 169.485 ;
        RECT -49.805 167.795 -49.475 168.125 ;
        RECT -49.805 166.435 -49.475 166.765 ;
        RECT -49.805 165.075 -49.475 165.405 ;
        RECT -49.805 163.715 -49.475 164.045 ;
        RECT -49.805 162.355 -49.475 162.685 ;
        RECT -49.805 160.995 -49.475 161.325 ;
        RECT -49.805 159.635 -49.475 159.965 ;
        RECT -49.805 158.275 -49.475 158.605 ;
        RECT -49.805 156.915 -49.475 157.245 ;
        RECT -49.805 155.555 -49.475 155.885 ;
        RECT -49.805 154.195 -49.475 154.525 ;
        RECT -49.805 152.835 -49.475 153.165 ;
        RECT -49.805 151.475 -49.475 151.805 ;
        RECT -49.805 150.115 -49.475 150.445 ;
        RECT -49.805 148.755 -49.475 149.085 ;
        RECT -49.805 147.395 -49.475 147.725 ;
        RECT -49.805 146.035 -49.475 146.365 ;
        RECT -49.805 144.675 -49.475 145.005 ;
        RECT -49.805 143.315 -49.475 143.645 ;
        RECT -49.805 141.955 -49.475 142.285 ;
        RECT -49.805 140.595 -49.475 140.925 ;
        RECT -49.805 139.235 -49.475 139.565 ;
        RECT -49.805 136.42 -49.475 136.75 ;
        RECT -49.805 134.245 -49.475 134.575 ;
        RECT -49.805 133.395 -49.475 133.725 ;
        RECT -49.805 131.085 -49.475 131.415 ;
        RECT -49.805 130.235 -49.475 130.565 ;
        RECT -49.805 127.925 -49.475 128.255 ;
        RECT -49.805 127.075 -49.475 127.405 ;
        RECT -49.805 124.765 -49.475 125.095 ;
        RECT -49.805 123.915 -49.475 124.245 ;
        RECT -49.805 121.605 -49.475 121.935 ;
        RECT -49.805 120.755 -49.475 121.085 ;
        RECT -49.805 118.445 -49.475 118.775 ;
        RECT -49.805 117.595 -49.475 117.925 ;
        RECT -49.805 115.285 -49.475 115.615 ;
        RECT -49.805 114.435 -49.475 114.765 ;
        RECT -49.805 112.125 -49.475 112.455 ;
        RECT -49.805 111.275 -49.475 111.605 ;
        RECT -49.805 108.965 -49.475 109.295 ;
        RECT -49.805 108.115 -49.475 108.445 ;
        RECT -49.805 105.805 -49.475 106.135 ;
        RECT -49.805 104.955 -49.475 105.285 ;
        RECT -49.805 102.645 -49.475 102.975 ;
        RECT -49.805 101.795 -49.475 102.125 ;
        RECT -49.805 99.62 -49.475 99.95 ;
        RECT -49.805 97.075 -49.475 97.405 ;
        RECT -49.805 95.715 -49.475 96.045 ;
        RECT -49.805 94.355 -49.475 94.685 ;
        RECT -49.805 92.995 -49.475 93.325 ;
        RECT -49.805 91.635 -49.475 91.965 ;
        RECT -49.805 90.275 -49.475 90.605 ;
        RECT -49.805 88.915 -49.475 89.245 ;
        RECT -49.805 87.555 -49.475 87.885 ;
        RECT -49.805 86.195 -49.475 86.525 ;
        RECT -49.805 84.835 -49.475 85.165 ;
        RECT -49.805 83.475 -49.475 83.805 ;
        RECT -49.805 82.115 -49.475 82.445 ;
        RECT -49.805 80.755 -49.475 81.085 ;
        RECT -49.805 79.395 -49.475 79.725 ;
        RECT -49.805 78.035 -49.475 78.365 ;
        RECT -49.805 76.675 -49.475 77.005 ;
        RECT -49.805 75.315 -49.475 75.645 ;
        RECT -49.805 73.955 -49.475 74.285 ;
        RECT -49.805 72.595 -49.475 72.925 ;
        RECT -49.805 71.235 -49.475 71.565 ;
        RECT -49.805 69.875 -49.475 70.205 ;
        RECT -49.805 68.515 -49.475 68.845 ;
        RECT -49.805 67.155 -49.475 67.485 ;
        RECT -49.805 65.795 -49.475 66.125 ;
        RECT -49.805 64.435 -49.475 64.765 ;
        RECT -49.805 63.075 -49.475 63.405 ;
        RECT -49.805 61.715 -49.475 62.045 ;
        RECT -49.805 60.355 -49.475 60.685 ;
        RECT -49.805 58.995 -49.475 59.325 ;
        RECT -49.805 57.635 -49.475 57.965 ;
        RECT -49.805 56.275 -49.475 56.605 ;
        RECT -49.805 54.915 -49.475 55.245 ;
        RECT -49.805 53.555 -49.475 53.885 ;
        RECT -49.805 52.195 -49.475 52.525 ;
        RECT -49.805 50.835 -49.475 51.165 ;
        RECT -49.805 49.475 -49.475 49.805 ;
        RECT -49.805 48.115 -49.475 48.445 ;
        RECT -49.805 46.755 -49.475 47.085 ;
        RECT -49.805 45.395 -49.475 45.725 ;
        RECT -49.805 44.035 -49.475 44.365 ;
        RECT -49.805 42.675 -49.475 43.005 ;
        RECT -49.805 41.315 -49.475 41.645 ;
        RECT -49.805 39.955 -49.475 40.285 ;
        RECT -49.805 38.595 -49.475 38.925 ;
        RECT -49.805 37.235 -49.475 37.565 ;
        RECT -49.805 35.875 -49.475 36.205 ;
        RECT -49.805 34.515 -49.475 34.845 ;
        RECT -49.805 33.155 -49.475 33.485 ;
        RECT -49.805 31.795 -49.475 32.125 ;
        RECT -49.805 30.435 -49.475 30.765 ;
        RECT -49.805 29.075 -49.475 29.405 ;
        RECT -49.805 27.715 -49.475 28.045 ;
        RECT -49.805 26.355 -49.475 26.685 ;
        RECT -49.805 24.995 -49.475 25.325 ;
        RECT -49.805 23.635 -49.475 23.965 ;
        RECT -49.805 22.275 -49.475 22.605 ;
        RECT -49.805 20.915 -49.475 21.245 ;
        RECT -49.805 19.555 -49.475 19.885 ;
        RECT -49.805 18.195 -49.475 18.525 ;
        RECT -49.805 16.835 -49.475 17.165 ;
        RECT -49.805 15.475 -49.475 15.805 ;
        RECT -49.805 14.115 -49.475 14.445 ;
        RECT -49.805 12.755 -49.475 13.085 ;
        RECT -49.805 11.395 -49.475 11.725 ;
        RECT -49.805 10.035 -49.475 10.365 ;
        RECT -49.805 8.675 -49.475 9.005 ;
        RECT -49.805 7.315 -49.475 7.645 ;
        RECT -49.805 5.955 -49.475 6.285 ;
        RECT -49.805 4.595 -49.475 4.925 ;
        RECT -49.805 3.235 -49.475 3.565 ;
        RECT -49.805 1.875 -49.475 2.205 ;
        RECT -49.805 0.515 -49.475 0.845 ;
        RECT -49.805 -0.845 -49.475 -0.515 ;
        RECT -49.805 -2.205 -49.475 -1.875 ;
        RECT -49.805 -3.565 -49.475 -3.235 ;
        RECT -49.805 -4.925 -49.475 -4.595 ;
        RECT -49.805 -6.285 -49.475 -5.955 ;
        RECT -49.805 -7.645 -49.475 -7.315 ;
        RECT -49.805 -9.005 -49.475 -8.675 ;
        RECT -49.805 -10.365 -49.475 -10.035 ;
        RECT -49.805 -11.725 -49.475 -11.395 ;
        RECT -49.805 -14.445 -49.475 -14.115 ;
        RECT -49.805 -15.805 -49.475 -15.475 ;
        RECT -49.805 -17.165 -49.475 -16.835 ;
        RECT -49.805 -18.525 -49.475 -18.195 ;
        RECT -49.805 -19.885 -49.475 -19.555 ;
        RECT -49.805 -21.245 -49.475 -20.915 ;
        RECT -49.805 -22.605 -49.475 -22.275 ;
        RECT -49.805 -23.965 -49.475 -23.635 ;
        RECT -49.805 -25.325 -49.475 -24.995 ;
        RECT -49.805 -29.405 -49.475 -29.075 ;
        RECT -49.805 -30.765 -49.475 -30.435 ;
        RECT -49.805 -32.125 -49.475 -31.795 ;
        RECT -49.805 -34.845 -49.475 -34.515 ;
        RECT -49.805 -36.205 -49.475 -35.875 ;
        RECT -49.805 -38.925 -49.475 -38.595 ;
        RECT -49.805 -41.645 -49.475 -41.315 ;
        RECT -49.805 -44.365 -49.475 -44.035 ;
        RECT -49.805 -49.805 -49.475 -49.475 ;
        RECT -49.805 -51.165 -49.475 -50.835 ;
        RECT -49.805 -53.885 -49.475 -53.555 ;
        RECT -49.805 -55.245 -49.475 -54.915 ;
        RECT -49.805 -59.325 -49.475 -58.995 ;
        RECT -49.805 -60.685 -49.475 -60.355 ;
        RECT -49.805 -63.405 -49.475 -63.075 ;
        RECT -49.805 -67.485 -49.475 -67.155 ;
        RECT -49.805 -68.845 -49.475 -68.515 ;
        RECT -49.805 -70.205 -49.475 -69.875 ;
        RECT -49.805 -71.565 -49.475 -71.235 ;
        RECT -49.805 -72.925 -49.475 -72.595 ;
        RECT -49.805 -74.285 -49.475 -73.955 ;
        RECT -49.805 -75.645 -49.475 -75.315 ;
        RECT -49.805 -77.005 -49.475 -76.675 ;
        RECT -49.805 -78.365 -49.475 -78.035 ;
        RECT -49.805 -79.725 -49.475 -79.395 ;
        RECT -49.805 -81.085 -49.475 -80.755 ;
        RECT -49.805 -82.445 -49.475 -82.115 ;
        RECT -49.805 -83.805 -49.475 -83.475 ;
        RECT -49.805 -85.165 -49.475 -84.835 ;
        RECT -49.805 -86.525 -49.475 -86.195 ;
        RECT -49.805 -87.885 -49.475 -87.555 ;
        RECT -49.805 -89.245 -49.475 -88.915 ;
        RECT -49.805 -90.81 -49.475 -90.48 ;
        RECT -49.805 -91.965 -49.475 -91.635 ;
        RECT -49.805 -93.325 -49.475 -92.995 ;
        RECT -49.805 -94.685 -49.475 -94.355 ;
        RECT -49.805 -96.045 -49.475 -95.715 ;
        RECT -49.805 -97.405 -49.475 -97.075 ;
        RECT -49.805 -100.125 -49.475 -99.795 ;
        RECT -49.805 -101.35 -49.475 -101.02 ;
        RECT -49.805 -102.845 -49.475 -102.515 ;
        RECT -49.805 -104.205 -49.475 -103.875 ;
        RECT -49.805 -105.565 -49.475 -105.235 ;
        RECT -49.805 -108.285 -49.475 -107.955 ;
        RECT -49.805 -109.645 -49.475 -109.315 ;
        RECT -49.805 -113.725 -49.475 -113.395 ;
        RECT -49.805 -115.085 -49.475 -114.755 ;
        RECT -49.805 -116.445 -49.475 -116.115 ;
        RECT -49.805 -117.805 -49.475 -117.475 ;
        RECT -49.805 -119.165 -49.475 -118.835 ;
        RECT -49.805 -120.525 -49.475 -120.195 ;
        RECT -49.805 -121.885 -49.475 -121.555 ;
        RECT -49.805 -123.245 -49.475 -122.915 ;
        RECT -49.805 -124.605 -49.475 -124.275 ;
        RECT -49.805 -125.965 -49.475 -125.635 ;
        RECT -49.805 -127.325 -49.475 -126.995 ;
        RECT -49.805 -128.685 -49.475 -128.355 ;
        RECT -49.805 -130.045 -49.475 -129.715 ;
        RECT -49.805 -131.405 -49.475 -131.075 ;
        RECT -49.805 -132.765 -49.475 -132.435 ;
        RECT -49.805 -134.125 -49.475 -133.795 ;
        RECT -49.805 -135.485 -49.475 -135.155 ;
        RECT -49.805 -136.845 -49.475 -136.515 ;
        RECT -49.805 -138.205 -49.475 -137.875 ;
        RECT -49.805 -139.565 -49.475 -139.235 ;
        RECT -49.805 -140.925 -49.475 -140.595 ;
        RECT -49.805 -142.285 -49.475 -141.955 ;
        RECT -49.805 -143.645 -49.475 -143.315 ;
        RECT -49.805 -145.005 -49.475 -144.675 ;
        RECT -49.805 -146.365 -49.475 -146.035 ;
        RECT -49.805 -147.725 -49.475 -147.395 ;
        RECT -49.805 -149.085 -49.475 -148.755 ;
        RECT -49.805 -150.445 -49.475 -150.115 ;
        RECT -49.805 -151.805 -49.475 -151.475 ;
        RECT -49.805 -153.165 -49.475 -152.835 ;
        RECT -49.805 -154.525 -49.475 -154.195 ;
        RECT -49.805 -155.885 -49.475 -155.555 ;
        RECT -49.805 -157.245 -49.475 -156.915 ;
        RECT -49.805 -158.605 -49.475 -158.275 ;
        RECT -49.805 -159.965 -49.475 -159.635 ;
        RECT -49.805 -161.325 -49.475 -160.995 ;
        RECT -49.805 -162.685 -49.475 -162.355 ;
        RECT -49.805 -164.045 -49.475 -163.715 ;
        RECT -49.805 -165.405 -49.475 -165.075 ;
        RECT -49.805 -166.765 -49.475 -166.435 ;
        RECT -49.805 -168.655 -49.475 -168.325 ;
        RECT -49.805 -169.485 -49.475 -169.155 ;
        RECT -49.805 -170.845 -49.475 -170.515 ;
        RECT -49.805 -172.205 -49.475 -171.875 ;
        RECT -49.805 -173.565 -49.475 -173.235 ;
        RECT -49.805 -174.925 -49.475 -174.595 ;
        RECT -49.805 -177.645 -49.475 -177.315 ;
        RECT -49.805 -183.29 -49.475 -182.16 ;
        RECT -49.8 -183.405 -49.48 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -48.445 244.04 -48.115 245.17 ;
        RECT -48.445 239.875 -48.115 240.205 ;
        RECT -48.445 238.515 -48.115 238.845 ;
        RECT -48.445 237.155 -48.115 237.485 ;
        RECT -48.445 235.795 -48.115 236.125 ;
        RECT -48.445 234.435 -48.115 234.765 ;
        RECT -48.445 233.075 -48.115 233.405 ;
        RECT -48.445 231.715 -48.115 232.045 ;
        RECT -48.445 230.355 -48.115 230.685 ;
        RECT -48.445 228.995 -48.115 229.325 ;
        RECT -48.445 227.635 -48.115 227.965 ;
        RECT -48.445 226.275 -48.115 226.605 ;
        RECT -48.445 224.915 -48.115 225.245 ;
        RECT -48.445 223.555 -48.115 223.885 ;
        RECT -48.445 222.195 -48.115 222.525 ;
        RECT -48.445 220.835 -48.115 221.165 ;
        RECT -48.445 219.475 -48.115 219.805 ;
        RECT -48.445 218.115 -48.115 218.445 ;
        RECT -48.445 216.755 -48.115 217.085 ;
        RECT -48.445 215.395 -48.115 215.725 ;
        RECT -48.445 214.035 -48.115 214.365 ;
        RECT -48.445 212.675 -48.115 213.005 ;
        RECT -48.445 211.315 -48.115 211.645 ;
        RECT -48.445 209.955 -48.115 210.285 ;
        RECT -48.445 208.595 -48.115 208.925 ;
        RECT -48.445 207.235 -48.115 207.565 ;
        RECT -48.445 205.875 -48.115 206.205 ;
        RECT -48.445 204.515 -48.115 204.845 ;
        RECT -48.445 203.155 -48.115 203.485 ;
        RECT -48.445 201.795 -48.115 202.125 ;
        RECT -48.445 200.435 -48.115 200.765 ;
        RECT -48.445 199.075 -48.115 199.405 ;
        RECT -48.445 197.715 -48.115 198.045 ;
        RECT -48.445 196.355 -48.115 196.685 ;
        RECT -48.445 194.995 -48.115 195.325 ;
        RECT -48.445 193.635 -48.115 193.965 ;
        RECT -48.445 192.275 -48.115 192.605 ;
        RECT -48.445 190.915 -48.115 191.245 ;
        RECT -48.445 189.555 -48.115 189.885 ;
        RECT -48.445 188.195 -48.115 188.525 ;
        RECT -48.445 186.835 -48.115 187.165 ;
        RECT -48.445 185.475 -48.115 185.805 ;
        RECT -48.445 184.115 -48.115 184.445 ;
        RECT -48.445 182.755 -48.115 183.085 ;
        RECT -48.445 181.395 -48.115 181.725 ;
        RECT -48.445 180.035 -48.115 180.365 ;
        RECT -48.445 178.675 -48.115 179.005 ;
        RECT -48.445 177.315 -48.115 177.645 ;
        RECT -48.445 175.955 -48.115 176.285 ;
        RECT -48.445 174.595 -48.115 174.925 ;
        RECT -48.445 173.235 -48.115 173.565 ;
        RECT -48.445 171.875 -48.115 172.205 ;
        RECT -48.445 170.515 -48.115 170.845 ;
        RECT -48.445 169.155 -48.115 169.485 ;
        RECT -48.445 167.795 -48.115 168.125 ;
        RECT -48.445 166.435 -48.115 166.765 ;
        RECT -48.445 165.075 -48.115 165.405 ;
        RECT -48.445 163.715 -48.115 164.045 ;
        RECT -48.445 162.355 -48.115 162.685 ;
        RECT -48.445 160.995 -48.115 161.325 ;
        RECT -48.445 159.635 -48.115 159.965 ;
        RECT -48.445 158.275 -48.115 158.605 ;
        RECT -48.445 156.915 -48.115 157.245 ;
        RECT -48.445 155.555 -48.115 155.885 ;
        RECT -48.445 154.195 -48.115 154.525 ;
        RECT -48.445 152.835 -48.115 153.165 ;
        RECT -48.445 151.475 -48.115 151.805 ;
        RECT -48.445 150.115 -48.115 150.445 ;
        RECT -48.445 148.755 -48.115 149.085 ;
        RECT -48.445 147.395 -48.115 147.725 ;
        RECT -48.445 146.035 -48.115 146.365 ;
        RECT -48.445 144.675 -48.115 145.005 ;
        RECT -48.445 143.315 -48.115 143.645 ;
        RECT -48.445 141.955 -48.115 142.285 ;
        RECT -48.445 140.595 -48.115 140.925 ;
        RECT -48.445 139.235 -48.115 139.565 ;
        RECT -48.445 136.42 -48.115 136.75 ;
        RECT -48.445 134.245 -48.115 134.575 ;
        RECT -48.445 133.395 -48.115 133.725 ;
        RECT -48.445 131.085 -48.115 131.415 ;
        RECT -48.445 130.235 -48.115 130.565 ;
        RECT -48.445 127.925 -48.115 128.255 ;
        RECT -48.445 127.075 -48.115 127.405 ;
        RECT -48.445 124.765 -48.115 125.095 ;
        RECT -48.445 123.915 -48.115 124.245 ;
        RECT -48.445 121.605 -48.115 121.935 ;
        RECT -48.445 120.755 -48.115 121.085 ;
        RECT -48.445 118.445 -48.115 118.775 ;
        RECT -48.445 117.595 -48.115 117.925 ;
        RECT -48.445 115.285 -48.115 115.615 ;
        RECT -48.445 114.435 -48.115 114.765 ;
        RECT -48.445 112.125 -48.115 112.455 ;
        RECT -48.445 111.275 -48.115 111.605 ;
        RECT -48.445 108.965 -48.115 109.295 ;
        RECT -48.445 108.115 -48.115 108.445 ;
        RECT -48.445 105.805 -48.115 106.135 ;
        RECT -48.445 104.955 -48.115 105.285 ;
        RECT -48.445 102.645 -48.115 102.975 ;
        RECT -48.445 101.795 -48.115 102.125 ;
        RECT -48.445 99.62 -48.115 99.95 ;
        RECT -48.445 97.075 -48.115 97.405 ;
        RECT -48.445 95.715 -48.115 96.045 ;
        RECT -48.445 94.355 -48.115 94.685 ;
        RECT -48.445 92.995 -48.115 93.325 ;
        RECT -48.445 91.635 -48.115 91.965 ;
        RECT -48.445 90.275 -48.115 90.605 ;
        RECT -48.445 88.915 -48.115 89.245 ;
        RECT -48.445 87.555 -48.115 87.885 ;
        RECT -48.445 86.195 -48.115 86.525 ;
        RECT -48.445 84.835 -48.115 85.165 ;
        RECT -48.445 83.475 -48.115 83.805 ;
        RECT -48.445 82.115 -48.115 82.445 ;
        RECT -48.445 80.755 -48.115 81.085 ;
        RECT -48.445 79.395 -48.115 79.725 ;
        RECT -48.445 78.035 -48.115 78.365 ;
        RECT -48.445 76.675 -48.115 77.005 ;
        RECT -48.445 75.315 -48.115 75.645 ;
        RECT -48.445 73.955 -48.115 74.285 ;
        RECT -48.445 72.595 -48.115 72.925 ;
        RECT -48.445 71.235 -48.115 71.565 ;
        RECT -48.445 69.875 -48.115 70.205 ;
        RECT -48.445 68.515 -48.115 68.845 ;
        RECT -48.445 67.155 -48.115 67.485 ;
        RECT -48.445 65.795 -48.115 66.125 ;
        RECT -48.445 64.435 -48.115 64.765 ;
        RECT -48.445 63.075 -48.115 63.405 ;
        RECT -48.445 61.715 -48.115 62.045 ;
        RECT -48.445 60.355 -48.115 60.685 ;
        RECT -48.445 58.995 -48.115 59.325 ;
        RECT -48.445 57.635 -48.115 57.965 ;
        RECT -48.445 56.275 -48.115 56.605 ;
        RECT -48.445 54.915 -48.115 55.245 ;
        RECT -48.445 53.555 -48.115 53.885 ;
        RECT -48.445 52.195 -48.115 52.525 ;
        RECT -48.445 50.835 -48.115 51.165 ;
        RECT -48.445 49.475 -48.115 49.805 ;
        RECT -48.445 48.115 -48.115 48.445 ;
        RECT -48.445 46.755 -48.115 47.085 ;
        RECT -48.445 45.395 -48.115 45.725 ;
        RECT -48.445 44.035 -48.115 44.365 ;
        RECT -48.445 42.675 -48.115 43.005 ;
        RECT -48.445 41.315 -48.115 41.645 ;
        RECT -48.445 39.955 -48.115 40.285 ;
        RECT -48.445 38.595 -48.115 38.925 ;
        RECT -48.445 37.235 -48.115 37.565 ;
        RECT -48.445 35.875 -48.115 36.205 ;
        RECT -48.445 34.515 -48.115 34.845 ;
        RECT -48.445 33.155 -48.115 33.485 ;
        RECT -48.445 31.795 -48.115 32.125 ;
        RECT -48.445 30.435 -48.115 30.765 ;
        RECT -48.445 29.075 -48.115 29.405 ;
        RECT -48.445 27.715 -48.115 28.045 ;
        RECT -48.445 26.355 -48.115 26.685 ;
        RECT -48.445 24.995 -48.115 25.325 ;
        RECT -48.445 23.635 -48.115 23.965 ;
        RECT -48.445 22.275 -48.115 22.605 ;
        RECT -48.445 20.915 -48.115 21.245 ;
        RECT -48.445 19.555 -48.115 19.885 ;
        RECT -48.445 18.195 -48.115 18.525 ;
        RECT -48.445 16.835 -48.115 17.165 ;
        RECT -48.445 15.475 -48.115 15.805 ;
        RECT -48.445 14.115 -48.115 14.445 ;
        RECT -48.445 12.755 -48.115 13.085 ;
        RECT -48.445 11.395 -48.115 11.725 ;
        RECT -48.445 10.035 -48.115 10.365 ;
        RECT -48.445 8.675 -48.115 9.005 ;
        RECT -48.445 7.315 -48.115 7.645 ;
        RECT -48.445 5.955 -48.115 6.285 ;
        RECT -48.445 4.595 -48.115 4.925 ;
        RECT -48.445 3.235 -48.115 3.565 ;
        RECT -48.445 1.875 -48.115 2.205 ;
        RECT -48.445 0.515 -48.115 0.845 ;
        RECT -48.445 -0.845 -48.115 -0.515 ;
        RECT -48.445 -2.205 -48.115 -1.875 ;
        RECT -48.445 -3.565 -48.115 -3.235 ;
        RECT -48.445 -4.925 -48.115 -4.595 ;
        RECT -48.445 -6.285 -48.115 -5.955 ;
        RECT -48.445 -7.645 -48.115 -7.315 ;
        RECT -48.445 -9.005 -48.115 -8.675 ;
        RECT -48.445 -10.365 -48.115 -10.035 ;
        RECT -48.445 -14.445 -48.115 -14.115 ;
        RECT -48.445 -15.805 -48.115 -15.475 ;
        RECT -48.445 -17.165 -48.115 -16.835 ;
        RECT -48.445 -18.525 -48.115 -18.195 ;
        RECT -48.445 -19.885 -48.115 -19.555 ;
        RECT -48.445 -21.245 -48.115 -20.915 ;
        RECT -48.445 -22.605 -48.115 -22.275 ;
        RECT -48.445 -23.965 -48.115 -23.635 ;
        RECT -48.445 -25.325 -48.115 -24.995 ;
        RECT -48.445 -29.405 -48.115 -29.075 ;
        RECT -48.445 -32.125 -48.115 -31.795 ;
        RECT -48.445 -33.71 -48.115 -33.38 ;
        RECT -48.445 -34.845 -48.115 -34.515 ;
        RECT -48.445 -36.205 -48.115 -35.875 ;
        RECT -48.445 -38.925 -48.115 -38.595 ;
        RECT -48.445 -39.75 -48.115 -39.42 ;
        RECT -48.445 -41.645 -48.115 -41.315 ;
        RECT -48.445 -44.365 -48.115 -44.035 ;
        RECT -48.445 -49.805 -48.115 -49.475 ;
        RECT -48.445 -51.165 -48.115 -50.835 ;
        RECT -48.445 -53.885 -48.115 -53.555 ;
        RECT -48.445 -55.245 -48.115 -54.915 ;
        RECT -48.445 -59.325 -48.115 -58.995 ;
        RECT -48.445 -60.685 -48.115 -60.355 ;
        RECT -48.445 -67.485 -48.115 -67.155 ;
        RECT -48.445 -68.845 -48.115 -68.515 ;
        RECT -48.445 -70.205 -48.115 -69.875 ;
        RECT -48.445 -71.565 -48.115 -71.235 ;
        RECT -48.445 -72.925 -48.115 -72.595 ;
        RECT -48.445 -74.285 -48.115 -73.955 ;
        RECT -48.445 -75.645 -48.115 -75.315 ;
        RECT -48.445 -77.005 -48.115 -76.675 ;
        RECT -48.445 -78.365 -48.115 -78.035 ;
        RECT -48.445 -79.725 -48.115 -79.395 ;
        RECT -48.445 -81.085 -48.115 -80.755 ;
        RECT -48.445 -82.445 -48.115 -82.115 ;
        RECT -48.445 -83.805 -48.115 -83.475 ;
        RECT -48.445 -85.165 -48.115 -84.835 ;
        RECT -48.445 -86.525 -48.115 -86.195 ;
        RECT -48.445 -87.885 -48.115 -87.555 ;
        RECT -48.445 -89.245 -48.115 -88.915 ;
        RECT -48.445 -90.81 -48.115 -90.48 ;
        RECT -48.445 -91.965 -48.115 -91.635 ;
        RECT -48.445 -93.325 -48.115 -92.995 ;
        RECT -48.445 -94.685 -48.115 -94.355 ;
        RECT -48.445 -96.045 -48.115 -95.715 ;
        RECT -48.445 -97.405 -48.115 -97.075 ;
        RECT -48.445 -100.125 -48.115 -99.795 ;
        RECT -48.445 -101.35 -48.115 -101.02 ;
        RECT -48.445 -102.845 -48.115 -102.515 ;
        RECT -48.445 -104.205 -48.115 -103.875 ;
        RECT -48.445 -105.565 -48.115 -105.235 ;
        RECT -48.445 -108.285 -48.115 -107.955 ;
        RECT -48.445 -109.645 -48.115 -109.315 ;
        RECT -48.445 -112.365 -48.115 -112.035 ;
        RECT -48.44 -113.04 -48.12 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -48.445 -174.925 -48.115 -174.595 ;
        RECT -48.445 -177.645 -48.115 -177.315 ;
        RECT -48.445 -183.29 -48.115 -182.16 ;
        RECT -48.44 -183.405 -48.12 -173.92 ;
    END
    PORT
      LAYER met3 ;
        RECT -47.085 244.04 -46.755 245.17 ;
        RECT -47.085 239.875 -46.755 240.205 ;
        RECT -47.085 238.515 -46.755 238.845 ;
        RECT -47.085 237.155 -46.755 237.485 ;
        RECT -47.085 235.795 -46.755 236.125 ;
        RECT -47.085 234.435 -46.755 234.765 ;
        RECT -47.085 233.075 -46.755 233.405 ;
        RECT -47.085 231.715 -46.755 232.045 ;
        RECT -47.085 230.355 -46.755 230.685 ;
        RECT -47.085 228.995 -46.755 229.325 ;
        RECT -47.085 227.635 -46.755 227.965 ;
        RECT -47.085 226.275 -46.755 226.605 ;
        RECT -47.085 224.915 -46.755 225.245 ;
        RECT -47.085 223.555 -46.755 223.885 ;
        RECT -47.085 222.195 -46.755 222.525 ;
        RECT -47.085 220.835 -46.755 221.165 ;
        RECT -47.085 219.475 -46.755 219.805 ;
        RECT -47.085 218.115 -46.755 218.445 ;
        RECT -47.085 216.755 -46.755 217.085 ;
        RECT -47.085 215.395 -46.755 215.725 ;
        RECT -47.085 214.035 -46.755 214.365 ;
        RECT -47.085 212.675 -46.755 213.005 ;
        RECT -47.085 211.315 -46.755 211.645 ;
        RECT -47.085 209.955 -46.755 210.285 ;
        RECT -47.085 208.595 -46.755 208.925 ;
        RECT -47.085 207.235 -46.755 207.565 ;
        RECT -47.085 205.875 -46.755 206.205 ;
        RECT -47.085 204.515 -46.755 204.845 ;
        RECT -47.085 203.155 -46.755 203.485 ;
        RECT -47.085 201.795 -46.755 202.125 ;
        RECT -47.085 200.435 -46.755 200.765 ;
        RECT -47.085 199.075 -46.755 199.405 ;
        RECT -47.085 197.715 -46.755 198.045 ;
        RECT -47.085 196.355 -46.755 196.685 ;
        RECT -47.085 194.995 -46.755 195.325 ;
        RECT -47.085 193.635 -46.755 193.965 ;
        RECT -47.085 192.275 -46.755 192.605 ;
        RECT -47.085 190.915 -46.755 191.245 ;
        RECT -47.085 189.555 -46.755 189.885 ;
        RECT -47.085 188.195 -46.755 188.525 ;
        RECT -47.085 186.835 -46.755 187.165 ;
        RECT -47.085 185.475 -46.755 185.805 ;
        RECT -47.085 184.115 -46.755 184.445 ;
        RECT -47.085 182.755 -46.755 183.085 ;
        RECT -47.085 181.395 -46.755 181.725 ;
        RECT -47.085 180.035 -46.755 180.365 ;
        RECT -47.085 178.675 -46.755 179.005 ;
        RECT -47.085 177.315 -46.755 177.645 ;
        RECT -47.085 175.955 -46.755 176.285 ;
        RECT -47.085 174.595 -46.755 174.925 ;
        RECT -47.085 173.235 -46.755 173.565 ;
        RECT -47.085 171.875 -46.755 172.205 ;
        RECT -47.085 170.515 -46.755 170.845 ;
        RECT -47.085 169.155 -46.755 169.485 ;
        RECT -47.085 167.795 -46.755 168.125 ;
        RECT -47.085 166.435 -46.755 166.765 ;
        RECT -47.085 165.075 -46.755 165.405 ;
        RECT -47.085 163.715 -46.755 164.045 ;
        RECT -47.085 162.355 -46.755 162.685 ;
        RECT -47.085 160.995 -46.755 161.325 ;
        RECT -47.085 159.635 -46.755 159.965 ;
        RECT -47.085 158.275 -46.755 158.605 ;
        RECT -47.085 156.915 -46.755 157.245 ;
        RECT -47.085 155.555 -46.755 155.885 ;
        RECT -47.085 154.195 -46.755 154.525 ;
        RECT -47.085 152.835 -46.755 153.165 ;
        RECT -47.085 151.475 -46.755 151.805 ;
        RECT -47.085 150.115 -46.755 150.445 ;
        RECT -47.085 148.755 -46.755 149.085 ;
        RECT -47.085 147.395 -46.755 147.725 ;
        RECT -47.085 146.035 -46.755 146.365 ;
        RECT -47.085 144.675 -46.755 145.005 ;
        RECT -47.085 143.315 -46.755 143.645 ;
        RECT -47.085 141.955 -46.755 142.285 ;
        RECT -47.085 140.595 -46.755 140.925 ;
        RECT -47.085 139.235 -46.755 139.565 ;
        RECT -47.085 137.875 -46.755 138.205 ;
        RECT -47.085 136.515 -46.755 136.845 ;
        RECT -47.085 135.155 -46.755 135.485 ;
        RECT -47.085 133.795 -46.755 134.125 ;
        RECT -47.085 132.435 -46.755 132.765 ;
        RECT -47.085 131.075 -46.755 131.405 ;
        RECT -47.085 129.715 -46.755 130.045 ;
        RECT -47.085 128.355 -46.755 128.685 ;
        RECT -47.085 126.995 -46.755 127.325 ;
        RECT -47.085 125.635 -46.755 125.965 ;
        RECT -47.085 124.275 -46.755 124.605 ;
        RECT -47.085 122.915 -46.755 123.245 ;
        RECT -47.085 121.555 -46.755 121.885 ;
        RECT -47.085 120.195 -46.755 120.525 ;
        RECT -47.085 118.835 -46.755 119.165 ;
        RECT -47.085 117.475 -46.755 117.805 ;
        RECT -47.085 116.115 -46.755 116.445 ;
        RECT -47.085 114.755 -46.755 115.085 ;
        RECT -47.085 113.395 -46.755 113.725 ;
        RECT -47.085 112.035 -46.755 112.365 ;
        RECT -47.085 110.675 -46.755 111.005 ;
        RECT -47.085 109.315 -46.755 109.645 ;
        RECT -47.085 107.955 -46.755 108.285 ;
        RECT -47.085 106.595 -46.755 106.925 ;
        RECT -47.085 105.235 -46.755 105.565 ;
        RECT -47.085 103.875 -46.755 104.205 ;
        RECT -47.085 102.515 -46.755 102.845 ;
        RECT -47.085 101.155 -46.755 101.485 ;
        RECT -47.085 99.795 -46.755 100.125 ;
        RECT -47.085 98.435 -46.755 98.765 ;
        RECT -47.085 97.075 -46.755 97.405 ;
        RECT -47.085 95.715 -46.755 96.045 ;
        RECT -47.085 94.355 -46.755 94.685 ;
        RECT -47.085 92.995 -46.755 93.325 ;
        RECT -47.085 91.635 -46.755 91.965 ;
        RECT -47.085 90.275 -46.755 90.605 ;
        RECT -47.085 88.915 -46.755 89.245 ;
        RECT -47.085 87.555 -46.755 87.885 ;
        RECT -47.085 86.195 -46.755 86.525 ;
        RECT -47.085 84.835 -46.755 85.165 ;
        RECT -47.085 83.475 -46.755 83.805 ;
        RECT -47.085 82.115 -46.755 82.445 ;
        RECT -47.085 80.755 -46.755 81.085 ;
        RECT -47.085 79.395 -46.755 79.725 ;
        RECT -47.085 78.035 -46.755 78.365 ;
        RECT -47.085 76.675 -46.755 77.005 ;
        RECT -47.085 75.315 -46.755 75.645 ;
        RECT -47.085 73.955 -46.755 74.285 ;
        RECT -47.085 72.595 -46.755 72.925 ;
        RECT -47.085 71.235 -46.755 71.565 ;
        RECT -47.085 69.875 -46.755 70.205 ;
        RECT -47.085 68.515 -46.755 68.845 ;
        RECT -47.085 67.155 -46.755 67.485 ;
        RECT -47.085 65.795 -46.755 66.125 ;
        RECT -47.085 64.435 -46.755 64.765 ;
        RECT -47.085 63.075 -46.755 63.405 ;
        RECT -47.085 61.715 -46.755 62.045 ;
        RECT -47.085 60.355 -46.755 60.685 ;
        RECT -47.085 58.995 -46.755 59.325 ;
        RECT -47.085 57.635 -46.755 57.965 ;
        RECT -47.085 56.275 -46.755 56.605 ;
        RECT -47.085 54.915 -46.755 55.245 ;
        RECT -47.085 53.555 -46.755 53.885 ;
        RECT -47.085 52.195 -46.755 52.525 ;
        RECT -47.085 50.835 -46.755 51.165 ;
        RECT -47.085 49.475 -46.755 49.805 ;
        RECT -47.085 48.115 -46.755 48.445 ;
        RECT -47.085 46.755 -46.755 47.085 ;
        RECT -47.085 45.395 -46.755 45.725 ;
        RECT -47.085 44.035 -46.755 44.365 ;
        RECT -47.085 42.675 -46.755 43.005 ;
        RECT -47.085 41.315 -46.755 41.645 ;
        RECT -47.085 39.955 -46.755 40.285 ;
        RECT -47.085 38.595 -46.755 38.925 ;
        RECT -47.085 37.235 -46.755 37.565 ;
        RECT -47.085 35.875 -46.755 36.205 ;
        RECT -47.085 34.515 -46.755 34.845 ;
        RECT -47.085 33.155 -46.755 33.485 ;
        RECT -47.085 31.795 -46.755 32.125 ;
        RECT -47.085 30.435 -46.755 30.765 ;
        RECT -47.085 29.075 -46.755 29.405 ;
        RECT -47.085 27.715 -46.755 28.045 ;
        RECT -47.085 26.355 -46.755 26.685 ;
        RECT -47.085 24.995 -46.755 25.325 ;
        RECT -47.085 23.635 -46.755 23.965 ;
        RECT -47.085 22.275 -46.755 22.605 ;
        RECT -47.085 20.915 -46.755 21.245 ;
        RECT -47.085 19.555 -46.755 19.885 ;
        RECT -47.085 18.195 -46.755 18.525 ;
        RECT -47.085 16.835 -46.755 17.165 ;
        RECT -47.085 15.475 -46.755 15.805 ;
        RECT -47.085 14.115 -46.755 14.445 ;
        RECT -47.085 12.755 -46.755 13.085 ;
        RECT -47.085 11.395 -46.755 11.725 ;
        RECT -47.085 10.035 -46.755 10.365 ;
        RECT -47.085 8.675 -46.755 9.005 ;
        RECT -47.085 7.315 -46.755 7.645 ;
        RECT -47.085 5.955 -46.755 6.285 ;
        RECT -47.085 4.595 -46.755 4.925 ;
        RECT -47.085 3.235 -46.755 3.565 ;
        RECT -47.085 1.875 -46.755 2.205 ;
        RECT -47.085 0.515 -46.755 0.845 ;
        RECT -47.085 -0.845 -46.755 -0.515 ;
        RECT -47.08 -1.52 -46.76 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -47.085 -59.325 -46.755 -58.995 ;
        RECT -47.085 -60.685 -46.755 -60.355 ;
        RECT -47.085 -67.485 -46.755 -67.155 ;
        RECT -47.085 -68.845 -46.755 -68.515 ;
        RECT -47.085 -70.205 -46.755 -69.875 ;
        RECT -47.085 -71.565 -46.755 -71.235 ;
        RECT -47.085 -72.925 -46.755 -72.595 ;
        RECT -47.085 -74.285 -46.755 -73.955 ;
        RECT -47.085 -75.645 -46.755 -75.315 ;
        RECT -47.085 -77.005 -46.755 -76.675 ;
        RECT -47.085 -78.365 -46.755 -78.035 ;
        RECT -47.085 -79.725 -46.755 -79.395 ;
        RECT -47.085 -81.085 -46.755 -80.755 ;
        RECT -47.085 -82.445 -46.755 -82.115 ;
        RECT -47.085 -83.805 -46.755 -83.475 ;
        RECT -47.085 -85.165 -46.755 -84.835 ;
        RECT -47.085 -86.525 -46.755 -86.195 ;
        RECT -47.085 -87.885 -46.755 -87.555 ;
        RECT -47.085 -89.245 -46.755 -88.915 ;
        RECT -47.085 -90.81 -46.755 -90.48 ;
        RECT -47.085 -91.965 -46.755 -91.635 ;
        RECT -47.085 -93.325 -46.755 -92.995 ;
        RECT -47.085 -94.685 -46.755 -94.355 ;
        RECT -47.085 -96.045 -46.755 -95.715 ;
        RECT -47.085 -97.405 -46.755 -97.075 ;
        RECT -47.085 -100.125 -46.755 -99.795 ;
        RECT -47.085 -101.35 -46.755 -101.02 ;
        RECT -47.085 -102.845 -46.755 -102.515 ;
        RECT -47.085 -104.205 -46.755 -103.875 ;
        RECT -47.085 -105.565 -46.755 -105.235 ;
        RECT -47.085 -108.285 -46.755 -107.955 ;
        RECT -47.085 -109.645 -46.755 -109.315 ;
        RECT -47.085 -112.365 -46.755 -112.035 ;
        RECT -47.085 -115.085 -46.755 -114.755 ;
        RECT -47.085 -116.445 -46.755 -116.115 ;
        RECT -47.085 -117.805 -46.755 -117.475 ;
        RECT -47.085 -119.165 -46.755 -118.835 ;
        RECT -47.085 -120.525 -46.755 -120.195 ;
        RECT -47.085 -121.885 -46.755 -121.555 ;
        RECT -47.085 -123.245 -46.755 -122.915 ;
        RECT -47.085 -124.605 -46.755 -124.275 ;
        RECT -47.085 -125.965 -46.755 -125.635 ;
        RECT -47.085 -127.325 -46.755 -126.995 ;
        RECT -47.085 -128.685 -46.755 -128.355 ;
        RECT -47.085 -130.045 -46.755 -129.715 ;
        RECT -47.085 -131.405 -46.755 -131.075 ;
        RECT -47.085 -132.765 -46.755 -132.435 ;
        RECT -47.085 -134.125 -46.755 -133.795 ;
        RECT -47.085 -135.485 -46.755 -135.155 ;
        RECT -47.085 -136.845 -46.755 -136.515 ;
        RECT -47.085 -138.205 -46.755 -137.875 ;
        RECT -47.085 -139.565 -46.755 -139.235 ;
        RECT -47.085 -140.925 -46.755 -140.595 ;
        RECT -47.085 -142.285 -46.755 -141.955 ;
        RECT -47.085 -143.645 -46.755 -143.315 ;
        RECT -47.085 -145.005 -46.755 -144.675 ;
        RECT -47.085 -146.365 -46.755 -146.035 ;
        RECT -47.085 -147.725 -46.755 -147.395 ;
        RECT -47.085 -149.085 -46.755 -148.755 ;
        RECT -47.085 -150.445 -46.755 -150.115 ;
        RECT -47.085 -151.805 -46.755 -151.475 ;
        RECT -47.085 -153.165 -46.755 -152.835 ;
        RECT -47.085 -154.525 -46.755 -154.195 ;
        RECT -47.085 -155.885 -46.755 -155.555 ;
        RECT -47.085 -157.245 -46.755 -156.915 ;
        RECT -47.085 -158.605 -46.755 -158.275 ;
        RECT -47.085 -159.965 -46.755 -159.635 ;
        RECT -47.085 -161.325 -46.755 -160.995 ;
        RECT -47.085 -162.685 -46.755 -162.355 ;
        RECT -47.085 -164.045 -46.755 -163.715 ;
        RECT -47.085 -165.405 -46.755 -165.075 ;
        RECT -47.085 -166.765 -46.755 -166.435 ;
        RECT -47.085 -169.485 -46.755 -169.155 ;
        RECT -47.085 -170.845 -46.755 -170.515 ;
        RECT -47.085 -173.565 -46.755 -173.235 ;
        RECT -47.085 -174.925 -46.755 -174.595 ;
        RECT -47.085 -177.645 -46.755 -177.315 ;
        RECT -47.085 -183.29 -46.755 -182.16 ;
        RECT -47.08 -183.405 -46.76 -29.76 ;
        RECT -47.085 -32.125 -46.755 -31.795 ;
        RECT -47.085 -33.71 -46.755 -33.38 ;
        RECT -47.085 -34.845 -46.755 -34.515 ;
        RECT -47.085 -36.205 -46.755 -35.875 ;
        RECT -47.085 -38.925 -46.755 -38.595 ;
        RECT -47.085 -39.75 -46.755 -39.42 ;
        RECT -47.085 -41.645 -46.755 -41.315 ;
        RECT -47.085 -44.365 -46.755 -44.035 ;
        RECT -47.085 -49.805 -46.755 -49.475 ;
        RECT -47.085 -51.165 -46.755 -50.835 ;
        RECT -47.085 -53.885 -46.755 -53.555 ;
        RECT -47.085 -55.245 -46.755 -54.915 ;
    END
    PORT
      LAYER met3 ;
        RECT -56.605 244.04 -56.275 245.17 ;
        RECT -56.605 239.875 -56.275 240.205 ;
        RECT -56.605 238.515 -56.275 238.845 ;
        RECT -56.605 237.155 -56.275 237.485 ;
        RECT -56.605 235.795 -56.275 236.125 ;
        RECT -56.605 234.435 -56.275 234.765 ;
        RECT -56.605 233.075 -56.275 233.405 ;
        RECT -56.605 231.715 -56.275 232.045 ;
        RECT -56.605 230.355 -56.275 230.685 ;
        RECT -56.605 228.995 -56.275 229.325 ;
        RECT -56.605 227.635 -56.275 227.965 ;
        RECT -56.605 226.275 -56.275 226.605 ;
        RECT -56.605 224.915 -56.275 225.245 ;
        RECT -56.605 223.555 -56.275 223.885 ;
        RECT -56.605 222.195 -56.275 222.525 ;
        RECT -56.605 220.835 -56.275 221.165 ;
        RECT -56.605 219.475 -56.275 219.805 ;
        RECT -56.605 218.115 -56.275 218.445 ;
        RECT -56.605 216.755 -56.275 217.085 ;
        RECT -56.605 215.395 -56.275 215.725 ;
        RECT -56.605 214.035 -56.275 214.365 ;
        RECT -56.605 212.675 -56.275 213.005 ;
        RECT -56.605 211.315 -56.275 211.645 ;
        RECT -56.605 209.955 -56.275 210.285 ;
        RECT -56.605 208.595 -56.275 208.925 ;
        RECT -56.605 207.235 -56.275 207.565 ;
        RECT -56.605 205.875 -56.275 206.205 ;
        RECT -56.605 204.515 -56.275 204.845 ;
        RECT -56.605 203.155 -56.275 203.485 ;
        RECT -56.605 201.795 -56.275 202.125 ;
        RECT -56.605 200.435 -56.275 200.765 ;
        RECT -56.605 199.075 -56.275 199.405 ;
        RECT -56.605 197.715 -56.275 198.045 ;
        RECT -56.605 196.355 -56.275 196.685 ;
        RECT -56.605 194.995 -56.275 195.325 ;
        RECT -56.605 193.635 -56.275 193.965 ;
        RECT -56.605 192.275 -56.275 192.605 ;
        RECT -56.605 190.915 -56.275 191.245 ;
        RECT -56.605 189.555 -56.275 189.885 ;
        RECT -56.605 188.195 -56.275 188.525 ;
        RECT -56.605 186.835 -56.275 187.165 ;
        RECT -56.605 185.475 -56.275 185.805 ;
        RECT -56.605 184.115 -56.275 184.445 ;
        RECT -56.605 182.755 -56.275 183.085 ;
        RECT -56.605 181.395 -56.275 181.725 ;
        RECT -56.605 180.035 -56.275 180.365 ;
        RECT -56.605 178.675 -56.275 179.005 ;
        RECT -56.605 177.315 -56.275 177.645 ;
        RECT -56.605 175.955 -56.275 176.285 ;
        RECT -56.605 174.595 -56.275 174.925 ;
        RECT -56.605 173.235 -56.275 173.565 ;
        RECT -56.605 171.875 -56.275 172.205 ;
        RECT -56.605 170.515 -56.275 170.845 ;
        RECT -56.605 169.155 -56.275 169.485 ;
        RECT -56.605 167.795 -56.275 168.125 ;
        RECT -56.605 166.435 -56.275 166.765 ;
        RECT -56.605 165.075 -56.275 165.405 ;
        RECT -56.605 163.715 -56.275 164.045 ;
        RECT -56.605 162.355 -56.275 162.685 ;
        RECT -56.605 160.995 -56.275 161.325 ;
        RECT -56.605 159.635 -56.275 159.965 ;
        RECT -56.605 158.275 -56.275 158.605 ;
        RECT -56.605 156.915 -56.275 157.245 ;
        RECT -56.605 155.555 -56.275 155.885 ;
        RECT -56.605 154.195 -56.275 154.525 ;
        RECT -56.605 152.835 -56.275 153.165 ;
        RECT -56.605 151.475 -56.275 151.805 ;
        RECT -56.605 150.115 -56.275 150.445 ;
        RECT -56.605 148.755 -56.275 149.085 ;
        RECT -56.605 147.395 -56.275 147.725 ;
        RECT -56.605 146.035 -56.275 146.365 ;
        RECT -56.605 144.675 -56.275 145.005 ;
        RECT -56.605 143.315 -56.275 143.645 ;
        RECT -56.605 141.955 -56.275 142.285 ;
        RECT -56.605 140.595 -56.275 140.925 ;
        RECT -56.605 139.235 -56.275 139.565 ;
        RECT -56.6 138.56 -56.28 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -56.605 97.075 -56.275 97.405 ;
        RECT -56.605 95.715 -56.275 96.045 ;
        RECT -56.605 94.355 -56.275 94.685 ;
        RECT -56.605 92.995 -56.275 93.325 ;
        RECT -56.605 88.915 -56.275 89.245 ;
        RECT -56.605 84.835 -56.275 85.165 ;
        RECT -56.605 83.475 -56.275 83.805 ;
        RECT -56.605 82.115 -56.275 82.445 ;
        RECT -56.605 80.755 -56.275 81.085 ;
        RECT -56.605 79.395 -56.275 79.725 ;
        RECT -56.605 78.035 -56.275 78.365 ;
        RECT -56.605 76.675 -56.275 77.005 ;
        RECT -56.605 75.315 -56.275 75.645 ;
        RECT -56.605 73.955 -56.275 74.285 ;
        RECT -56.605 72.595 -56.275 72.925 ;
        RECT -56.605 71.235 -56.275 71.565 ;
        RECT -56.605 69.875 -56.275 70.205 ;
        RECT -56.605 68.515 -56.275 68.845 ;
        RECT -56.605 67.155 -56.275 67.485 ;
        RECT -56.605 65.795 -56.275 66.125 ;
        RECT -56.605 64.435 -56.275 64.765 ;
        RECT -56.605 63.075 -56.275 63.405 ;
        RECT -56.605 61.715 -56.275 62.045 ;
        RECT -56.605 60.355 -56.275 60.685 ;
        RECT -56.605 58.995 -56.275 59.325 ;
        RECT -56.605 57.635 -56.275 57.965 ;
        RECT -56.605 56.275 -56.275 56.605 ;
        RECT -56.605 54.915 -56.275 55.245 ;
        RECT -56.605 53.555 -56.275 53.885 ;
        RECT -56.605 52.195 -56.275 52.525 ;
        RECT -56.605 50.835 -56.275 51.165 ;
        RECT -56.605 49.475 -56.275 49.805 ;
        RECT -56.605 48.115 -56.275 48.445 ;
        RECT -56.605 46.755 -56.275 47.085 ;
        RECT -56.605 45.395 -56.275 45.725 ;
        RECT -56.605 44.035 -56.275 44.365 ;
        RECT -56.605 42.675 -56.275 43.005 ;
        RECT -56.605 41.315 -56.275 41.645 ;
        RECT -56.605 39.955 -56.275 40.285 ;
        RECT -56.605 38.595 -56.275 38.925 ;
        RECT -56.605 37.235 -56.275 37.565 ;
        RECT -56.605 35.875 -56.275 36.205 ;
        RECT -56.605 34.515 -56.275 34.845 ;
        RECT -56.605 33.155 -56.275 33.485 ;
        RECT -56.605 31.795 -56.275 32.125 ;
        RECT -56.605 30.435 -56.275 30.765 ;
        RECT -56.605 29.075 -56.275 29.405 ;
        RECT -56.605 27.715 -56.275 28.045 ;
        RECT -56.605 26.355 -56.275 26.685 ;
        RECT -56.605 24.995 -56.275 25.325 ;
        RECT -56.605 23.635 -56.275 23.965 ;
        RECT -56.605 22.275 -56.275 22.605 ;
        RECT -56.605 20.915 -56.275 21.245 ;
        RECT -56.605 19.555 -56.275 19.885 ;
        RECT -56.605 18.195 -56.275 18.525 ;
        RECT -56.605 16.835 -56.275 17.165 ;
        RECT -56.605 15.475 -56.275 15.805 ;
        RECT -56.605 14.115 -56.275 14.445 ;
        RECT -56.605 12.755 -56.275 13.085 ;
        RECT -56.605 11.395 -56.275 11.725 ;
        RECT -56.605 10.035 -56.275 10.365 ;
        RECT -56.605 8.675 -56.275 9.005 ;
        RECT -56.605 7.315 -56.275 7.645 ;
        RECT -56.605 5.955 -56.275 6.285 ;
        RECT -56.605 4.595 -56.275 4.925 ;
        RECT -56.605 3.235 -56.275 3.565 ;
        RECT -56.605 1.875 -56.275 2.205 ;
        RECT -56.605 0.515 -56.275 0.845 ;
        RECT -56.605 -0.845 -56.275 -0.515 ;
        RECT -56.605 -2.205 -56.275 -1.875 ;
        RECT -56.605 -3.565 -56.275 -3.235 ;
        RECT -56.605 -4.925 -56.275 -4.595 ;
        RECT -56.605 -6.285 -56.275 -5.955 ;
        RECT -56.605 -7.645 -56.275 -7.315 ;
        RECT -56.605 -9.005 -56.275 -8.675 ;
        RECT -56.605 -10.365 -56.275 -10.035 ;
        RECT -56.605 -11.725 -56.275 -11.395 ;
        RECT -56.605 -13.085 -56.275 -12.755 ;
        RECT -56.605 -14.445 -56.275 -14.115 ;
        RECT -56.605 -15.805 -56.275 -15.475 ;
        RECT -56.605 -17.165 -56.275 -16.835 ;
        RECT -56.605 -18.525 -56.275 -18.195 ;
        RECT -56.605 -19.885 -56.275 -19.555 ;
        RECT -56.605 -21.245 -56.275 -20.915 ;
        RECT -56.605 -22.605 -56.275 -22.275 ;
        RECT -56.605 -23.965 -56.275 -23.635 ;
        RECT -56.605 -25.325 -56.275 -24.995 ;
        RECT -56.605 -28.045 -56.275 -27.715 ;
        RECT -56.605 -29.405 -56.275 -29.075 ;
        RECT -56.605 -30.765 -56.275 -30.435 ;
        RECT -56.605 -32.125 -56.275 -31.795 ;
        RECT -56.605 -33.485 -56.275 -33.155 ;
        RECT -56.605 -34.845 -56.275 -34.515 ;
        RECT -56.605 -36.205 -56.275 -35.875 ;
        RECT -56.605 -37.565 -56.275 -37.235 ;
        RECT -56.605 -38.925 -56.275 -38.595 ;
        RECT -56.605 -40.285 -56.275 -39.955 ;
        RECT -56.605 -41.645 -56.275 -41.315 ;
        RECT -56.605 -43.005 -56.275 -42.675 ;
        RECT -56.605 -44.365 -56.275 -44.035 ;
        RECT -56.605 -45.725 -56.275 -45.395 ;
        RECT -56.605 -47.085 -56.275 -46.755 ;
        RECT -56.605 -48.445 -56.275 -48.115 ;
        RECT -56.605 -49.805 -56.275 -49.475 ;
        RECT -56.605 -51.165 -56.275 -50.835 ;
        RECT -56.605 -52.525 -56.275 -52.195 ;
        RECT -56.605 -53.885 -56.275 -53.555 ;
        RECT -56.605 -55.245 -56.275 -54.915 ;
        RECT -56.605 -56.605 -56.275 -56.275 ;
        RECT -56.605 -57.965 -56.275 -57.635 ;
        RECT -56.605 -59.325 -56.275 -58.995 ;
        RECT -56.605 -60.685 -56.275 -60.355 ;
        RECT -56.605 -62.045 -56.275 -61.715 ;
        RECT -56.605 -63.405 -56.275 -63.075 ;
        RECT -56.605 -64.765 -56.275 -64.435 ;
        RECT -56.605 -66.125 -56.275 -65.795 ;
        RECT -56.605 -67.485 -56.275 -67.155 ;
        RECT -56.605 -68.845 -56.275 -68.515 ;
        RECT -56.605 -70.205 -56.275 -69.875 ;
        RECT -56.605 -71.565 -56.275 -71.235 ;
        RECT -56.605 -72.925 -56.275 -72.595 ;
        RECT -56.605 -74.285 -56.275 -73.955 ;
        RECT -56.605 -75.645 -56.275 -75.315 ;
        RECT -56.605 -77.005 -56.275 -76.675 ;
        RECT -56.605 -78.365 -56.275 -78.035 ;
        RECT -56.605 -79.725 -56.275 -79.395 ;
        RECT -56.605 -81.085 -56.275 -80.755 ;
        RECT -56.605 -82.445 -56.275 -82.115 ;
        RECT -56.605 -83.805 -56.275 -83.475 ;
        RECT -56.605 -85.165 -56.275 -84.835 ;
        RECT -56.605 -86.525 -56.275 -86.195 ;
        RECT -56.605 -87.885 -56.275 -87.555 ;
        RECT -56.605 -89.245 -56.275 -88.915 ;
        RECT -56.605 -90.81 -56.275 -90.48 ;
        RECT -56.605 -91.965 -56.275 -91.635 ;
        RECT -56.605 -93.325 -56.275 -92.995 ;
        RECT -56.605 -94.685 -56.275 -94.355 ;
        RECT -56.605 -96.045 -56.275 -95.715 ;
        RECT -56.605 -97.405 -56.275 -97.075 ;
        RECT -56.605 -100.125 -56.275 -99.795 ;
        RECT -56.605 -101.35 -56.275 -101.02 ;
        RECT -56.605 -102.845 -56.275 -102.515 ;
        RECT -56.605 -104.205 -56.275 -103.875 ;
        RECT -56.605 -105.565 -56.275 -105.235 ;
        RECT -56.605 -108.285 -56.275 -107.955 ;
        RECT -56.605 -109.645 -56.275 -109.315 ;
        RECT -56.605 -112.365 -56.275 -112.035 ;
        RECT -56.605 -115.085 -56.275 -114.755 ;
        RECT -56.605 -116.445 -56.275 -116.115 ;
        RECT -56.605 -117.805 -56.275 -117.475 ;
        RECT -56.605 -119.165 -56.275 -118.835 ;
        RECT -56.605 -120.525 -56.275 -120.195 ;
        RECT -56.605 -121.885 -56.275 -121.555 ;
        RECT -56.605 -123.245 -56.275 -122.915 ;
        RECT -56.605 -124.605 -56.275 -124.275 ;
        RECT -56.605 -125.965 -56.275 -125.635 ;
        RECT -56.605 -127.325 -56.275 -126.995 ;
        RECT -56.605 -128.685 -56.275 -128.355 ;
        RECT -56.605 -130.045 -56.275 -129.715 ;
        RECT -56.605 -131.405 -56.275 -131.075 ;
        RECT -56.605 -132.765 -56.275 -132.435 ;
        RECT -56.605 -134.125 -56.275 -133.795 ;
        RECT -56.605 -135.485 -56.275 -135.155 ;
        RECT -56.605 -136.845 -56.275 -136.515 ;
        RECT -56.605 -138.205 -56.275 -137.875 ;
        RECT -56.605 -139.565 -56.275 -139.235 ;
        RECT -56.605 -140.925 -56.275 -140.595 ;
        RECT -56.605 -142.285 -56.275 -141.955 ;
        RECT -56.605 -143.645 -56.275 -143.315 ;
        RECT -56.605 -145.005 -56.275 -144.675 ;
        RECT -56.605 -146.365 -56.275 -146.035 ;
        RECT -56.605 -147.725 -56.275 -147.395 ;
        RECT -56.605 -149.085 -56.275 -148.755 ;
        RECT -56.605 -150.445 -56.275 -150.115 ;
        RECT -56.605 -151.805 -56.275 -151.475 ;
        RECT -56.605 -153.165 -56.275 -152.835 ;
        RECT -56.605 -154.525 -56.275 -154.195 ;
        RECT -56.605 -155.885 -56.275 -155.555 ;
        RECT -56.605 -157.245 -56.275 -156.915 ;
        RECT -56.605 -158.605 -56.275 -158.275 ;
        RECT -56.605 -159.965 -56.275 -159.635 ;
        RECT -56.605 -161.325 -56.275 -160.995 ;
        RECT -56.605 -162.685 -56.275 -162.355 ;
        RECT -56.605 -164.045 -56.275 -163.715 ;
        RECT -56.605 -165.405 -56.275 -165.075 ;
        RECT -56.605 -166.765 -56.275 -166.435 ;
        RECT -56.605 -168.655 -56.275 -168.325 ;
        RECT -56.605 -169.485 -56.275 -169.155 ;
        RECT -56.605 -170.845 -56.275 -170.515 ;
        RECT -56.605 -172.205 -56.275 -171.875 ;
        RECT -56.605 -173.565 -56.275 -173.235 ;
        RECT -56.605 -174.925 -56.275 -174.595 ;
        RECT -56.605 -177.645 -56.275 -177.315 ;
        RECT -56.605 -183.29 -56.275 -182.16 ;
        RECT -56.6 -183.405 -56.28 98.08 ;
    END
    PORT
      LAYER met3 ;
        RECT -55.245 244.04 -54.915 245.17 ;
        RECT -55.245 239.875 -54.915 240.205 ;
        RECT -55.245 238.515 -54.915 238.845 ;
        RECT -55.245 237.155 -54.915 237.485 ;
        RECT -55.245 235.795 -54.915 236.125 ;
        RECT -55.245 234.435 -54.915 234.765 ;
        RECT -55.245 233.075 -54.915 233.405 ;
        RECT -55.245 231.715 -54.915 232.045 ;
        RECT -55.245 230.355 -54.915 230.685 ;
        RECT -55.245 228.995 -54.915 229.325 ;
        RECT -55.245 227.635 -54.915 227.965 ;
        RECT -55.245 226.275 -54.915 226.605 ;
        RECT -55.245 224.915 -54.915 225.245 ;
        RECT -55.245 223.555 -54.915 223.885 ;
        RECT -55.245 222.195 -54.915 222.525 ;
        RECT -55.245 220.835 -54.915 221.165 ;
        RECT -55.245 219.475 -54.915 219.805 ;
        RECT -55.245 218.115 -54.915 218.445 ;
        RECT -55.245 216.755 -54.915 217.085 ;
        RECT -55.245 215.395 -54.915 215.725 ;
        RECT -55.245 214.035 -54.915 214.365 ;
        RECT -55.245 212.675 -54.915 213.005 ;
        RECT -55.245 211.315 -54.915 211.645 ;
        RECT -55.245 209.955 -54.915 210.285 ;
        RECT -55.245 208.595 -54.915 208.925 ;
        RECT -55.245 207.235 -54.915 207.565 ;
        RECT -55.245 205.875 -54.915 206.205 ;
        RECT -55.245 204.515 -54.915 204.845 ;
        RECT -55.245 203.155 -54.915 203.485 ;
        RECT -55.245 201.795 -54.915 202.125 ;
        RECT -55.245 200.435 -54.915 200.765 ;
        RECT -55.245 199.075 -54.915 199.405 ;
        RECT -55.245 197.715 -54.915 198.045 ;
        RECT -55.245 196.355 -54.915 196.685 ;
        RECT -55.245 194.995 -54.915 195.325 ;
        RECT -55.245 193.635 -54.915 193.965 ;
        RECT -55.245 192.275 -54.915 192.605 ;
        RECT -55.245 190.915 -54.915 191.245 ;
        RECT -55.245 189.555 -54.915 189.885 ;
        RECT -55.245 188.195 -54.915 188.525 ;
        RECT -55.245 186.835 -54.915 187.165 ;
        RECT -55.245 185.475 -54.915 185.805 ;
        RECT -55.245 184.115 -54.915 184.445 ;
        RECT -55.245 182.755 -54.915 183.085 ;
        RECT -55.245 181.395 -54.915 181.725 ;
        RECT -55.245 180.035 -54.915 180.365 ;
        RECT -55.245 178.675 -54.915 179.005 ;
        RECT -55.245 177.315 -54.915 177.645 ;
        RECT -55.245 175.955 -54.915 176.285 ;
        RECT -55.245 174.595 -54.915 174.925 ;
        RECT -55.245 173.235 -54.915 173.565 ;
        RECT -55.245 171.875 -54.915 172.205 ;
        RECT -55.245 170.515 -54.915 170.845 ;
        RECT -55.245 169.155 -54.915 169.485 ;
        RECT -55.245 167.795 -54.915 168.125 ;
        RECT -55.245 166.435 -54.915 166.765 ;
        RECT -55.245 165.075 -54.915 165.405 ;
        RECT -55.245 163.715 -54.915 164.045 ;
        RECT -55.245 162.355 -54.915 162.685 ;
        RECT -55.245 160.995 -54.915 161.325 ;
        RECT -55.245 159.635 -54.915 159.965 ;
        RECT -55.245 158.275 -54.915 158.605 ;
        RECT -55.245 156.915 -54.915 157.245 ;
        RECT -55.245 155.555 -54.915 155.885 ;
        RECT -55.245 154.195 -54.915 154.525 ;
        RECT -55.245 152.835 -54.915 153.165 ;
        RECT -55.245 151.475 -54.915 151.805 ;
        RECT -55.245 150.115 -54.915 150.445 ;
        RECT -55.245 148.755 -54.915 149.085 ;
        RECT -55.245 147.395 -54.915 147.725 ;
        RECT -55.245 146.035 -54.915 146.365 ;
        RECT -55.245 144.675 -54.915 145.005 ;
        RECT -55.245 143.315 -54.915 143.645 ;
        RECT -55.245 141.955 -54.915 142.285 ;
        RECT -55.245 140.595 -54.915 140.925 ;
        RECT -55.245 139.235 -54.915 139.565 ;
        RECT -55.24 138.56 -54.92 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -55.245 97.075 -54.915 97.405 ;
        RECT -55.245 95.715 -54.915 96.045 ;
        RECT -55.245 94.355 -54.915 94.685 ;
        RECT -55.245 92.995 -54.915 93.325 ;
        RECT -55.245 88.915 -54.915 89.245 ;
        RECT -55.245 84.835 -54.915 85.165 ;
        RECT -55.245 83.475 -54.915 83.805 ;
        RECT -55.245 82.115 -54.915 82.445 ;
        RECT -55.245 80.755 -54.915 81.085 ;
        RECT -55.245 79.395 -54.915 79.725 ;
        RECT -55.245 78.035 -54.915 78.365 ;
        RECT -55.245 76.675 -54.915 77.005 ;
        RECT -55.245 75.315 -54.915 75.645 ;
        RECT -55.245 73.955 -54.915 74.285 ;
        RECT -55.245 72.595 -54.915 72.925 ;
        RECT -55.245 71.235 -54.915 71.565 ;
        RECT -55.245 69.875 -54.915 70.205 ;
        RECT -55.245 68.515 -54.915 68.845 ;
        RECT -55.245 67.155 -54.915 67.485 ;
        RECT -55.245 65.795 -54.915 66.125 ;
        RECT -55.245 64.435 -54.915 64.765 ;
        RECT -55.245 63.075 -54.915 63.405 ;
        RECT -55.245 61.715 -54.915 62.045 ;
        RECT -55.245 60.355 -54.915 60.685 ;
        RECT -55.245 58.995 -54.915 59.325 ;
        RECT -55.245 57.635 -54.915 57.965 ;
        RECT -55.245 56.275 -54.915 56.605 ;
        RECT -55.245 54.915 -54.915 55.245 ;
        RECT -55.245 53.555 -54.915 53.885 ;
        RECT -55.245 52.195 -54.915 52.525 ;
        RECT -55.245 50.835 -54.915 51.165 ;
        RECT -55.245 49.475 -54.915 49.805 ;
        RECT -55.245 48.115 -54.915 48.445 ;
        RECT -55.245 46.755 -54.915 47.085 ;
        RECT -55.245 45.395 -54.915 45.725 ;
        RECT -55.245 44.035 -54.915 44.365 ;
        RECT -55.245 42.675 -54.915 43.005 ;
        RECT -55.245 41.315 -54.915 41.645 ;
        RECT -55.245 39.955 -54.915 40.285 ;
        RECT -55.245 38.595 -54.915 38.925 ;
        RECT -55.245 37.235 -54.915 37.565 ;
        RECT -55.245 35.875 -54.915 36.205 ;
        RECT -55.245 34.515 -54.915 34.845 ;
        RECT -55.245 33.155 -54.915 33.485 ;
        RECT -55.245 31.795 -54.915 32.125 ;
        RECT -55.245 30.435 -54.915 30.765 ;
        RECT -55.245 29.075 -54.915 29.405 ;
        RECT -55.245 27.715 -54.915 28.045 ;
        RECT -55.245 26.355 -54.915 26.685 ;
        RECT -55.245 24.995 -54.915 25.325 ;
        RECT -55.245 23.635 -54.915 23.965 ;
        RECT -55.245 22.275 -54.915 22.605 ;
        RECT -55.245 20.915 -54.915 21.245 ;
        RECT -55.245 19.555 -54.915 19.885 ;
        RECT -55.245 18.195 -54.915 18.525 ;
        RECT -55.245 16.835 -54.915 17.165 ;
        RECT -55.245 15.475 -54.915 15.805 ;
        RECT -55.245 14.115 -54.915 14.445 ;
        RECT -55.245 12.755 -54.915 13.085 ;
        RECT -55.245 11.395 -54.915 11.725 ;
        RECT -55.245 10.035 -54.915 10.365 ;
        RECT -55.245 8.675 -54.915 9.005 ;
        RECT -55.245 7.315 -54.915 7.645 ;
        RECT -55.245 5.955 -54.915 6.285 ;
        RECT -55.245 4.595 -54.915 4.925 ;
        RECT -55.245 3.235 -54.915 3.565 ;
        RECT -55.245 1.875 -54.915 2.205 ;
        RECT -55.245 0.515 -54.915 0.845 ;
        RECT -55.245 -0.845 -54.915 -0.515 ;
        RECT -55.245 -2.205 -54.915 -1.875 ;
        RECT -55.245 -3.565 -54.915 -3.235 ;
        RECT -55.245 -4.925 -54.915 -4.595 ;
        RECT -55.245 -6.285 -54.915 -5.955 ;
        RECT -55.245 -7.645 -54.915 -7.315 ;
        RECT -55.245 -9.005 -54.915 -8.675 ;
        RECT -55.245 -10.365 -54.915 -10.035 ;
        RECT -55.245 -11.725 -54.915 -11.395 ;
        RECT -55.245 -13.085 -54.915 -12.755 ;
        RECT -55.245 -14.445 -54.915 -14.115 ;
        RECT -55.245 -15.805 -54.915 -15.475 ;
        RECT -55.245 -17.165 -54.915 -16.835 ;
        RECT -55.245 -18.525 -54.915 -18.195 ;
        RECT -55.245 -19.885 -54.915 -19.555 ;
        RECT -55.245 -21.245 -54.915 -20.915 ;
        RECT -55.245 -22.605 -54.915 -22.275 ;
        RECT -55.245 -23.965 -54.915 -23.635 ;
        RECT -55.245 -25.325 -54.915 -24.995 ;
        RECT -55.245 -28.045 -54.915 -27.715 ;
        RECT -55.245 -29.405 -54.915 -29.075 ;
        RECT -55.245 -30.765 -54.915 -30.435 ;
        RECT -55.245 -32.125 -54.915 -31.795 ;
        RECT -55.245 -33.485 -54.915 -33.155 ;
        RECT -55.245 -34.845 -54.915 -34.515 ;
        RECT -55.245 -36.205 -54.915 -35.875 ;
        RECT -55.245 -37.565 -54.915 -37.235 ;
        RECT -55.245 -38.925 -54.915 -38.595 ;
        RECT -55.245 -40.285 -54.915 -39.955 ;
        RECT -55.245 -41.645 -54.915 -41.315 ;
        RECT -55.245 -43.005 -54.915 -42.675 ;
        RECT -55.245 -44.365 -54.915 -44.035 ;
        RECT -55.245 -45.725 -54.915 -45.395 ;
        RECT -55.245 -47.085 -54.915 -46.755 ;
        RECT -55.245 -48.445 -54.915 -48.115 ;
        RECT -55.245 -49.805 -54.915 -49.475 ;
        RECT -55.245 -51.165 -54.915 -50.835 ;
        RECT -55.245 -52.525 -54.915 -52.195 ;
        RECT -55.245 -53.885 -54.915 -53.555 ;
        RECT -55.245 -55.245 -54.915 -54.915 ;
        RECT -55.245 -56.605 -54.915 -56.275 ;
        RECT -55.245 -57.965 -54.915 -57.635 ;
        RECT -55.245 -59.325 -54.915 -58.995 ;
        RECT -55.245 -60.685 -54.915 -60.355 ;
        RECT -55.245 -62.045 -54.915 -61.715 ;
        RECT -55.245 -63.405 -54.915 -63.075 ;
        RECT -55.245 -64.765 -54.915 -64.435 ;
        RECT -55.245 -66.125 -54.915 -65.795 ;
        RECT -55.245 -67.485 -54.915 -67.155 ;
        RECT -55.245 -68.845 -54.915 -68.515 ;
        RECT -55.245 -70.205 -54.915 -69.875 ;
        RECT -55.245 -71.565 -54.915 -71.235 ;
        RECT -55.245 -72.925 -54.915 -72.595 ;
        RECT -55.245 -74.285 -54.915 -73.955 ;
        RECT -55.245 -75.645 -54.915 -75.315 ;
        RECT -55.245 -77.005 -54.915 -76.675 ;
        RECT -55.245 -78.365 -54.915 -78.035 ;
        RECT -55.245 -79.725 -54.915 -79.395 ;
        RECT -55.245 -81.085 -54.915 -80.755 ;
        RECT -55.245 -82.445 -54.915 -82.115 ;
        RECT -55.245 -83.805 -54.915 -83.475 ;
        RECT -55.245 -85.165 -54.915 -84.835 ;
        RECT -55.245 -86.525 -54.915 -86.195 ;
        RECT -55.245 -87.885 -54.915 -87.555 ;
        RECT -55.245 -89.245 -54.915 -88.915 ;
        RECT -55.245 -90.81 -54.915 -90.48 ;
        RECT -55.245 -91.965 -54.915 -91.635 ;
        RECT -55.245 -93.325 -54.915 -92.995 ;
        RECT -55.245 -94.685 -54.915 -94.355 ;
        RECT -55.245 -96.045 -54.915 -95.715 ;
        RECT -55.245 -97.405 -54.915 -97.075 ;
        RECT -55.245 -100.125 -54.915 -99.795 ;
        RECT -55.245 -101.35 -54.915 -101.02 ;
        RECT -55.245 -102.845 -54.915 -102.515 ;
        RECT -55.245 -104.205 -54.915 -103.875 ;
        RECT -55.245 -105.565 -54.915 -105.235 ;
        RECT -55.245 -108.285 -54.915 -107.955 ;
        RECT -55.245 -109.645 -54.915 -109.315 ;
        RECT -55.245 -112.365 -54.915 -112.035 ;
        RECT -55.245 -115.085 -54.915 -114.755 ;
        RECT -55.245 -116.445 -54.915 -116.115 ;
        RECT -55.245 -117.805 -54.915 -117.475 ;
        RECT -55.245 -119.165 -54.915 -118.835 ;
        RECT -55.245 -120.525 -54.915 -120.195 ;
        RECT -55.245 -121.885 -54.915 -121.555 ;
        RECT -55.245 -123.245 -54.915 -122.915 ;
        RECT -55.245 -124.605 -54.915 -124.275 ;
        RECT -55.245 -125.965 -54.915 -125.635 ;
        RECT -55.245 -127.325 -54.915 -126.995 ;
        RECT -55.245 -128.685 -54.915 -128.355 ;
        RECT -55.245 -130.045 -54.915 -129.715 ;
        RECT -55.245 -131.405 -54.915 -131.075 ;
        RECT -55.245 -132.765 -54.915 -132.435 ;
        RECT -55.245 -134.125 -54.915 -133.795 ;
        RECT -55.245 -135.485 -54.915 -135.155 ;
        RECT -55.245 -136.845 -54.915 -136.515 ;
        RECT -55.245 -138.205 -54.915 -137.875 ;
        RECT -55.245 -139.565 -54.915 -139.235 ;
        RECT -55.245 -140.925 -54.915 -140.595 ;
        RECT -55.245 -142.285 -54.915 -141.955 ;
        RECT -55.245 -143.645 -54.915 -143.315 ;
        RECT -55.245 -145.005 -54.915 -144.675 ;
        RECT -55.245 -146.365 -54.915 -146.035 ;
        RECT -55.245 -147.725 -54.915 -147.395 ;
        RECT -55.245 -149.085 -54.915 -148.755 ;
        RECT -55.245 -150.445 -54.915 -150.115 ;
        RECT -55.245 -151.805 -54.915 -151.475 ;
        RECT -55.245 -153.165 -54.915 -152.835 ;
        RECT -55.245 -154.525 -54.915 -154.195 ;
        RECT -55.245 -155.885 -54.915 -155.555 ;
        RECT -55.245 -157.245 -54.915 -156.915 ;
        RECT -55.245 -158.605 -54.915 -158.275 ;
        RECT -55.245 -159.965 -54.915 -159.635 ;
        RECT -55.245 -161.325 -54.915 -160.995 ;
        RECT -55.245 -162.685 -54.915 -162.355 ;
        RECT -55.245 -164.045 -54.915 -163.715 ;
        RECT -55.245 -165.405 -54.915 -165.075 ;
        RECT -55.245 -166.765 -54.915 -166.435 ;
        RECT -55.245 -168.655 -54.915 -168.325 ;
        RECT -55.245 -169.485 -54.915 -169.155 ;
        RECT -55.245 -170.845 -54.915 -170.515 ;
        RECT -55.245 -172.205 -54.915 -171.875 ;
        RECT -55.245 -173.565 -54.915 -173.235 ;
        RECT -55.245 -174.925 -54.915 -174.595 ;
        RECT -55.245 -177.645 -54.915 -177.315 ;
        RECT -55.245 -183.29 -54.915 -182.16 ;
        RECT -55.24 -183.405 -54.92 98.08 ;
    END
    PORT
      LAYER met3 ;
        RECT -53.885 244.04 -53.555 245.17 ;
        RECT -53.885 239.875 -53.555 240.205 ;
        RECT -53.885 238.515 -53.555 238.845 ;
        RECT -53.885 237.155 -53.555 237.485 ;
        RECT -53.885 235.795 -53.555 236.125 ;
        RECT -53.885 234.435 -53.555 234.765 ;
        RECT -53.885 233.075 -53.555 233.405 ;
        RECT -53.885 231.715 -53.555 232.045 ;
        RECT -53.885 230.355 -53.555 230.685 ;
        RECT -53.885 228.995 -53.555 229.325 ;
        RECT -53.885 227.635 -53.555 227.965 ;
        RECT -53.885 226.275 -53.555 226.605 ;
        RECT -53.885 224.915 -53.555 225.245 ;
        RECT -53.885 223.555 -53.555 223.885 ;
        RECT -53.885 222.195 -53.555 222.525 ;
        RECT -53.885 220.835 -53.555 221.165 ;
        RECT -53.885 219.475 -53.555 219.805 ;
        RECT -53.885 218.115 -53.555 218.445 ;
        RECT -53.885 216.755 -53.555 217.085 ;
        RECT -53.885 215.395 -53.555 215.725 ;
        RECT -53.885 214.035 -53.555 214.365 ;
        RECT -53.885 212.675 -53.555 213.005 ;
        RECT -53.885 211.315 -53.555 211.645 ;
        RECT -53.885 209.955 -53.555 210.285 ;
        RECT -53.885 208.595 -53.555 208.925 ;
        RECT -53.885 207.235 -53.555 207.565 ;
        RECT -53.885 205.875 -53.555 206.205 ;
        RECT -53.885 204.515 -53.555 204.845 ;
        RECT -53.885 203.155 -53.555 203.485 ;
        RECT -53.885 201.795 -53.555 202.125 ;
        RECT -53.885 200.435 -53.555 200.765 ;
        RECT -53.885 199.075 -53.555 199.405 ;
        RECT -53.885 197.715 -53.555 198.045 ;
        RECT -53.885 196.355 -53.555 196.685 ;
        RECT -53.885 194.995 -53.555 195.325 ;
        RECT -53.885 193.635 -53.555 193.965 ;
        RECT -53.885 192.275 -53.555 192.605 ;
        RECT -53.885 190.915 -53.555 191.245 ;
        RECT -53.885 189.555 -53.555 189.885 ;
        RECT -53.885 188.195 -53.555 188.525 ;
        RECT -53.885 186.835 -53.555 187.165 ;
        RECT -53.885 185.475 -53.555 185.805 ;
        RECT -53.885 184.115 -53.555 184.445 ;
        RECT -53.885 182.755 -53.555 183.085 ;
        RECT -53.885 181.395 -53.555 181.725 ;
        RECT -53.885 180.035 -53.555 180.365 ;
        RECT -53.885 178.675 -53.555 179.005 ;
        RECT -53.885 177.315 -53.555 177.645 ;
        RECT -53.885 175.955 -53.555 176.285 ;
        RECT -53.885 174.595 -53.555 174.925 ;
        RECT -53.885 173.235 -53.555 173.565 ;
        RECT -53.885 171.875 -53.555 172.205 ;
        RECT -53.885 170.515 -53.555 170.845 ;
        RECT -53.885 169.155 -53.555 169.485 ;
        RECT -53.885 167.795 -53.555 168.125 ;
        RECT -53.885 166.435 -53.555 166.765 ;
        RECT -53.885 165.075 -53.555 165.405 ;
        RECT -53.885 163.715 -53.555 164.045 ;
        RECT -53.885 162.355 -53.555 162.685 ;
        RECT -53.885 160.995 -53.555 161.325 ;
        RECT -53.885 159.635 -53.555 159.965 ;
        RECT -53.885 158.275 -53.555 158.605 ;
        RECT -53.885 156.915 -53.555 157.245 ;
        RECT -53.885 155.555 -53.555 155.885 ;
        RECT -53.885 154.195 -53.555 154.525 ;
        RECT -53.885 152.835 -53.555 153.165 ;
        RECT -53.885 151.475 -53.555 151.805 ;
        RECT -53.885 150.115 -53.555 150.445 ;
        RECT -53.885 148.755 -53.555 149.085 ;
        RECT -53.885 147.395 -53.555 147.725 ;
        RECT -53.885 146.035 -53.555 146.365 ;
        RECT -53.885 144.675 -53.555 145.005 ;
        RECT -53.885 143.315 -53.555 143.645 ;
        RECT -53.885 141.955 -53.555 142.285 ;
        RECT -53.885 140.595 -53.555 140.925 ;
        RECT -53.885 139.235 -53.555 139.565 ;
        RECT -53.88 138.56 -53.56 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -53.885 97.075 -53.555 97.405 ;
        RECT -53.885 95.715 -53.555 96.045 ;
        RECT -53.885 94.355 -53.555 94.685 ;
        RECT -53.885 92.995 -53.555 93.325 ;
        RECT -53.885 88.915 -53.555 89.245 ;
        RECT -53.885 84.835 -53.555 85.165 ;
        RECT -53.885 83.475 -53.555 83.805 ;
        RECT -53.885 82.115 -53.555 82.445 ;
        RECT -53.885 80.755 -53.555 81.085 ;
        RECT -53.885 79.395 -53.555 79.725 ;
        RECT -53.885 78.035 -53.555 78.365 ;
        RECT -53.885 76.675 -53.555 77.005 ;
        RECT -53.885 75.315 -53.555 75.645 ;
        RECT -53.885 73.955 -53.555 74.285 ;
        RECT -53.885 72.595 -53.555 72.925 ;
        RECT -53.885 71.235 -53.555 71.565 ;
        RECT -53.885 69.875 -53.555 70.205 ;
        RECT -53.885 68.515 -53.555 68.845 ;
        RECT -53.885 67.155 -53.555 67.485 ;
        RECT -53.885 65.795 -53.555 66.125 ;
        RECT -53.885 64.435 -53.555 64.765 ;
        RECT -53.885 63.075 -53.555 63.405 ;
        RECT -53.885 61.715 -53.555 62.045 ;
        RECT -53.885 60.355 -53.555 60.685 ;
        RECT -53.885 58.995 -53.555 59.325 ;
        RECT -53.885 57.635 -53.555 57.965 ;
        RECT -53.885 56.275 -53.555 56.605 ;
        RECT -53.885 54.915 -53.555 55.245 ;
        RECT -53.885 53.555 -53.555 53.885 ;
        RECT -53.885 52.195 -53.555 52.525 ;
        RECT -53.885 50.835 -53.555 51.165 ;
        RECT -53.885 49.475 -53.555 49.805 ;
        RECT -53.885 48.115 -53.555 48.445 ;
        RECT -53.885 46.755 -53.555 47.085 ;
        RECT -53.885 45.395 -53.555 45.725 ;
        RECT -53.885 44.035 -53.555 44.365 ;
        RECT -53.885 42.675 -53.555 43.005 ;
        RECT -53.885 41.315 -53.555 41.645 ;
        RECT -53.885 39.955 -53.555 40.285 ;
        RECT -53.885 38.595 -53.555 38.925 ;
        RECT -53.885 37.235 -53.555 37.565 ;
        RECT -53.885 35.875 -53.555 36.205 ;
        RECT -53.885 34.515 -53.555 34.845 ;
        RECT -53.885 33.155 -53.555 33.485 ;
        RECT -53.885 31.795 -53.555 32.125 ;
        RECT -53.885 30.435 -53.555 30.765 ;
        RECT -53.885 29.075 -53.555 29.405 ;
        RECT -53.885 27.715 -53.555 28.045 ;
        RECT -53.885 26.355 -53.555 26.685 ;
        RECT -53.885 24.995 -53.555 25.325 ;
        RECT -53.885 23.635 -53.555 23.965 ;
        RECT -53.885 22.275 -53.555 22.605 ;
        RECT -53.885 20.915 -53.555 21.245 ;
        RECT -53.885 19.555 -53.555 19.885 ;
        RECT -53.885 18.195 -53.555 18.525 ;
        RECT -53.885 16.835 -53.555 17.165 ;
        RECT -53.885 15.475 -53.555 15.805 ;
        RECT -53.885 14.115 -53.555 14.445 ;
        RECT -53.885 12.755 -53.555 13.085 ;
        RECT -53.885 11.395 -53.555 11.725 ;
        RECT -53.885 10.035 -53.555 10.365 ;
        RECT -53.885 8.675 -53.555 9.005 ;
        RECT -53.885 7.315 -53.555 7.645 ;
        RECT -53.885 5.955 -53.555 6.285 ;
        RECT -53.885 4.595 -53.555 4.925 ;
        RECT -53.885 3.235 -53.555 3.565 ;
        RECT -53.885 1.875 -53.555 2.205 ;
        RECT -53.885 0.515 -53.555 0.845 ;
        RECT -53.885 -0.845 -53.555 -0.515 ;
        RECT -53.885 -2.205 -53.555 -1.875 ;
        RECT -53.885 -3.565 -53.555 -3.235 ;
        RECT -53.885 -4.925 -53.555 -4.595 ;
        RECT -53.885 -6.285 -53.555 -5.955 ;
        RECT -53.885 -7.645 -53.555 -7.315 ;
        RECT -53.885 -9.005 -53.555 -8.675 ;
        RECT -53.885 -10.365 -53.555 -10.035 ;
        RECT -53.885 -11.725 -53.555 -11.395 ;
        RECT -53.885 -13.085 -53.555 -12.755 ;
        RECT -53.885 -14.445 -53.555 -14.115 ;
        RECT -53.885 -15.805 -53.555 -15.475 ;
        RECT -53.885 -17.165 -53.555 -16.835 ;
        RECT -53.885 -18.525 -53.555 -18.195 ;
        RECT -53.885 -19.885 -53.555 -19.555 ;
        RECT -53.885 -21.245 -53.555 -20.915 ;
        RECT -53.885 -22.605 -53.555 -22.275 ;
        RECT -53.885 -23.965 -53.555 -23.635 ;
        RECT -53.885 -25.325 -53.555 -24.995 ;
        RECT -53.885 -28.045 -53.555 -27.715 ;
        RECT -53.885 -29.405 -53.555 -29.075 ;
        RECT -53.885 -30.765 -53.555 -30.435 ;
        RECT -53.885 -32.125 -53.555 -31.795 ;
        RECT -53.885 -33.485 -53.555 -33.155 ;
        RECT -53.885 -34.845 -53.555 -34.515 ;
        RECT -53.885 -36.205 -53.555 -35.875 ;
        RECT -53.885 -37.565 -53.555 -37.235 ;
        RECT -53.885 -38.925 -53.555 -38.595 ;
        RECT -53.885 -40.285 -53.555 -39.955 ;
        RECT -53.885 -41.645 -53.555 -41.315 ;
        RECT -53.885 -43.005 -53.555 -42.675 ;
        RECT -53.885 -44.365 -53.555 -44.035 ;
        RECT -53.885 -45.725 -53.555 -45.395 ;
        RECT -53.885 -47.085 -53.555 -46.755 ;
        RECT -53.885 -48.445 -53.555 -48.115 ;
        RECT -53.885 -49.805 -53.555 -49.475 ;
        RECT -53.885 -51.165 -53.555 -50.835 ;
        RECT -53.885 -52.525 -53.555 -52.195 ;
        RECT -53.885 -53.885 -53.555 -53.555 ;
        RECT -53.885 -55.245 -53.555 -54.915 ;
        RECT -53.885 -56.605 -53.555 -56.275 ;
        RECT -53.885 -57.965 -53.555 -57.635 ;
        RECT -53.885 -59.325 -53.555 -58.995 ;
        RECT -53.885 -60.685 -53.555 -60.355 ;
        RECT -53.885 -62.045 -53.555 -61.715 ;
        RECT -53.885 -63.405 -53.555 -63.075 ;
        RECT -53.885 -64.765 -53.555 -64.435 ;
        RECT -53.885 -66.125 -53.555 -65.795 ;
        RECT -53.885 -67.485 -53.555 -67.155 ;
        RECT -53.885 -68.845 -53.555 -68.515 ;
        RECT -53.885 -70.205 -53.555 -69.875 ;
        RECT -53.885 -71.565 -53.555 -71.235 ;
        RECT -53.885 -72.925 -53.555 -72.595 ;
        RECT -53.885 -74.285 -53.555 -73.955 ;
        RECT -53.885 -75.645 -53.555 -75.315 ;
        RECT -53.885 -77.005 -53.555 -76.675 ;
        RECT -53.885 -78.365 -53.555 -78.035 ;
        RECT -53.885 -79.725 -53.555 -79.395 ;
        RECT -53.885 -81.085 -53.555 -80.755 ;
        RECT -53.885 -82.445 -53.555 -82.115 ;
        RECT -53.885 -83.805 -53.555 -83.475 ;
        RECT -53.885 -85.165 -53.555 -84.835 ;
        RECT -53.885 -86.525 -53.555 -86.195 ;
        RECT -53.885 -87.885 -53.555 -87.555 ;
        RECT -53.885 -89.245 -53.555 -88.915 ;
        RECT -53.885 -90.81 -53.555 -90.48 ;
        RECT -53.885 -91.965 -53.555 -91.635 ;
        RECT -53.885 -93.325 -53.555 -92.995 ;
        RECT -53.885 -94.685 -53.555 -94.355 ;
        RECT -53.885 -96.045 -53.555 -95.715 ;
        RECT -53.885 -97.405 -53.555 -97.075 ;
        RECT -53.885 -100.125 -53.555 -99.795 ;
        RECT -53.885 -101.35 -53.555 -101.02 ;
        RECT -53.885 -102.845 -53.555 -102.515 ;
        RECT -53.885 -104.205 -53.555 -103.875 ;
        RECT -53.885 -105.565 -53.555 -105.235 ;
        RECT -53.885 -108.285 -53.555 -107.955 ;
        RECT -53.885 -109.645 -53.555 -109.315 ;
        RECT -53.885 -112.365 -53.555 -112.035 ;
        RECT -53.885 -115.085 -53.555 -114.755 ;
        RECT -53.885 -116.445 -53.555 -116.115 ;
        RECT -53.885 -117.805 -53.555 -117.475 ;
        RECT -53.885 -119.165 -53.555 -118.835 ;
        RECT -53.885 -120.525 -53.555 -120.195 ;
        RECT -53.885 -121.885 -53.555 -121.555 ;
        RECT -53.885 -123.245 -53.555 -122.915 ;
        RECT -53.885 -124.605 -53.555 -124.275 ;
        RECT -53.885 -125.965 -53.555 -125.635 ;
        RECT -53.885 -127.325 -53.555 -126.995 ;
        RECT -53.885 -128.685 -53.555 -128.355 ;
        RECT -53.885 -130.045 -53.555 -129.715 ;
        RECT -53.885 -131.405 -53.555 -131.075 ;
        RECT -53.885 -132.765 -53.555 -132.435 ;
        RECT -53.885 -134.125 -53.555 -133.795 ;
        RECT -53.885 -135.485 -53.555 -135.155 ;
        RECT -53.885 -136.845 -53.555 -136.515 ;
        RECT -53.885 -138.205 -53.555 -137.875 ;
        RECT -53.885 -139.565 -53.555 -139.235 ;
        RECT -53.885 -140.925 -53.555 -140.595 ;
        RECT -53.885 -142.285 -53.555 -141.955 ;
        RECT -53.885 -143.645 -53.555 -143.315 ;
        RECT -53.885 -145.005 -53.555 -144.675 ;
        RECT -53.885 -146.365 -53.555 -146.035 ;
        RECT -53.885 -147.725 -53.555 -147.395 ;
        RECT -53.885 -149.085 -53.555 -148.755 ;
        RECT -53.885 -150.445 -53.555 -150.115 ;
        RECT -53.885 -151.805 -53.555 -151.475 ;
        RECT -53.885 -153.165 -53.555 -152.835 ;
        RECT -53.885 -154.525 -53.555 -154.195 ;
        RECT -53.885 -155.885 -53.555 -155.555 ;
        RECT -53.885 -157.245 -53.555 -156.915 ;
        RECT -53.885 -158.605 -53.555 -158.275 ;
        RECT -53.885 -159.965 -53.555 -159.635 ;
        RECT -53.885 -161.325 -53.555 -160.995 ;
        RECT -53.885 -162.685 -53.555 -162.355 ;
        RECT -53.885 -164.045 -53.555 -163.715 ;
        RECT -53.885 -165.405 -53.555 -165.075 ;
        RECT -53.885 -166.765 -53.555 -166.435 ;
        RECT -53.885 -169.485 -53.555 -169.155 ;
        RECT -53.885 -170.845 -53.555 -170.515 ;
        RECT -53.885 -174.925 -53.555 -174.595 ;
        RECT -53.885 -177.645 -53.555 -177.315 ;
        RECT -53.885 -183.29 -53.555 -182.16 ;
        RECT -53.88 -183.405 -53.56 98.08 ;
    END
    PORT
      LAYER met3 ;
        RECT -52.525 244.04 -52.195 245.17 ;
        RECT -52.525 239.875 -52.195 240.205 ;
        RECT -52.525 238.515 -52.195 238.845 ;
        RECT -52.525 237.155 -52.195 237.485 ;
        RECT -52.525 235.795 -52.195 236.125 ;
        RECT -52.525 234.435 -52.195 234.765 ;
        RECT -52.525 233.075 -52.195 233.405 ;
        RECT -52.525 231.715 -52.195 232.045 ;
        RECT -52.525 230.355 -52.195 230.685 ;
        RECT -52.525 228.995 -52.195 229.325 ;
        RECT -52.525 227.635 -52.195 227.965 ;
        RECT -52.525 226.275 -52.195 226.605 ;
        RECT -52.525 224.915 -52.195 225.245 ;
        RECT -52.525 223.555 -52.195 223.885 ;
        RECT -52.525 222.195 -52.195 222.525 ;
        RECT -52.525 220.835 -52.195 221.165 ;
        RECT -52.525 219.475 -52.195 219.805 ;
        RECT -52.525 218.115 -52.195 218.445 ;
        RECT -52.525 216.755 -52.195 217.085 ;
        RECT -52.525 215.395 -52.195 215.725 ;
        RECT -52.525 214.035 -52.195 214.365 ;
        RECT -52.525 212.675 -52.195 213.005 ;
        RECT -52.525 211.315 -52.195 211.645 ;
        RECT -52.525 209.955 -52.195 210.285 ;
        RECT -52.525 208.595 -52.195 208.925 ;
        RECT -52.525 207.235 -52.195 207.565 ;
        RECT -52.525 205.875 -52.195 206.205 ;
        RECT -52.525 204.515 -52.195 204.845 ;
        RECT -52.525 203.155 -52.195 203.485 ;
        RECT -52.525 201.795 -52.195 202.125 ;
        RECT -52.525 200.435 -52.195 200.765 ;
        RECT -52.525 199.075 -52.195 199.405 ;
        RECT -52.525 197.715 -52.195 198.045 ;
        RECT -52.525 196.355 -52.195 196.685 ;
        RECT -52.525 194.995 -52.195 195.325 ;
        RECT -52.525 193.635 -52.195 193.965 ;
        RECT -52.525 192.275 -52.195 192.605 ;
        RECT -52.525 190.915 -52.195 191.245 ;
        RECT -52.525 189.555 -52.195 189.885 ;
        RECT -52.525 188.195 -52.195 188.525 ;
        RECT -52.525 186.835 -52.195 187.165 ;
        RECT -52.525 185.475 -52.195 185.805 ;
        RECT -52.525 184.115 -52.195 184.445 ;
        RECT -52.525 182.755 -52.195 183.085 ;
        RECT -52.525 181.395 -52.195 181.725 ;
        RECT -52.525 180.035 -52.195 180.365 ;
        RECT -52.525 178.675 -52.195 179.005 ;
        RECT -52.525 177.315 -52.195 177.645 ;
        RECT -52.525 175.955 -52.195 176.285 ;
        RECT -52.525 174.595 -52.195 174.925 ;
        RECT -52.525 173.235 -52.195 173.565 ;
        RECT -52.525 171.875 -52.195 172.205 ;
        RECT -52.525 170.515 -52.195 170.845 ;
        RECT -52.525 169.155 -52.195 169.485 ;
        RECT -52.525 167.795 -52.195 168.125 ;
        RECT -52.525 166.435 -52.195 166.765 ;
        RECT -52.525 165.075 -52.195 165.405 ;
        RECT -52.525 163.715 -52.195 164.045 ;
        RECT -52.525 162.355 -52.195 162.685 ;
        RECT -52.525 160.995 -52.195 161.325 ;
        RECT -52.525 159.635 -52.195 159.965 ;
        RECT -52.525 158.275 -52.195 158.605 ;
        RECT -52.525 156.915 -52.195 157.245 ;
        RECT -52.525 155.555 -52.195 155.885 ;
        RECT -52.525 154.195 -52.195 154.525 ;
        RECT -52.525 152.835 -52.195 153.165 ;
        RECT -52.525 151.475 -52.195 151.805 ;
        RECT -52.525 150.115 -52.195 150.445 ;
        RECT -52.525 148.755 -52.195 149.085 ;
        RECT -52.525 147.395 -52.195 147.725 ;
        RECT -52.525 146.035 -52.195 146.365 ;
        RECT -52.525 144.675 -52.195 145.005 ;
        RECT -52.525 143.315 -52.195 143.645 ;
        RECT -52.525 141.955 -52.195 142.285 ;
        RECT -52.525 140.595 -52.195 140.925 ;
        RECT -52.525 139.235 -52.195 139.565 ;
        RECT -52.525 136.42 -52.195 136.75 ;
        RECT -52.525 134.245 -52.195 134.575 ;
        RECT -52.525 133.395 -52.195 133.725 ;
        RECT -52.525 131.085 -52.195 131.415 ;
        RECT -52.525 130.235 -52.195 130.565 ;
        RECT -52.525 127.925 -52.195 128.255 ;
        RECT -52.525 127.075 -52.195 127.405 ;
        RECT -52.525 124.765 -52.195 125.095 ;
        RECT -52.525 123.915 -52.195 124.245 ;
        RECT -52.525 121.605 -52.195 121.935 ;
        RECT -52.525 120.755 -52.195 121.085 ;
        RECT -52.525 118.445 -52.195 118.775 ;
        RECT -52.525 117.595 -52.195 117.925 ;
        RECT -52.52 117.48 -52.2 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -51.165 -64.765 -50.835 -64.435 ;
        RECT -51.165 -66.125 -50.835 -65.795 ;
        RECT -51.165 -67.485 -50.835 -67.155 ;
        RECT -51.165 -68.845 -50.835 -68.515 ;
        RECT -51.165 -70.205 -50.835 -69.875 ;
        RECT -51.165 -71.565 -50.835 -71.235 ;
        RECT -51.165 -72.925 -50.835 -72.595 ;
        RECT -51.165 -74.285 -50.835 -73.955 ;
        RECT -51.165 -75.645 -50.835 -75.315 ;
        RECT -51.165 -77.005 -50.835 -76.675 ;
        RECT -51.165 -78.365 -50.835 -78.035 ;
        RECT -51.165 -79.725 -50.835 -79.395 ;
        RECT -51.165 -81.085 -50.835 -80.755 ;
        RECT -51.165 -82.445 -50.835 -82.115 ;
        RECT -51.165 -83.805 -50.835 -83.475 ;
        RECT -51.165 -85.165 -50.835 -84.835 ;
        RECT -51.165 -86.525 -50.835 -86.195 ;
        RECT -51.165 -87.885 -50.835 -87.555 ;
        RECT -51.165 -89.245 -50.835 -88.915 ;
        RECT -51.165 -90.81 -50.835 -90.48 ;
        RECT -51.165 -91.965 -50.835 -91.635 ;
        RECT -51.165 -93.325 -50.835 -92.995 ;
        RECT -51.165 -94.685 -50.835 -94.355 ;
        RECT -51.165 -96.045 -50.835 -95.715 ;
        RECT -51.165 -97.405 -50.835 -97.075 ;
        RECT -51.165 -100.125 -50.835 -99.795 ;
        RECT -51.165 -101.35 -50.835 -101.02 ;
        RECT -51.165 -102.845 -50.835 -102.515 ;
        RECT -51.165 -104.205 -50.835 -103.875 ;
        RECT -51.165 -105.565 -50.835 -105.235 ;
        RECT -51.165 -108.285 -50.835 -107.955 ;
        RECT -51.165 -109.645 -50.835 -109.315 ;
        RECT -51.165 -113.725 -50.835 -113.395 ;
        RECT -51.165 -115.085 -50.835 -114.755 ;
        RECT -51.165 -116.445 -50.835 -116.115 ;
        RECT -51.165 -117.805 -50.835 -117.475 ;
        RECT -51.165 -119.165 -50.835 -118.835 ;
        RECT -51.165 -120.525 -50.835 -120.195 ;
        RECT -51.165 -121.885 -50.835 -121.555 ;
        RECT -51.165 -123.245 -50.835 -122.915 ;
        RECT -51.165 -124.605 -50.835 -124.275 ;
        RECT -51.165 -125.965 -50.835 -125.635 ;
        RECT -51.165 -127.325 -50.835 -126.995 ;
        RECT -51.165 -128.685 -50.835 -128.355 ;
        RECT -51.165 -130.045 -50.835 -129.715 ;
        RECT -51.165 -131.405 -50.835 -131.075 ;
        RECT -51.165 -132.765 -50.835 -132.435 ;
        RECT -51.165 -134.125 -50.835 -133.795 ;
        RECT -51.165 -135.485 -50.835 -135.155 ;
        RECT -51.165 -136.845 -50.835 -136.515 ;
        RECT -51.165 -138.205 -50.835 -137.875 ;
        RECT -51.165 -139.565 -50.835 -139.235 ;
        RECT -51.165 -140.925 -50.835 -140.595 ;
        RECT -51.165 -142.285 -50.835 -141.955 ;
        RECT -51.165 -143.645 -50.835 -143.315 ;
        RECT -51.165 -145.005 -50.835 -144.675 ;
        RECT -51.165 -146.365 -50.835 -146.035 ;
        RECT -51.165 -147.725 -50.835 -147.395 ;
        RECT -51.165 -149.085 -50.835 -148.755 ;
        RECT -51.165 -150.445 -50.835 -150.115 ;
        RECT -51.165 -151.805 -50.835 -151.475 ;
        RECT -51.165 -153.165 -50.835 -152.835 ;
        RECT -51.165 -154.525 -50.835 -154.195 ;
        RECT -51.165 -155.885 -50.835 -155.555 ;
        RECT -51.165 -157.245 -50.835 -156.915 ;
        RECT -51.165 -158.605 -50.835 -158.275 ;
        RECT -51.165 -159.965 -50.835 -159.635 ;
        RECT -51.165 -161.325 -50.835 -160.995 ;
        RECT -51.165 -162.685 -50.835 -162.355 ;
        RECT -51.165 -164.045 -50.835 -163.715 ;
        RECT -51.165 -165.405 -50.835 -165.075 ;
        RECT -51.165 -166.765 -50.835 -166.435 ;
        RECT -51.165 -168.655 -50.835 -168.325 ;
        RECT -51.165 -169.485 -50.835 -169.155 ;
        RECT -51.165 -170.845 -50.835 -170.515 ;
        RECT -51.165 -173.565 -50.835 -173.235 ;
        RECT -51.165 -174.925 -50.835 -174.595 ;
        RECT -51.165 -177.645 -50.835 -177.315 ;
        RECT -51.165 -183.29 -50.835 -182.16 ;
        RECT -51.16 -183.405 -50.84 245.285 ;
        RECT -51.165 244.04 -50.835 245.17 ;
        RECT -51.165 239.875 -50.835 240.205 ;
        RECT -51.165 238.515 -50.835 238.845 ;
        RECT -51.165 237.155 -50.835 237.485 ;
        RECT -51.165 235.795 -50.835 236.125 ;
        RECT -51.165 234.435 -50.835 234.765 ;
        RECT -51.165 233.075 -50.835 233.405 ;
        RECT -51.165 231.715 -50.835 232.045 ;
        RECT -51.165 230.355 -50.835 230.685 ;
        RECT -51.165 228.995 -50.835 229.325 ;
        RECT -51.165 227.635 -50.835 227.965 ;
        RECT -51.165 226.275 -50.835 226.605 ;
        RECT -51.165 224.915 -50.835 225.245 ;
        RECT -51.165 223.555 -50.835 223.885 ;
        RECT -51.165 222.195 -50.835 222.525 ;
        RECT -51.165 220.835 -50.835 221.165 ;
        RECT -51.165 219.475 -50.835 219.805 ;
        RECT -51.165 218.115 -50.835 218.445 ;
        RECT -51.165 216.755 -50.835 217.085 ;
        RECT -51.165 215.395 -50.835 215.725 ;
        RECT -51.165 214.035 -50.835 214.365 ;
        RECT -51.165 212.675 -50.835 213.005 ;
        RECT -51.165 211.315 -50.835 211.645 ;
        RECT -51.165 209.955 -50.835 210.285 ;
        RECT -51.165 208.595 -50.835 208.925 ;
        RECT -51.165 207.235 -50.835 207.565 ;
        RECT -51.165 205.875 -50.835 206.205 ;
        RECT -51.165 204.515 -50.835 204.845 ;
        RECT -51.165 203.155 -50.835 203.485 ;
        RECT -51.165 201.795 -50.835 202.125 ;
        RECT -51.165 200.435 -50.835 200.765 ;
        RECT -51.165 199.075 -50.835 199.405 ;
        RECT -51.165 197.715 -50.835 198.045 ;
        RECT -51.165 196.355 -50.835 196.685 ;
        RECT -51.165 194.995 -50.835 195.325 ;
        RECT -51.165 193.635 -50.835 193.965 ;
        RECT -51.165 192.275 -50.835 192.605 ;
        RECT -51.165 190.915 -50.835 191.245 ;
        RECT -51.165 189.555 -50.835 189.885 ;
        RECT -51.165 188.195 -50.835 188.525 ;
        RECT -51.165 186.835 -50.835 187.165 ;
        RECT -51.165 185.475 -50.835 185.805 ;
        RECT -51.165 184.115 -50.835 184.445 ;
        RECT -51.165 182.755 -50.835 183.085 ;
        RECT -51.165 181.395 -50.835 181.725 ;
        RECT -51.165 180.035 -50.835 180.365 ;
        RECT -51.165 178.675 -50.835 179.005 ;
        RECT -51.165 177.315 -50.835 177.645 ;
        RECT -51.165 175.955 -50.835 176.285 ;
        RECT -51.165 174.595 -50.835 174.925 ;
        RECT -51.165 173.235 -50.835 173.565 ;
        RECT -51.165 171.875 -50.835 172.205 ;
        RECT -51.165 170.515 -50.835 170.845 ;
        RECT -51.165 169.155 -50.835 169.485 ;
        RECT -51.165 167.795 -50.835 168.125 ;
        RECT -51.165 166.435 -50.835 166.765 ;
        RECT -51.165 165.075 -50.835 165.405 ;
        RECT -51.165 163.715 -50.835 164.045 ;
        RECT -51.165 162.355 -50.835 162.685 ;
        RECT -51.165 160.995 -50.835 161.325 ;
        RECT -51.165 159.635 -50.835 159.965 ;
        RECT -51.165 158.275 -50.835 158.605 ;
        RECT -51.165 156.915 -50.835 157.245 ;
        RECT -51.165 155.555 -50.835 155.885 ;
        RECT -51.165 154.195 -50.835 154.525 ;
        RECT -51.165 152.835 -50.835 153.165 ;
        RECT -51.165 151.475 -50.835 151.805 ;
        RECT -51.165 150.115 -50.835 150.445 ;
        RECT -51.165 148.755 -50.835 149.085 ;
        RECT -51.165 147.395 -50.835 147.725 ;
        RECT -51.165 146.035 -50.835 146.365 ;
        RECT -51.165 144.675 -50.835 145.005 ;
        RECT -51.165 143.315 -50.835 143.645 ;
        RECT -51.165 141.955 -50.835 142.285 ;
        RECT -51.165 140.595 -50.835 140.925 ;
        RECT -51.165 139.235 -50.835 139.565 ;
        RECT -51.165 136.42 -50.835 136.75 ;
        RECT -51.165 134.245 -50.835 134.575 ;
        RECT -51.165 133.395 -50.835 133.725 ;
        RECT -51.165 131.085 -50.835 131.415 ;
        RECT -51.165 130.235 -50.835 130.565 ;
        RECT -51.165 127.925 -50.835 128.255 ;
        RECT -51.165 127.075 -50.835 127.405 ;
        RECT -51.165 124.765 -50.835 125.095 ;
        RECT -51.165 123.915 -50.835 124.245 ;
        RECT -51.165 121.605 -50.835 121.935 ;
        RECT -51.165 120.755 -50.835 121.085 ;
        RECT -51.165 118.445 -50.835 118.775 ;
        RECT -51.165 117.595 -50.835 117.925 ;
        RECT -51.165 115.285 -50.835 115.615 ;
        RECT -51.165 114.435 -50.835 114.765 ;
        RECT -51.165 112.125 -50.835 112.455 ;
        RECT -51.165 111.275 -50.835 111.605 ;
        RECT -51.165 108.965 -50.835 109.295 ;
        RECT -51.165 108.115 -50.835 108.445 ;
        RECT -51.165 105.805 -50.835 106.135 ;
        RECT -51.165 104.955 -50.835 105.285 ;
        RECT -51.165 102.645 -50.835 102.975 ;
        RECT -51.165 101.795 -50.835 102.125 ;
        RECT -51.165 99.62 -50.835 99.95 ;
        RECT -51.165 97.075 -50.835 97.405 ;
        RECT -51.165 95.715 -50.835 96.045 ;
        RECT -51.165 94.355 -50.835 94.685 ;
        RECT -51.165 92.995 -50.835 93.325 ;
        RECT -51.165 91.635 -50.835 91.965 ;
        RECT -51.165 90.275 -50.835 90.605 ;
        RECT -51.165 88.915 -50.835 89.245 ;
        RECT -51.165 87.555 -50.835 87.885 ;
        RECT -51.165 86.195 -50.835 86.525 ;
        RECT -51.165 84.835 -50.835 85.165 ;
        RECT -51.165 83.475 -50.835 83.805 ;
        RECT -51.165 82.115 -50.835 82.445 ;
        RECT -51.165 80.755 -50.835 81.085 ;
        RECT -51.165 79.395 -50.835 79.725 ;
        RECT -51.165 78.035 -50.835 78.365 ;
        RECT -51.165 76.675 -50.835 77.005 ;
        RECT -51.165 75.315 -50.835 75.645 ;
        RECT -51.165 73.955 -50.835 74.285 ;
        RECT -51.165 72.595 -50.835 72.925 ;
        RECT -51.165 71.235 -50.835 71.565 ;
        RECT -51.165 69.875 -50.835 70.205 ;
        RECT -51.165 68.515 -50.835 68.845 ;
        RECT -51.165 67.155 -50.835 67.485 ;
        RECT -51.165 65.795 -50.835 66.125 ;
        RECT -51.165 64.435 -50.835 64.765 ;
        RECT -51.165 63.075 -50.835 63.405 ;
        RECT -51.165 61.715 -50.835 62.045 ;
        RECT -51.165 60.355 -50.835 60.685 ;
        RECT -51.165 58.995 -50.835 59.325 ;
        RECT -51.165 57.635 -50.835 57.965 ;
        RECT -51.165 56.275 -50.835 56.605 ;
        RECT -51.165 54.915 -50.835 55.245 ;
        RECT -51.165 53.555 -50.835 53.885 ;
        RECT -51.165 52.195 -50.835 52.525 ;
        RECT -51.165 50.835 -50.835 51.165 ;
        RECT -51.165 49.475 -50.835 49.805 ;
        RECT -51.165 48.115 -50.835 48.445 ;
        RECT -51.165 46.755 -50.835 47.085 ;
        RECT -51.165 45.395 -50.835 45.725 ;
        RECT -51.165 44.035 -50.835 44.365 ;
        RECT -51.165 42.675 -50.835 43.005 ;
        RECT -51.165 41.315 -50.835 41.645 ;
        RECT -51.165 39.955 -50.835 40.285 ;
        RECT -51.165 38.595 -50.835 38.925 ;
        RECT -51.165 37.235 -50.835 37.565 ;
        RECT -51.165 35.875 -50.835 36.205 ;
        RECT -51.165 34.515 -50.835 34.845 ;
        RECT -51.165 33.155 -50.835 33.485 ;
        RECT -51.165 31.795 -50.835 32.125 ;
        RECT -51.165 30.435 -50.835 30.765 ;
        RECT -51.165 29.075 -50.835 29.405 ;
        RECT -51.165 27.715 -50.835 28.045 ;
        RECT -51.165 26.355 -50.835 26.685 ;
        RECT -51.165 24.995 -50.835 25.325 ;
        RECT -51.165 23.635 -50.835 23.965 ;
        RECT -51.165 22.275 -50.835 22.605 ;
        RECT -51.165 20.915 -50.835 21.245 ;
        RECT -51.165 19.555 -50.835 19.885 ;
        RECT -51.165 18.195 -50.835 18.525 ;
        RECT -51.165 16.835 -50.835 17.165 ;
        RECT -51.165 15.475 -50.835 15.805 ;
        RECT -51.165 14.115 -50.835 14.445 ;
        RECT -51.165 12.755 -50.835 13.085 ;
        RECT -51.165 11.395 -50.835 11.725 ;
        RECT -51.165 10.035 -50.835 10.365 ;
        RECT -51.165 8.675 -50.835 9.005 ;
        RECT -51.165 7.315 -50.835 7.645 ;
        RECT -51.165 5.955 -50.835 6.285 ;
        RECT -51.165 4.595 -50.835 4.925 ;
        RECT -51.165 3.235 -50.835 3.565 ;
        RECT -51.165 1.875 -50.835 2.205 ;
        RECT -51.165 0.515 -50.835 0.845 ;
        RECT -51.165 -0.845 -50.835 -0.515 ;
        RECT -51.165 -2.205 -50.835 -1.875 ;
        RECT -51.165 -3.565 -50.835 -3.235 ;
        RECT -51.165 -4.925 -50.835 -4.595 ;
        RECT -51.165 -6.285 -50.835 -5.955 ;
        RECT -51.165 -7.645 -50.835 -7.315 ;
        RECT -51.165 -9.005 -50.835 -8.675 ;
        RECT -51.165 -10.365 -50.835 -10.035 ;
        RECT -51.165 -11.725 -50.835 -11.395 ;
        RECT -51.165 -13.085 -50.835 -12.755 ;
        RECT -51.165 -14.445 -50.835 -14.115 ;
        RECT -51.165 -15.805 -50.835 -15.475 ;
        RECT -51.165 -17.165 -50.835 -16.835 ;
        RECT -51.165 -18.525 -50.835 -18.195 ;
        RECT -51.165 -19.885 -50.835 -19.555 ;
        RECT -51.165 -21.245 -50.835 -20.915 ;
        RECT -51.165 -22.605 -50.835 -22.275 ;
        RECT -51.165 -23.965 -50.835 -23.635 ;
        RECT -51.165 -25.325 -50.835 -24.995 ;
        RECT -51.165 -29.405 -50.835 -29.075 ;
        RECT -51.165 -30.765 -50.835 -30.435 ;
        RECT -51.165 -32.125 -50.835 -31.795 ;
        RECT -51.165 -33.485 -50.835 -33.155 ;
        RECT -51.165 -34.845 -50.835 -34.515 ;
        RECT -51.165 -36.205 -50.835 -35.875 ;
        RECT -51.165 -37.565 -50.835 -37.235 ;
        RECT -51.165 -38.925 -50.835 -38.595 ;
        RECT -51.165 -40.285 -50.835 -39.955 ;
        RECT -51.165 -41.645 -50.835 -41.315 ;
        RECT -51.165 -43.005 -50.835 -42.675 ;
        RECT -51.165 -44.365 -50.835 -44.035 ;
        RECT -51.165 -45.725 -50.835 -45.395 ;
        RECT -51.165 -47.085 -50.835 -46.755 ;
        RECT -51.165 -48.445 -50.835 -48.115 ;
        RECT -51.165 -49.805 -50.835 -49.475 ;
        RECT -51.165 -51.165 -50.835 -50.835 ;
        RECT -51.165 -52.525 -50.835 -52.195 ;
        RECT -51.165 -53.885 -50.835 -53.555 ;
        RECT -51.165 -55.245 -50.835 -54.915 ;
        RECT -51.165 -56.605 -50.835 -56.275 ;
        RECT -51.165 -57.965 -50.835 -57.635 ;
        RECT -51.165 -59.325 -50.835 -58.995 ;
        RECT -51.165 -60.685 -50.835 -60.355 ;
        RECT -51.165 -62.045 -50.835 -61.715 ;
        RECT -51.165 -63.405 -50.835 -63.075 ;
    END
    PORT
      LAYER met3 ;
        RECT -62.045 -120.525 -61.715 -120.195 ;
        RECT -62.045 -121.885 -61.715 -121.555 ;
        RECT -62.045 -123.245 -61.715 -122.915 ;
        RECT -62.045 -124.605 -61.715 -124.275 ;
        RECT -62.045 -125.965 -61.715 -125.635 ;
        RECT -62.045 -127.325 -61.715 -126.995 ;
        RECT -62.045 -128.685 -61.715 -128.355 ;
        RECT -62.045 -130.045 -61.715 -129.715 ;
        RECT -62.045 -131.405 -61.715 -131.075 ;
        RECT -62.045 -132.765 -61.715 -132.435 ;
        RECT -62.045 -134.125 -61.715 -133.795 ;
        RECT -62.045 -135.485 -61.715 -135.155 ;
        RECT -62.045 -136.845 -61.715 -136.515 ;
        RECT -62.045 -138.205 -61.715 -137.875 ;
        RECT -62.045 -139.565 -61.715 -139.235 ;
        RECT -62.045 -140.925 -61.715 -140.595 ;
        RECT -62.045 -142.285 -61.715 -141.955 ;
        RECT -62.045 -143.645 -61.715 -143.315 ;
        RECT -62.045 -145.005 -61.715 -144.675 ;
        RECT -62.045 -146.365 -61.715 -146.035 ;
        RECT -62.045 -147.725 -61.715 -147.395 ;
        RECT -62.045 -149.085 -61.715 -148.755 ;
        RECT -62.045 -150.445 -61.715 -150.115 ;
        RECT -62.045 -151.805 -61.715 -151.475 ;
        RECT -62.045 -153.165 -61.715 -152.835 ;
        RECT -62.045 -154.525 -61.715 -154.195 ;
        RECT -62.045 -155.885 -61.715 -155.555 ;
        RECT -62.045 -157.245 -61.715 -156.915 ;
        RECT -62.045 -158.605 -61.715 -158.275 ;
        RECT -62.045 -159.965 -61.715 -159.635 ;
        RECT -62.045 -161.325 -61.715 -160.995 ;
        RECT -62.045 -162.685 -61.715 -162.355 ;
        RECT -62.045 -164.045 -61.715 -163.715 ;
        RECT -62.045 -165.405 -61.715 -165.075 ;
        RECT -62.045 -166.765 -61.715 -166.435 ;
        RECT -62.045 -168.655 -61.715 -168.325 ;
        RECT -62.045 -169.485 -61.715 -169.155 ;
        RECT -62.045 -170.845 -61.715 -170.515 ;
        RECT -62.045 -172.205 -61.715 -171.875 ;
        RECT -62.045 -174.925 -61.715 -174.595 ;
        RECT -62.045 -177.645 -61.715 -177.315 ;
        RECT -62.045 -183.29 -61.715 -182.16 ;
        RECT -62.04 -183.405 -61.72 -120.195 ;
    END
    PORT
      LAYER met3 ;
        RECT -60.685 244.04 -60.355 245.17 ;
        RECT -60.685 239.875 -60.355 240.205 ;
        RECT -60.685 238.515 -60.355 238.845 ;
        RECT -60.685 237.155 -60.355 237.485 ;
        RECT -60.685 235.795 -60.355 236.125 ;
        RECT -60.685 234.435 -60.355 234.765 ;
        RECT -60.685 233.075 -60.355 233.405 ;
        RECT -60.685 231.715 -60.355 232.045 ;
        RECT -60.685 230.355 -60.355 230.685 ;
        RECT -60.685 228.995 -60.355 229.325 ;
        RECT -60.685 227.635 -60.355 227.965 ;
        RECT -60.685 226.275 -60.355 226.605 ;
        RECT -60.685 224.915 -60.355 225.245 ;
        RECT -60.685 223.555 -60.355 223.885 ;
        RECT -60.685 222.195 -60.355 222.525 ;
        RECT -60.685 220.835 -60.355 221.165 ;
        RECT -60.685 219.475 -60.355 219.805 ;
        RECT -60.685 218.115 -60.355 218.445 ;
        RECT -60.685 216.755 -60.355 217.085 ;
        RECT -60.685 215.395 -60.355 215.725 ;
        RECT -60.685 214.035 -60.355 214.365 ;
        RECT -60.685 212.675 -60.355 213.005 ;
        RECT -60.685 211.315 -60.355 211.645 ;
        RECT -60.685 209.955 -60.355 210.285 ;
        RECT -60.685 208.595 -60.355 208.925 ;
        RECT -60.685 207.235 -60.355 207.565 ;
        RECT -60.685 205.875 -60.355 206.205 ;
        RECT -60.685 204.515 -60.355 204.845 ;
        RECT -60.685 203.155 -60.355 203.485 ;
        RECT -60.685 201.795 -60.355 202.125 ;
        RECT -60.685 200.435 -60.355 200.765 ;
        RECT -60.685 199.075 -60.355 199.405 ;
        RECT -60.685 197.715 -60.355 198.045 ;
        RECT -60.685 196.355 -60.355 196.685 ;
        RECT -60.685 194.995 -60.355 195.325 ;
        RECT -60.685 193.635 -60.355 193.965 ;
        RECT -60.685 192.275 -60.355 192.605 ;
        RECT -60.685 190.915 -60.355 191.245 ;
        RECT -60.685 189.555 -60.355 189.885 ;
        RECT -60.685 188.195 -60.355 188.525 ;
        RECT -60.685 186.835 -60.355 187.165 ;
        RECT -60.685 185.475 -60.355 185.805 ;
        RECT -60.685 184.115 -60.355 184.445 ;
        RECT -60.685 182.755 -60.355 183.085 ;
        RECT -60.685 181.395 -60.355 181.725 ;
        RECT -60.685 180.035 -60.355 180.365 ;
        RECT -60.685 178.675 -60.355 179.005 ;
        RECT -60.685 177.315 -60.355 177.645 ;
        RECT -60.685 175.955 -60.355 176.285 ;
        RECT -60.685 174.595 -60.355 174.925 ;
        RECT -60.685 173.235 -60.355 173.565 ;
        RECT -60.685 171.875 -60.355 172.205 ;
        RECT -60.685 170.515 -60.355 170.845 ;
        RECT -60.685 169.155 -60.355 169.485 ;
        RECT -60.685 167.795 -60.355 168.125 ;
        RECT -60.685 166.435 -60.355 166.765 ;
        RECT -60.685 165.075 -60.355 165.405 ;
        RECT -60.685 163.715 -60.355 164.045 ;
        RECT -60.685 162.355 -60.355 162.685 ;
        RECT -60.685 160.995 -60.355 161.325 ;
        RECT -60.685 159.635 -60.355 159.965 ;
        RECT -60.685 158.275 -60.355 158.605 ;
        RECT -60.685 156.915 -60.355 157.245 ;
        RECT -60.685 155.555 -60.355 155.885 ;
        RECT -60.685 154.195 -60.355 154.525 ;
        RECT -60.685 152.835 -60.355 153.165 ;
        RECT -60.685 151.475 -60.355 151.805 ;
        RECT -60.685 150.115 -60.355 150.445 ;
        RECT -60.685 148.755 -60.355 149.085 ;
        RECT -60.685 147.395 -60.355 147.725 ;
        RECT -60.685 146.035 -60.355 146.365 ;
        RECT -60.685 144.675 -60.355 145.005 ;
        RECT -60.685 143.315 -60.355 143.645 ;
        RECT -60.685 141.955 -60.355 142.285 ;
        RECT -60.685 140.595 -60.355 140.925 ;
        RECT -60.685 139.235 -60.355 139.565 ;
        RECT -60.685 136.42 -60.355 136.75 ;
        RECT -60.685 134.245 -60.355 134.575 ;
        RECT -60.685 133.395 -60.355 133.725 ;
        RECT -60.685 131.085 -60.355 131.415 ;
        RECT -60.685 130.235 -60.355 130.565 ;
        RECT -60.685 127.925 -60.355 128.255 ;
        RECT -60.685 127.075 -60.355 127.405 ;
        RECT -60.685 124.765 -60.355 125.095 ;
        RECT -60.685 123.915 -60.355 124.245 ;
        RECT -60.685 121.605 -60.355 121.935 ;
        RECT -60.685 120.755 -60.355 121.085 ;
        RECT -60.685 118.445 -60.355 118.775 ;
        RECT -60.685 117.595 -60.355 117.925 ;
        RECT -60.685 115.285 -60.355 115.615 ;
        RECT -60.685 114.435 -60.355 114.765 ;
        RECT -60.685 112.125 -60.355 112.455 ;
        RECT -60.685 111.275 -60.355 111.605 ;
        RECT -60.685 108.965 -60.355 109.295 ;
        RECT -60.685 108.115 -60.355 108.445 ;
        RECT -60.685 105.805 -60.355 106.135 ;
        RECT -60.685 104.955 -60.355 105.285 ;
        RECT -60.685 102.645 -60.355 102.975 ;
        RECT -60.685 101.795 -60.355 102.125 ;
        RECT -60.685 99.62 -60.355 99.95 ;
        RECT -60.685 97.075 -60.355 97.405 ;
        RECT -60.685 95.715 -60.355 96.045 ;
        RECT -60.685 94.355 -60.355 94.685 ;
        RECT -60.685 92.995 -60.355 93.325 ;
        RECT -60.685 91.635 -60.355 91.965 ;
        RECT -60.685 90.275 -60.355 90.605 ;
        RECT -60.685 88.915 -60.355 89.245 ;
        RECT -60.685 87.555 -60.355 87.885 ;
        RECT -60.685 86.195 -60.355 86.525 ;
        RECT -60.685 84.835 -60.355 85.165 ;
        RECT -60.685 83.475 -60.355 83.805 ;
        RECT -60.685 82.115 -60.355 82.445 ;
        RECT -60.685 80.755 -60.355 81.085 ;
        RECT -60.685 79.395 -60.355 79.725 ;
        RECT -60.685 78.035 -60.355 78.365 ;
        RECT -60.685 76.675 -60.355 77.005 ;
        RECT -60.685 75.315 -60.355 75.645 ;
        RECT -60.685 73.955 -60.355 74.285 ;
        RECT -60.685 72.595 -60.355 72.925 ;
        RECT -60.685 71.235 -60.355 71.565 ;
        RECT -60.685 69.875 -60.355 70.205 ;
        RECT -60.685 68.515 -60.355 68.845 ;
        RECT -60.685 67.155 -60.355 67.485 ;
        RECT -60.685 65.795 -60.355 66.125 ;
        RECT -60.685 64.435 -60.355 64.765 ;
        RECT -60.685 63.075 -60.355 63.405 ;
        RECT -60.685 61.715 -60.355 62.045 ;
        RECT -60.685 60.355 -60.355 60.685 ;
        RECT -60.685 58.995 -60.355 59.325 ;
        RECT -60.685 57.635 -60.355 57.965 ;
        RECT -60.685 56.275 -60.355 56.605 ;
        RECT -60.685 54.915 -60.355 55.245 ;
        RECT -60.685 53.555 -60.355 53.885 ;
        RECT -60.685 52.195 -60.355 52.525 ;
        RECT -60.685 50.835 -60.355 51.165 ;
        RECT -60.685 49.475 -60.355 49.805 ;
        RECT -60.685 48.115 -60.355 48.445 ;
        RECT -60.685 46.755 -60.355 47.085 ;
        RECT -60.685 45.395 -60.355 45.725 ;
        RECT -60.685 44.035 -60.355 44.365 ;
        RECT -60.685 42.675 -60.355 43.005 ;
        RECT -60.685 41.315 -60.355 41.645 ;
        RECT -60.685 39.955 -60.355 40.285 ;
        RECT -60.685 38.595 -60.355 38.925 ;
        RECT -60.685 37.235 -60.355 37.565 ;
        RECT -60.685 35.875 -60.355 36.205 ;
        RECT -60.685 34.515 -60.355 34.845 ;
        RECT -60.685 33.155 -60.355 33.485 ;
        RECT -60.685 31.795 -60.355 32.125 ;
        RECT -60.685 30.435 -60.355 30.765 ;
        RECT -60.685 29.075 -60.355 29.405 ;
        RECT -60.685 27.715 -60.355 28.045 ;
        RECT -60.685 26.355 -60.355 26.685 ;
        RECT -60.685 24.995 -60.355 25.325 ;
        RECT -60.685 23.635 -60.355 23.965 ;
        RECT -60.685 22.275 -60.355 22.605 ;
        RECT -60.685 20.915 -60.355 21.245 ;
        RECT -60.685 19.555 -60.355 19.885 ;
        RECT -60.685 18.195 -60.355 18.525 ;
        RECT -60.685 16.835 -60.355 17.165 ;
        RECT -60.685 15.475 -60.355 15.805 ;
        RECT -60.685 14.115 -60.355 14.445 ;
        RECT -60.685 12.755 -60.355 13.085 ;
        RECT -60.685 11.395 -60.355 11.725 ;
        RECT -60.685 10.035 -60.355 10.365 ;
        RECT -60.685 8.675 -60.355 9.005 ;
        RECT -60.685 7.315 -60.355 7.645 ;
        RECT -60.685 5.955 -60.355 6.285 ;
        RECT -60.685 4.595 -60.355 4.925 ;
        RECT -60.685 3.235 -60.355 3.565 ;
        RECT -60.685 1.875 -60.355 2.205 ;
        RECT -60.685 0.515 -60.355 0.845 ;
        RECT -60.685 -0.845 -60.355 -0.515 ;
        RECT -60.685 -2.205 -60.355 -1.875 ;
        RECT -60.685 -3.565 -60.355 -3.235 ;
        RECT -60.685 -4.925 -60.355 -4.595 ;
        RECT -60.685 -6.285 -60.355 -5.955 ;
        RECT -60.685 -7.645 -60.355 -7.315 ;
        RECT -60.685 -9.005 -60.355 -8.675 ;
        RECT -60.685 -10.365 -60.355 -10.035 ;
        RECT -60.685 -11.725 -60.355 -11.395 ;
        RECT -60.685 -13.085 -60.355 -12.755 ;
        RECT -60.685 -14.445 -60.355 -14.115 ;
        RECT -60.685 -15.805 -60.355 -15.475 ;
        RECT -60.685 -17.165 -60.355 -16.835 ;
        RECT -60.685 -18.525 -60.355 -18.195 ;
        RECT -60.685 -19.885 -60.355 -19.555 ;
        RECT -60.685 -21.245 -60.355 -20.915 ;
        RECT -60.685 -22.605 -60.355 -22.275 ;
        RECT -60.685 -23.965 -60.355 -23.635 ;
        RECT -60.685 -25.325 -60.355 -24.995 ;
        RECT -60.685 -26.685 -60.355 -26.355 ;
        RECT -60.685 -28.045 -60.355 -27.715 ;
        RECT -60.685 -29.405 -60.355 -29.075 ;
        RECT -60.685 -30.765 -60.355 -30.435 ;
        RECT -60.685 -32.125 -60.355 -31.795 ;
        RECT -60.685 -33.485 -60.355 -33.155 ;
        RECT -60.685 -34.845 -60.355 -34.515 ;
        RECT -60.685 -36.205 -60.355 -35.875 ;
        RECT -60.685 -37.565 -60.355 -37.235 ;
        RECT -60.685 -38.925 -60.355 -38.595 ;
        RECT -60.685 -40.285 -60.355 -39.955 ;
        RECT -60.685 -41.645 -60.355 -41.315 ;
        RECT -60.685 -43.005 -60.355 -42.675 ;
        RECT -60.685 -44.365 -60.355 -44.035 ;
        RECT -60.685 -45.725 -60.355 -45.395 ;
        RECT -60.685 -47.085 -60.355 -46.755 ;
        RECT -60.685 -48.445 -60.355 -48.115 ;
        RECT -60.685 -49.805 -60.355 -49.475 ;
        RECT -60.685 -51.165 -60.355 -50.835 ;
        RECT -60.685 -52.525 -60.355 -52.195 ;
        RECT -60.685 -53.885 -60.355 -53.555 ;
        RECT -60.685 -55.245 -60.355 -54.915 ;
        RECT -60.685 -56.605 -60.355 -56.275 ;
        RECT -60.685 -57.965 -60.355 -57.635 ;
        RECT -60.685 -59.325 -60.355 -58.995 ;
        RECT -60.685 -60.685 -60.355 -60.355 ;
        RECT -60.685 -62.045 -60.355 -61.715 ;
        RECT -60.685 -63.405 -60.355 -63.075 ;
        RECT -60.685 -64.765 -60.355 -64.435 ;
        RECT -60.685 -66.125 -60.355 -65.795 ;
        RECT -60.685 -67.485 -60.355 -67.155 ;
        RECT -60.685 -68.845 -60.355 -68.515 ;
        RECT -60.685 -70.205 -60.355 -69.875 ;
        RECT -60.685 -71.565 -60.355 -71.235 ;
        RECT -60.685 -72.925 -60.355 -72.595 ;
        RECT -60.685 -74.285 -60.355 -73.955 ;
        RECT -60.685 -75.645 -60.355 -75.315 ;
        RECT -60.685 -77.005 -60.355 -76.675 ;
        RECT -60.685 -78.365 -60.355 -78.035 ;
        RECT -60.685 -79.725 -60.355 -79.395 ;
        RECT -60.685 -81.085 -60.355 -80.755 ;
        RECT -60.685 -82.445 -60.355 -82.115 ;
        RECT -60.685 -83.805 -60.355 -83.475 ;
        RECT -60.685 -85.165 -60.355 -84.835 ;
        RECT -60.685 -86.525 -60.355 -86.195 ;
        RECT -60.685 -87.885 -60.355 -87.555 ;
        RECT -60.685 -89.245 -60.355 -88.915 ;
        RECT -60.685 -90.81 -60.355 -90.48 ;
        RECT -60.685 -91.965 -60.355 -91.635 ;
        RECT -60.685 -93.325 -60.355 -92.995 ;
        RECT -60.685 -94.685 -60.355 -94.355 ;
        RECT -60.685 -96.045 -60.355 -95.715 ;
        RECT -60.685 -97.405 -60.355 -97.075 ;
        RECT -60.685 -100.125 -60.355 -99.795 ;
        RECT -60.685 -101.35 -60.355 -101.02 ;
        RECT -60.685 -102.845 -60.355 -102.515 ;
        RECT -60.685 -104.205 -60.355 -103.875 ;
        RECT -60.685 -105.565 -60.355 -105.235 ;
        RECT -60.685 -108.285 -60.355 -107.955 ;
        RECT -60.685 -109.645 -60.355 -109.315 ;
        RECT -60.685 -113.725 -60.355 -113.395 ;
        RECT -60.68 -113.725 -60.36 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -60.685 -174.925 -60.355 -174.595 ;
        RECT -60.685 -177.645 -60.355 -177.315 ;
        RECT -60.685 -183.29 -60.355 -182.16 ;
        RECT -60.68 -183.405 -60.36 -173.92 ;
    END
    PORT
      LAYER met3 ;
        RECT -59.325 244.04 -58.995 245.17 ;
        RECT -59.325 239.875 -58.995 240.205 ;
        RECT -59.325 238.515 -58.995 238.845 ;
        RECT -59.325 237.155 -58.995 237.485 ;
        RECT -59.325 235.795 -58.995 236.125 ;
        RECT -59.325 234.435 -58.995 234.765 ;
        RECT -59.325 233.075 -58.995 233.405 ;
        RECT -59.325 231.715 -58.995 232.045 ;
        RECT -59.325 230.355 -58.995 230.685 ;
        RECT -59.325 228.995 -58.995 229.325 ;
        RECT -59.325 227.635 -58.995 227.965 ;
        RECT -59.325 226.275 -58.995 226.605 ;
        RECT -59.325 224.915 -58.995 225.245 ;
        RECT -59.325 223.555 -58.995 223.885 ;
        RECT -59.325 222.195 -58.995 222.525 ;
        RECT -59.325 220.835 -58.995 221.165 ;
        RECT -59.325 219.475 -58.995 219.805 ;
        RECT -59.325 218.115 -58.995 218.445 ;
        RECT -59.325 216.755 -58.995 217.085 ;
        RECT -59.325 215.395 -58.995 215.725 ;
        RECT -59.325 214.035 -58.995 214.365 ;
        RECT -59.325 212.675 -58.995 213.005 ;
        RECT -59.325 211.315 -58.995 211.645 ;
        RECT -59.325 209.955 -58.995 210.285 ;
        RECT -59.325 208.595 -58.995 208.925 ;
        RECT -59.325 207.235 -58.995 207.565 ;
        RECT -59.325 205.875 -58.995 206.205 ;
        RECT -59.325 204.515 -58.995 204.845 ;
        RECT -59.325 203.155 -58.995 203.485 ;
        RECT -59.325 201.795 -58.995 202.125 ;
        RECT -59.325 200.435 -58.995 200.765 ;
        RECT -59.325 199.075 -58.995 199.405 ;
        RECT -59.325 197.715 -58.995 198.045 ;
        RECT -59.325 196.355 -58.995 196.685 ;
        RECT -59.325 194.995 -58.995 195.325 ;
        RECT -59.325 193.635 -58.995 193.965 ;
        RECT -59.325 192.275 -58.995 192.605 ;
        RECT -59.325 190.915 -58.995 191.245 ;
        RECT -59.325 189.555 -58.995 189.885 ;
        RECT -59.325 188.195 -58.995 188.525 ;
        RECT -59.325 186.835 -58.995 187.165 ;
        RECT -59.325 185.475 -58.995 185.805 ;
        RECT -59.325 184.115 -58.995 184.445 ;
        RECT -59.325 182.755 -58.995 183.085 ;
        RECT -59.325 181.395 -58.995 181.725 ;
        RECT -59.325 180.035 -58.995 180.365 ;
        RECT -59.325 178.675 -58.995 179.005 ;
        RECT -59.325 177.315 -58.995 177.645 ;
        RECT -59.325 175.955 -58.995 176.285 ;
        RECT -59.325 174.595 -58.995 174.925 ;
        RECT -59.325 173.235 -58.995 173.565 ;
        RECT -59.325 171.875 -58.995 172.205 ;
        RECT -59.325 170.515 -58.995 170.845 ;
        RECT -59.325 169.155 -58.995 169.485 ;
        RECT -59.325 167.795 -58.995 168.125 ;
        RECT -59.325 166.435 -58.995 166.765 ;
        RECT -59.325 165.075 -58.995 165.405 ;
        RECT -59.325 163.715 -58.995 164.045 ;
        RECT -59.325 162.355 -58.995 162.685 ;
        RECT -59.325 160.995 -58.995 161.325 ;
        RECT -59.325 159.635 -58.995 159.965 ;
        RECT -59.325 158.275 -58.995 158.605 ;
        RECT -59.325 156.915 -58.995 157.245 ;
        RECT -59.325 155.555 -58.995 155.885 ;
        RECT -59.325 154.195 -58.995 154.525 ;
        RECT -59.325 152.835 -58.995 153.165 ;
        RECT -59.325 151.475 -58.995 151.805 ;
        RECT -59.325 150.115 -58.995 150.445 ;
        RECT -59.325 148.755 -58.995 149.085 ;
        RECT -59.325 147.395 -58.995 147.725 ;
        RECT -59.325 146.035 -58.995 146.365 ;
        RECT -59.325 144.675 -58.995 145.005 ;
        RECT -59.325 143.315 -58.995 143.645 ;
        RECT -59.325 141.955 -58.995 142.285 ;
        RECT -59.325 140.595 -58.995 140.925 ;
        RECT -59.325 139.235 -58.995 139.565 ;
        RECT -59.325 136.42 -58.995 136.75 ;
        RECT -59.325 134.245 -58.995 134.575 ;
        RECT -59.325 133.395 -58.995 133.725 ;
        RECT -59.325 131.085 -58.995 131.415 ;
        RECT -59.325 130.235 -58.995 130.565 ;
        RECT -59.325 127.925 -58.995 128.255 ;
        RECT -59.325 127.075 -58.995 127.405 ;
        RECT -59.325 124.765 -58.995 125.095 ;
        RECT -59.325 123.915 -58.995 124.245 ;
        RECT -59.325 121.605 -58.995 121.935 ;
        RECT -59.325 120.755 -58.995 121.085 ;
        RECT -59.325 118.445 -58.995 118.775 ;
        RECT -59.325 117.595 -58.995 117.925 ;
        RECT -59.325 115.285 -58.995 115.615 ;
        RECT -59.325 114.435 -58.995 114.765 ;
        RECT -59.325 112.125 -58.995 112.455 ;
        RECT -59.325 111.275 -58.995 111.605 ;
        RECT -59.325 108.965 -58.995 109.295 ;
        RECT -59.325 108.115 -58.995 108.445 ;
        RECT -59.325 105.805 -58.995 106.135 ;
        RECT -59.325 104.955 -58.995 105.285 ;
        RECT -59.325 102.645 -58.995 102.975 ;
        RECT -59.325 101.795 -58.995 102.125 ;
        RECT -59.325 99.62 -58.995 99.95 ;
        RECT -59.325 97.075 -58.995 97.405 ;
        RECT -59.325 95.715 -58.995 96.045 ;
        RECT -59.325 94.355 -58.995 94.685 ;
        RECT -59.325 92.995 -58.995 93.325 ;
        RECT -59.325 91.635 -58.995 91.965 ;
        RECT -59.325 90.275 -58.995 90.605 ;
        RECT -59.325 88.915 -58.995 89.245 ;
        RECT -59.32 87.56 -59 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -59.325 -2.205 -58.995 -1.875 ;
        RECT -59.325 -3.565 -58.995 -3.235 ;
        RECT -59.325 -4.925 -58.995 -4.595 ;
        RECT -59.325 -6.285 -58.995 -5.955 ;
        RECT -59.325 -7.645 -58.995 -7.315 ;
        RECT -59.325 -9.005 -58.995 -8.675 ;
        RECT -59.325 -10.365 -58.995 -10.035 ;
        RECT -59.325 -11.725 -58.995 -11.395 ;
        RECT -59.325 -13.085 -58.995 -12.755 ;
        RECT -59.325 -14.445 -58.995 -14.115 ;
        RECT -59.325 -15.805 -58.995 -15.475 ;
        RECT -59.325 -17.165 -58.995 -16.835 ;
        RECT -59.325 -18.525 -58.995 -18.195 ;
        RECT -59.325 -19.885 -58.995 -19.555 ;
        RECT -59.325 -21.245 -58.995 -20.915 ;
        RECT -59.325 -22.605 -58.995 -22.275 ;
        RECT -59.325 -23.965 -58.995 -23.635 ;
        RECT -59.325 -25.325 -58.995 -24.995 ;
        RECT -59.325 -26.685 -58.995 -26.355 ;
        RECT -59.325 -28.045 -58.995 -27.715 ;
        RECT -59.325 -29.405 -58.995 -29.075 ;
        RECT -59.325 -30.765 -58.995 -30.435 ;
        RECT -59.325 -32.125 -58.995 -31.795 ;
        RECT -59.325 -33.485 -58.995 -33.155 ;
        RECT -59.325 -34.845 -58.995 -34.515 ;
        RECT -59.325 -36.205 -58.995 -35.875 ;
        RECT -59.325 -37.565 -58.995 -37.235 ;
        RECT -59.325 -38.925 -58.995 -38.595 ;
        RECT -59.325 -40.285 -58.995 -39.955 ;
        RECT -59.325 -41.645 -58.995 -41.315 ;
        RECT -59.325 -43.005 -58.995 -42.675 ;
        RECT -59.325 -44.365 -58.995 -44.035 ;
        RECT -59.325 -45.725 -58.995 -45.395 ;
        RECT -59.325 -47.085 -58.995 -46.755 ;
        RECT -59.325 -48.445 -58.995 -48.115 ;
        RECT -59.325 -49.805 -58.995 -49.475 ;
        RECT -59.325 -51.165 -58.995 -50.835 ;
        RECT -59.325 -52.525 -58.995 -52.195 ;
        RECT -59.325 -53.885 -58.995 -53.555 ;
        RECT -59.325 -55.245 -58.995 -54.915 ;
        RECT -59.325 -56.605 -58.995 -56.275 ;
        RECT -59.325 -57.965 -58.995 -57.635 ;
        RECT -59.325 -59.325 -58.995 -58.995 ;
        RECT -59.325 -60.685 -58.995 -60.355 ;
        RECT -59.325 -62.045 -58.995 -61.715 ;
        RECT -59.325 -63.405 -58.995 -63.075 ;
        RECT -59.325 -64.765 -58.995 -64.435 ;
        RECT -59.325 -66.125 -58.995 -65.795 ;
        RECT -59.325 -67.485 -58.995 -67.155 ;
        RECT -59.325 -68.845 -58.995 -68.515 ;
        RECT -59.325 -70.205 -58.995 -69.875 ;
        RECT -59.325 -71.565 -58.995 -71.235 ;
        RECT -59.325 -72.925 -58.995 -72.595 ;
        RECT -59.325 -74.285 -58.995 -73.955 ;
        RECT -59.325 -75.645 -58.995 -75.315 ;
        RECT -59.325 -77.005 -58.995 -76.675 ;
        RECT -59.325 -78.365 -58.995 -78.035 ;
        RECT -59.325 -79.725 -58.995 -79.395 ;
        RECT -59.325 -81.085 -58.995 -80.755 ;
        RECT -59.325 -82.445 -58.995 -82.115 ;
        RECT -59.325 -83.805 -58.995 -83.475 ;
        RECT -59.325 -85.165 -58.995 -84.835 ;
        RECT -59.325 -86.525 -58.995 -86.195 ;
        RECT -59.325 -87.885 -58.995 -87.555 ;
        RECT -59.325 -89.245 -58.995 -88.915 ;
        RECT -59.325 -90.81 -58.995 -90.48 ;
        RECT -59.325 -91.965 -58.995 -91.635 ;
        RECT -59.325 -93.325 -58.995 -92.995 ;
        RECT -59.325 -94.685 -58.995 -94.355 ;
        RECT -59.325 -96.045 -58.995 -95.715 ;
        RECT -59.325 -97.405 -58.995 -97.075 ;
        RECT -59.325 -100.125 -58.995 -99.795 ;
        RECT -59.325 -101.35 -58.995 -101.02 ;
        RECT -59.325 -102.845 -58.995 -102.515 ;
        RECT -59.325 -104.205 -58.995 -103.875 ;
        RECT -59.325 -105.565 -58.995 -105.235 ;
        RECT -59.325 -108.285 -58.995 -107.955 ;
        RECT -59.325 -109.645 -58.995 -109.315 ;
        RECT -59.325 -113.725 -58.995 -113.395 ;
        RECT -59.325 -115.085 -58.995 -114.755 ;
        RECT -59.325 -116.445 -58.995 -116.115 ;
        RECT -59.325 -117.805 -58.995 -117.475 ;
        RECT -59.325 -119.165 -58.995 -118.835 ;
        RECT -59.325 -120.525 -58.995 -120.195 ;
        RECT -59.325 -121.885 -58.995 -121.555 ;
        RECT -59.325 -123.245 -58.995 -122.915 ;
        RECT -59.325 -124.605 -58.995 -124.275 ;
        RECT -59.325 -125.965 -58.995 -125.635 ;
        RECT -59.325 -127.325 -58.995 -126.995 ;
        RECT -59.325 -128.685 -58.995 -128.355 ;
        RECT -59.325 -130.045 -58.995 -129.715 ;
        RECT -59.325 -131.405 -58.995 -131.075 ;
        RECT -59.325 -132.765 -58.995 -132.435 ;
        RECT -59.325 -134.125 -58.995 -133.795 ;
        RECT -59.325 -135.485 -58.995 -135.155 ;
        RECT -59.325 -136.845 -58.995 -136.515 ;
        RECT -59.325 -138.205 -58.995 -137.875 ;
        RECT -59.325 -139.565 -58.995 -139.235 ;
        RECT -59.325 -140.925 -58.995 -140.595 ;
        RECT -59.325 -142.285 -58.995 -141.955 ;
        RECT -59.325 -143.645 -58.995 -143.315 ;
        RECT -59.325 -145.005 -58.995 -144.675 ;
        RECT -59.325 -146.365 -58.995 -146.035 ;
        RECT -59.325 -147.725 -58.995 -147.395 ;
        RECT -59.325 -149.085 -58.995 -148.755 ;
        RECT -59.325 -150.445 -58.995 -150.115 ;
        RECT -59.325 -151.805 -58.995 -151.475 ;
        RECT -59.325 -153.165 -58.995 -152.835 ;
        RECT -59.325 -154.525 -58.995 -154.195 ;
        RECT -59.325 -155.885 -58.995 -155.555 ;
        RECT -59.325 -157.245 -58.995 -156.915 ;
        RECT -59.325 -158.605 -58.995 -158.275 ;
        RECT -59.325 -159.965 -58.995 -159.635 ;
        RECT -59.325 -161.325 -58.995 -160.995 ;
        RECT -59.325 -162.685 -58.995 -162.355 ;
        RECT -59.325 -164.045 -58.995 -163.715 ;
        RECT -59.325 -165.405 -58.995 -165.075 ;
        RECT -59.325 -166.765 -58.995 -166.435 ;
        RECT -59.325 -168.655 -58.995 -168.325 ;
        RECT -59.325 -169.485 -58.995 -169.155 ;
        RECT -59.325 -170.845 -58.995 -170.515 ;
        RECT -59.325 -173.565 -58.995 -173.235 ;
        RECT -59.325 -174.925 -58.995 -174.595 ;
        RECT -59.325 -177.645 -58.995 -177.315 ;
        RECT -59.325 -183.29 -58.995 -182.16 ;
        RECT -59.32 -183.405 -59 -1.875 ;
    END
    PORT
      LAYER met3 ;
        RECT -57.965 244.04 -57.635 245.17 ;
        RECT -57.965 239.875 -57.635 240.205 ;
        RECT -57.965 238.515 -57.635 238.845 ;
        RECT -57.965 237.155 -57.635 237.485 ;
        RECT -57.965 235.795 -57.635 236.125 ;
        RECT -57.965 234.435 -57.635 234.765 ;
        RECT -57.965 233.075 -57.635 233.405 ;
        RECT -57.965 231.715 -57.635 232.045 ;
        RECT -57.965 230.355 -57.635 230.685 ;
        RECT -57.965 228.995 -57.635 229.325 ;
        RECT -57.965 227.635 -57.635 227.965 ;
        RECT -57.965 226.275 -57.635 226.605 ;
        RECT -57.965 224.915 -57.635 225.245 ;
        RECT -57.965 223.555 -57.635 223.885 ;
        RECT -57.965 222.195 -57.635 222.525 ;
        RECT -57.965 220.835 -57.635 221.165 ;
        RECT -57.965 219.475 -57.635 219.805 ;
        RECT -57.965 218.115 -57.635 218.445 ;
        RECT -57.965 216.755 -57.635 217.085 ;
        RECT -57.965 215.395 -57.635 215.725 ;
        RECT -57.965 214.035 -57.635 214.365 ;
        RECT -57.965 212.675 -57.635 213.005 ;
        RECT -57.965 211.315 -57.635 211.645 ;
        RECT -57.965 209.955 -57.635 210.285 ;
        RECT -57.965 208.595 -57.635 208.925 ;
        RECT -57.965 207.235 -57.635 207.565 ;
        RECT -57.965 205.875 -57.635 206.205 ;
        RECT -57.965 204.515 -57.635 204.845 ;
        RECT -57.965 203.155 -57.635 203.485 ;
        RECT -57.965 201.795 -57.635 202.125 ;
        RECT -57.965 200.435 -57.635 200.765 ;
        RECT -57.965 199.075 -57.635 199.405 ;
        RECT -57.965 197.715 -57.635 198.045 ;
        RECT -57.965 196.355 -57.635 196.685 ;
        RECT -57.965 194.995 -57.635 195.325 ;
        RECT -57.965 193.635 -57.635 193.965 ;
        RECT -57.965 192.275 -57.635 192.605 ;
        RECT -57.965 190.915 -57.635 191.245 ;
        RECT -57.965 189.555 -57.635 189.885 ;
        RECT -57.965 188.195 -57.635 188.525 ;
        RECT -57.965 186.835 -57.635 187.165 ;
        RECT -57.965 185.475 -57.635 185.805 ;
        RECT -57.965 184.115 -57.635 184.445 ;
        RECT -57.965 182.755 -57.635 183.085 ;
        RECT -57.965 181.395 -57.635 181.725 ;
        RECT -57.965 180.035 -57.635 180.365 ;
        RECT -57.965 178.675 -57.635 179.005 ;
        RECT -57.965 177.315 -57.635 177.645 ;
        RECT -57.965 175.955 -57.635 176.285 ;
        RECT -57.965 174.595 -57.635 174.925 ;
        RECT -57.965 173.235 -57.635 173.565 ;
        RECT -57.965 171.875 -57.635 172.205 ;
        RECT -57.965 170.515 -57.635 170.845 ;
        RECT -57.965 169.155 -57.635 169.485 ;
        RECT -57.965 167.795 -57.635 168.125 ;
        RECT -57.965 166.435 -57.635 166.765 ;
        RECT -57.965 165.075 -57.635 165.405 ;
        RECT -57.965 163.715 -57.635 164.045 ;
        RECT -57.965 162.355 -57.635 162.685 ;
        RECT -57.965 160.995 -57.635 161.325 ;
        RECT -57.965 159.635 -57.635 159.965 ;
        RECT -57.965 158.275 -57.635 158.605 ;
        RECT -57.965 156.915 -57.635 157.245 ;
        RECT -57.965 155.555 -57.635 155.885 ;
        RECT -57.965 154.195 -57.635 154.525 ;
        RECT -57.965 152.835 -57.635 153.165 ;
        RECT -57.965 151.475 -57.635 151.805 ;
        RECT -57.965 150.115 -57.635 150.445 ;
        RECT -57.965 148.755 -57.635 149.085 ;
        RECT -57.965 147.395 -57.635 147.725 ;
        RECT -57.965 146.035 -57.635 146.365 ;
        RECT -57.965 144.675 -57.635 145.005 ;
        RECT -57.965 143.315 -57.635 143.645 ;
        RECT -57.965 141.955 -57.635 142.285 ;
        RECT -57.965 140.595 -57.635 140.925 ;
        RECT -57.965 139.235 -57.635 139.565 ;
        RECT -57.96 138.56 -57.64 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -57.965 68.515 -57.635 68.845 ;
        RECT -57.965 67.155 -57.635 67.485 ;
        RECT -57.965 65.795 -57.635 66.125 ;
        RECT -57.965 64.435 -57.635 64.765 ;
        RECT -57.965 63.075 -57.635 63.405 ;
        RECT -57.965 61.715 -57.635 62.045 ;
        RECT -57.965 60.355 -57.635 60.685 ;
        RECT -57.965 58.995 -57.635 59.325 ;
        RECT -57.965 57.635 -57.635 57.965 ;
        RECT -57.965 56.275 -57.635 56.605 ;
        RECT -57.965 54.915 -57.635 55.245 ;
        RECT -57.965 53.555 -57.635 53.885 ;
        RECT -57.965 52.195 -57.635 52.525 ;
        RECT -57.965 50.835 -57.635 51.165 ;
        RECT -57.965 49.475 -57.635 49.805 ;
        RECT -57.965 48.115 -57.635 48.445 ;
        RECT -57.965 46.755 -57.635 47.085 ;
        RECT -57.965 45.395 -57.635 45.725 ;
        RECT -57.965 44.035 -57.635 44.365 ;
        RECT -57.965 42.675 -57.635 43.005 ;
        RECT -57.965 41.315 -57.635 41.645 ;
        RECT -57.965 39.955 -57.635 40.285 ;
        RECT -57.965 38.595 -57.635 38.925 ;
        RECT -57.965 37.235 -57.635 37.565 ;
        RECT -57.965 35.875 -57.635 36.205 ;
        RECT -57.965 34.515 -57.635 34.845 ;
        RECT -57.965 33.155 -57.635 33.485 ;
        RECT -57.965 31.795 -57.635 32.125 ;
        RECT -57.965 30.435 -57.635 30.765 ;
        RECT -57.965 29.075 -57.635 29.405 ;
        RECT -57.965 27.715 -57.635 28.045 ;
        RECT -57.965 26.355 -57.635 26.685 ;
        RECT -57.965 24.995 -57.635 25.325 ;
        RECT -57.965 23.635 -57.635 23.965 ;
        RECT -57.965 22.275 -57.635 22.605 ;
        RECT -57.965 20.915 -57.635 21.245 ;
        RECT -57.965 19.555 -57.635 19.885 ;
        RECT -57.965 18.195 -57.635 18.525 ;
        RECT -57.965 16.835 -57.635 17.165 ;
        RECT -57.965 15.475 -57.635 15.805 ;
        RECT -57.965 14.115 -57.635 14.445 ;
        RECT -57.965 12.755 -57.635 13.085 ;
        RECT -57.965 11.395 -57.635 11.725 ;
        RECT -57.965 10.035 -57.635 10.365 ;
        RECT -57.965 8.675 -57.635 9.005 ;
        RECT -57.965 7.315 -57.635 7.645 ;
        RECT -57.965 5.955 -57.635 6.285 ;
        RECT -57.965 4.595 -57.635 4.925 ;
        RECT -57.965 3.235 -57.635 3.565 ;
        RECT -57.965 1.875 -57.635 2.205 ;
        RECT -57.965 0.515 -57.635 0.845 ;
        RECT -57.965 -0.845 -57.635 -0.515 ;
        RECT -57.965 -2.205 -57.635 -1.875 ;
        RECT -57.965 -3.565 -57.635 -3.235 ;
        RECT -57.965 -4.925 -57.635 -4.595 ;
        RECT -57.965 -6.285 -57.635 -5.955 ;
        RECT -57.965 -7.645 -57.635 -7.315 ;
        RECT -57.965 -9.005 -57.635 -8.675 ;
        RECT -57.965 -10.365 -57.635 -10.035 ;
        RECT -57.965 -11.725 -57.635 -11.395 ;
        RECT -57.965 -13.085 -57.635 -12.755 ;
        RECT -57.965 -14.445 -57.635 -14.115 ;
        RECT -57.965 -15.805 -57.635 -15.475 ;
        RECT -57.965 -17.165 -57.635 -16.835 ;
        RECT -57.965 -18.525 -57.635 -18.195 ;
        RECT -57.965 -19.885 -57.635 -19.555 ;
        RECT -57.965 -21.245 -57.635 -20.915 ;
        RECT -57.965 -22.605 -57.635 -22.275 ;
        RECT -57.965 -23.965 -57.635 -23.635 ;
        RECT -57.965 -25.325 -57.635 -24.995 ;
        RECT -57.965 -28.045 -57.635 -27.715 ;
        RECT -57.965 -29.405 -57.635 -29.075 ;
        RECT -57.965 -30.765 -57.635 -30.435 ;
        RECT -57.965 -32.125 -57.635 -31.795 ;
        RECT -57.965 -33.485 -57.635 -33.155 ;
        RECT -57.965 -34.845 -57.635 -34.515 ;
        RECT -57.965 -36.205 -57.635 -35.875 ;
        RECT -57.965 -37.565 -57.635 -37.235 ;
        RECT -57.965 -38.925 -57.635 -38.595 ;
        RECT -57.965 -40.285 -57.635 -39.955 ;
        RECT -57.965 -41.645 -57.635 -41.315 ;
        RECT -57.965 -43.005 -57.635 -42.675 ;
        RECT -57.965 -44.365 -57.635 -44.035 ;
        RECT -57.965 -45.725 -57.635 -45.395 ;
        RECT -57.965 -47.085 -57.635 -46.755 ;
        RECT -57.965 -48.445 -57.635 -48.115 ;
        RECT -57.965 -49.805 -57.635 -49.475 ;
        RECT -57.965 -51.165 -57.635 -50.835 ;
        RECT -57.965 -52.525 -57.635 -52.195 ;
        RECT -57.965 -53.885 -57.635 -53.555 ;
        RECT -57.965 -55.245 -57.635 -54.915 ;
        RECT -57.965 -56.605 -57.635 -56.275 ;
        RECT -57.965 -57.965 -57.635 -57.635 ;
        RECT -57.965 -59.325 -57.635 -58.995 ;
        RECT -57.965 -60.685 -57.635 -60.355 ;
        RECT -57.965 -62.045 -57.635 -61.715 ;
        RECT -57.965 -63.405 -57.635 -63.075 ;
        RECT -57.965 -64.765 -57.635 -64.435 ;
        RECT -57.965 -66.125 -57.635 -65.795 ;
        RECT -57.965 -67.485 -57.635 -67.155 ;
        RECT -57.965 -68.845 -57.635 -68.515 ;
        RECT -57.965 -70.205 -57.635 -69.875 ;
        RECT -57.965 -71.565 -57.635 -71.235 ;
        RECT -57.965 -72.925 -57.635 -72.595 ;
        RECT -57.965 -74.285 -57.635 -73.955 ;
        RECT -57.965 -75.645 -57.635 -75.315 ;
        RECT -57.965 -77.005 -57.635 -76.675 ;
        RECT -57.965 -78.365 -57.635 -78.035 ;
        RECT -57.965 -79.725 -57.635 -79.395 ;
        RECT -57.965 -81.085 -57.635 -80.755 ;
        RECT -57.965 -82.445 -57.635 -82.115 ;
        RECT -57.965 -83.805 -57.635 -83.475 ;
        RECT -57.965 -85.165 -57.635 -84.835 ;
        RECT -57.965 -86.525 -57.635 -86.195 ;
        RECT -57.965 -87.885 -57.635 -87.555 ;
        RECT -57.965 -89.245 -57.635 -88.915 ;
        RECT -57.965 -90.81 -57.635 -90.48 ;
        RECT -57.965 -91.965 -57.635 -91.635 ;
        RECT -57.965 -93.325 -57.635 -92.995 ;
        RECT -57.965 -94.685 -57.635 -94.355 ;
        RECT -57.965 -96.045 -57.635 -95.715 ;
        RECT -57.965 -97.405 -57.635 -97.075 ;
        RECT -57.965 -100.125 -57.635 -99.795 ;
        RECT -57.965 -101.35 -57.635 -101.02 ;
        RECT -57.965 -102.845 -57.635 -102.515 ;
        RECT -57.965 -104.205 -57.635 -103.875 ;
        RECT -57.965 -105.565 -57.635 -105.235 ;
        RECT -57.965 -108.285 -57.635 -107.955 ;
        RECT -57.965 -109.645 -57.635 -109.315 ;
        RECT -57.965 -112.365 -57.635 -112.035 ;
        RECT -57.965 -115.085 -57.635 -114.755 ;
        RECT -57.965 -116.445 -57.635 -116.115 ;
        RECT -57.965 -117.805 -57.635 -117.475 ;
        RECT -57.965 -119.165 -57.635 -118.835 ;
        RECT -57.965 -120.525 -57.635 -120.195 ;
        RECT -57.965 -121.885 -57.635 -121.555 ;
        RECT -57.965 -123.245 -57.635 -122.915 ;
        RECT -57.965 -124.605 -57.635 -124.275 ;
        RECT -57.965 -125.965 -57.635 -125.635 ;
        RECT -57.965 -127.325 -57.635 -126.995 ;
        RECT -57.965 -128.685 -57.635 -128.355 ;
        RECT -57.965 -130.045 -57.635 -129.715 ;
        RECT -57.965 -131.405 -57.635 -131.075 ;
        RECT -57.965 -132.765 -57.635 -132.435 ;
        RECT -57.965 -134.125 -57.635 -133.795 ;
        RECT -57.965 -135.485 -57.635 -135.155 ;
        RECT -57.965 -136.845 -57.635 -136.515 ;
        RECT -57.965 -138.205 -57.635 -137.875 ;
        RECT -57.965 -139.565 -57.635 -139.235 ;
        RECT -57.965 -140.925 -57.635 -140.595 ;
        RECT -57.965 -142.285 -57.635 -141.955 ;
        RECT -57.965 -143.645 -57.635 -143.315 ;
        RECT -57.965 -145.005 -57.635 -144.675 ;
        RECT -57.965 -146.365 -57.635 -146.035 ;
        RECT -57.965 -147.725 -57.635 -147.395 ;
        RECT -57.965 -149.085 -57.635 -148.755 ;
        RECT -57.965 -150.445 -57.635 -150.115 ;
        RECT -57.965 -151.805 -57.635 -151.475 ;
        RECT -57.965 -153.165 -57.635 -152.835 ;
        RECT -57.965 -154.525 -57.635 -154.195 ;
        RECT -57.965 -155.885 -57.635 -155.555 ;
        RECT -57.965 -157.245 -57.635 -156.915 ;
        RECT -57.965 -158.605 -57.635 -158.275 ;
        RECT -57.965 -159.965 -57.635 -159.635 ;
        RECT -57.965 -161.325 -57.635 -160.995 ;
        RECT -57.965 -162.685 -57.635 -162.355 ;
        RECT -57.965 -164.045 -57.635 -163.715 ;
        RECT -57.965 -165.405 -57.635 -165.075 ;
        RECT -57.965 -166.765 -57.635 -166.435 ;
        RECT -57.965 -168.655 -57.635 -168.325 ;
        RECT -57.965 -169.485 -57.635 -169.155 ;
        RECT -57.965 -170.845 -57.635 -170.515 ;
        RECT -57.965 -173.565 -57.635 -173.235 ;
        RECT -57.965 -174.925 -57.635 -174.595 ;
        RECT -57.965 -177.645 -57.635 -177.315 ;
        RECT -57.965 -183.29 -57.635 -182.16 ;
        RECT -57.96 -183.405 -57.64 98.08 ;
        RECT -57.965 97.075 -57.635 97.405 ;
        RECT -57.965 95.715 -57.635 96.045 ;
        RECT -57.965 94.355 -57.635 94.685 ;
        RECT -57.965 92.995 -57.635 93.325 ;
        RECT -57.965 88.915 -57.635 89.245 ;
        RECT -57.965 84.835 -57.635 85.165 ;
        RECT -57.965 83.475 -57.635 83.805 ;
        RECT -57.965 82.115 -57.635 82.445 ;
        RECT -57.965 80.755 -57.635 81.085 ;
        RECT -57.965 79.395 -57.635 79.725 ;
        RECT -57.965 78.035 -57.635 78.365 ;
        RECT -57.965 76.675 -57.635 77.005 ;
        RECT -57.965 75.315 -57.635 75.645 ;
        RECT -57.965 73.955 -57.635 74.285 ;
        RECT -57.965 72.595 -57.635 72.925 ;
        RECT -57.965 71.235 -57.635 71.565 ;
        RECT -57.965 69.875 -57.635 70.205 ;
    END
    PORT
      LAYER met3 ;
        RECT -66.125 244.04 -65.795 245.17 ;
        RECT -66.125 239.875 -65.795 240.205 ;
        RECT -66.125 238.515 -65.795 238.845 ;
        RECT -66.125 237.155 -65.795 237.485 ;
        RECT -66.125 235.795 -65.795 236.125 ;
        RECT -66.125 234.435 -65.795 234.765 ;
        RECT -66.125 233.075 -65.795 233.405 ;
        RECT -66.125 231.715 -65.795 232.045 ;
        RECT -66.125 230.355 -65.795 230.685 ;
        RECT -66.125 228.995 -65.795 229.325 ;
        RECT -66.125 227.635 -65.795 227.965 ;
        RECT -66.125 226.275 -65.795 226.605 ;
        RECT -66.125 224.915 -65.795 225.245 ;
        RECT -66.125 223.555 -65.795 223.885 ;
        RECT -66.125 222.195 -65.795 222.525 ;
        RECT -66.125 220.835 -65.795 221.165 ;
        RECT -66.125 219.475 -65.795 219.805 ;
        RECT -66.125 218.115 -65.795 218.445 ;
        RECT -66.125 216.755 -65.795 217.085 ;
        RECT -66.125 215.395 -65.795 215.725 ;
        RECT -66.125 214.035 -65.795 214.365 ;
        RECT -66.125 212.675 -65.795 213.005 ;
        RECT -66.125 211.315 -65.795 211.645 ;
        RECT -66.125 209.955 -65.795 210.285 ;
        RECT -66.125 208.595 -65.795 208.925 ;
        RECT -66.125 207.235 -65.795 207.565 ;
        RECT -66.125 205.875 -65.795 206.205 ;
        RECT -66.125 204.515 -65.795 204.845 ;
        RECT -66.125 203.155 -65.795 203.485 ;
        RECT -66.125 201.795 -65.795 202.125 ;
        RECT -66.125 200.435 -65.795 200.765 ;
        RECT -66.125 199.075 -65.795 199.405 ;
        RECT -66.125 197.715 -65.795 198.045 ;
        RECT -66.125 196.355 -65.795 196.685 ;
        RECT -66.125 194.995 -65.795 195.325 ;
        RECT -66.125 193.635 -65.795 193.965 ;
        RECT -66.125 192.275 -65.795 192.605 ;
        RECT -66.125 190.915 -65.795 191.245 ;
        RECT -66.125 189.555 -65.795 189.885 ;
        RECT -66.125 188.195 -65.795 188.525 ;
        RECT -66.125 186.835 -65.795 187.165 ;
        RECT -66.125 185.475 -65.795 185.805 ;
        RECT -66.125 184.115 -65.795 184.445 ;
        RECT -66.125 182.755 -65.795 183.085 ;
        RECT -66.125 181.395 -65.795 181.725 ;
        RECT -66.125 180.035 -65.795 180.365 ;
        RECT -66.125 178.675 -65.795 179.005 ;
        RECT -66.125 177.315 -65.795 177.645 ;
        RECT -66.125 175.955 -65.795 176.285 ;
        RECT -66.125 174.595 -65.795 174.925 ;
        RECT -66.125 173.235 -65.795 173.565 ;
        RECT -66.125 171.875 -65.795 172.205 ;
        RECT -66.125 170.515 -65.795 170.845 ;
        RECT -66.125 169.155 -65.795 169.485 ;
        RECT -66.125 167.795 -65.795 168.125 ;
        RECT -66.125 166.435 -65.795 166.765 ;
        RECT -66.125 165.075 -65.795 165.405 ;
        RECT -66.125 163.715 -65.795 164.045 ;
        RECT -66.125 162.355 -65.795 162.685 ;
        RECT -66.125 160.995 -65.795 161.325 ;
        RECT -66.125 159.635 -65.795 159.965 ;
        RECT -66.125 158.275 -65.795 158.605 ;
        RECT -66.125 156.915 -65.795 157.245 ;
        RECT -66.125 155.555 -65.795 155.885 ;
        RECT -66.125 154.195 -65.795 154.525 ;
        RECT -66.125 152.835 -65.795 153.165 ;
        RECT -66.125 151.475 -65.795 151.805 ;
        RECT -66.125 150.115 -65.795 150.445 ;
        RECT -66.125 148.755 -65.795 149.085 ;
        RECT -66.125 147.395 -65.795 147.725 ;
        RECT -66.125 146.035 -65.795 146.365 ;
        RECT -66.125 144.675 -65.795 145.005 ;
        RECT -66.125 143.315 -65.795 143.645 ;
        RECT -66.125 141.955 -65.795 142.285 ;
        RECT -66.125 140.595 -65.795 140.925 ;
        RECT -66.125 139.235 -65.795 139.565 ;
        RECT -66.125 137.875 -65.795 138.205 ;
        RECT -66.125 136.515 -65.795 136.845 ;
        RECT -66.125 135.155 -65.795 135.485 ;
        RECT -66.125 133.795 -65.795 134.125 ;
        RECT -66.125 132.435 -65.795 132.765 ;
        RECT -66.125 131.075 -65.795 131.405 ;
        RECT -66.125 129.715 -65.795 130.045 ;
        RECT -66.125 128.355 -65.795 128.685 ;
        RECT -66.125 126.995 -65.795 127.325 ;
        RECT -66.125 125.635 -65.795 125.965 ;
        RECT -66.125 124.275 -65.795 124.605 ;
        RECT -66.125 122.915 -65.795 123.245 ;
        RECT -66.125 121.555 -65.795 121.885 ;
        RECT -66.125 120.195 -65.795 120.525 ;
        RECT -66.125 118.835 -65.795 119.165 ;
        RECT -66.125 117.475 -65.795 117.805 ;
        RECT -66.125 116.115 -65.795 116.445 ;
        RECT -66.125 114.755 -65.795 115.085 ;
        RECT -66.125 113.395 -65.795 113.725 ;
        RECT -66.125 112.035 -65.795 112.365 ;
        RECT -66.125 110.675 -65.795 111.005 ;
        RECT -66.125 109.315 -65.795 109.645 ;
        RECT -66.125 107.955 -65.795 108.285 ;
        RECT -66.125 106.595 -65.795 106.925 ;
        RECT -66.125 105.235 -65.795 105.565 ;
        RECT -66.125 103.875 -65.795 104.205 ;
        RECT -66.125 102.515 -65.795 102.845 ;
        RECT -66.125 101.155 -65.795 101.485 ;
        RECT -66.125 99.795 -65.795 100.125 ;
        RECT -66.125 98.435 -65.795 98.765 ;
        RECT -66.125 97.075 -65.795 97.405 ;
        RECT -66.125 95.715 -65.795 96.045 ;
        RECT -66.125 94.355 -65.795 94.685 ;
        RECT -66.125 92.995 -65.795 93.325 ;
        RECT -66.125 91.635 -65.795 91.965 ;
        RECT -66.125 90.275 -65.795 90.605 ;
        RECT -66.125 88.915 -65.795 89.245 ;
        RECT -66.125 87.555 -65.795 87.885 ;
        RECT -66.125 86.195 -65.795 86.525 ;
        RECT -66.125 84.835 -65.795 85.165 ;
        RECT -66.125 83.475 -65.795 83.805 ;
        RECT -66.125 82.115 -65.795 82.445 ;
        RECT -66.125 80.755 -65.795 81.085 ;
        RECT -66.125 79.395 -65.795 79.725 ;
        RECT -66.125 78.035 -65.795 78.365 ;
        RECT -66.125 76.675 -65.795 77.005 ;
        RECT -66.125 75.315 -65.795 75.645 ;
        RECT -66.125 73.955 -65.795 74.285 ;
        RECT -66.125 72.595 -65.795 72.925 ;
        RECT -66.125 71.235 -65.795 71.565 ;
        RECT -66.125 69.875 -65.795 70.205 ;
        RECT -66.125 68.515 -65.795 68.845 ;
        RECT -66.125 67.155 -65.795 67.485 ;
        RECT -66.125 65.795 -65.795 66.125 ;
        RECT -66.125 64.435 -65.795 64.765 ;
        RECT -66.125 63.075 -65.795 63.405 ;
        RECT -66.125 61.715 -65.795 62.045 ;
        RECT -66.125 60.355 -65.795 60.685 ;
        RECT -66.125 58.995 -65.795 59.325 ;
        RECT -66.125 57.635 -65.795 57.965 ;
        RECT -66.125 56.275 -65.795 56.605 ;
        RECT -66.125 54.915 -65.795 55.245 ;
        RECT -66.125 53.555 -65.795 53.885 ;
        RECT -66.125 52.195 -65.795 52.525 ;
        RECT -66.125 50.835 -65.795 51.165 ;
        RECT -66.125 49.475 -65.795 49.805 ;
        RECT -66.125 48.115 -65.795 48.445 ;
        RECT -66.125 46.755 -65.795 47.085 ;
        RECT -66.125 45.395 -65.795 45.725 ;
        RECT -66.125 44.035 -65.795 44.365 ;
        RECT -66.125 42.675 -65.795 43.005 ;
        RECT -66.125 41.315 -65.795 41.645 ;
        RECT -66.125 39.955 -65.795 40.285 ;
        RECT -66.125 38.595 -65.795 38.925 ;
        RECT -66.125 37.235 -65.795 37.565 ;
        RECT -66.125 35.875 -65.795 36.205 ;
        RECT -66.125 34.515 -65.795 34.845 ;
        RECT -66.125 33.155 -65.795 33.485 ;
        RECT -66.125 31.795 -65.795 32.125 ;
        RECT -66.125 30.435 -65.795 30.765 ;
        RECT -66.125 29.075 -65.795 29.405 ;
        RECT -66.125 27.715 -65.795 28.045 ;
        RECT -66.125 26.355 -65.795 26.685 ;
        RECT -66.125 24.995 -65.795 25.325 ;
        RECT -66.125 23.635 -65.795 23.965 ;
        RECT -66.125 22.275 -65.795 22.605 ;
        RECT -66.125 20.915 -65.795 21.245 ;
        RECT -66.125 19.555 -65.795 19.885 ;
        RECT -66.125 18.195 -65.795 18.525 ;
        RECT -66.125 16.835 -65.795 17.165 ;
        RECT -66.125 15.475 -65.795 15.805 ;
        RECT -66.125 14.115 -65.795 14.445 ;
        RECT -66.125 12.755 -65.795 13.085 ;
        RECT -66.125 11.395 -65.795 11.725 ;
        RECT -66.125 10.035 -65.795 10.365 ;
        RECT -66.125 8.675 -65.795 9.005 ;
        RECT -66.125 7.315 -65.795 7.645 ;
        RECT -66.125 5.955 -65.795 6.285 ;
        RECT -66.125 4.595 -65.795 4.925 ;
        RECT -66.125 3.235 -65.795 3.565 ;
        RECT -66.125 1.875 -65.795 2.205 ;
        RECT -66.125 0.515 -65.795 0.845 ;
        RECT -66.125 -0.845 -65.795 -0.515 ;
        RECT -66.125 -2.205 -65.795 -1.875 ;
        RECT -66.125 -3.565 -65.795 -3.235 ;
        RECT -66.125 -4.925 -65.795 -4.595 ;
        RECT -66.125 -6.285 -65.795 -5.955 ;
        RECT -66.125 -7.645 -65.795 -7.315 ;
        RECT -66.125 -9.005 -65.795 -8.675 ;
        RECT -66.125 -10.365 -65.795 -10.035 ;
        RECT -66.125 -11.725 -65.795 -11.395 ;
        RECT -66.125 -13.085 -65.795 -12.755 ;
        RECT -66.125 -14.445 -65.795 -14.115 ;
        RECT -66.125 -15.805 -65.795 -15.475 ;
        RECT -66.125 -17.165 -65.795 -16.835 ;
        RECT -66.125 -18.525 -65.795 -18.195 ;
        RECT -66.125 -19.885 -65.795 -19.555 ;
        RECT -66.125 -21.245 -65.795 -20.915 ;
        RECT -66.125 -22.605 -65.795 -22.275 ;
        RECT -66.125 -23.965 -65.795 -23.635 ;
        RECT -66.125 -25.325 -65.795 -24.995 ;
        RECT -66.125 -26.685 -65.795 -26.355 ;
        RECT -66.125 -28.045 -65.795 -27.715 ;
        RECT -66.125 -29.405 -65.795 -29.075 ;
        RECT -66.125 -30.765 -65.795 -30.435 ;
        RECT -66.125 -32.125 -65.795 -31.795 ;
        RECT -66.125 -33.485 -65.795 -33.155 ;
        RECT -66.125 -34.845 -65.795 -34.515 ;
        RECT -66.125 -36.205 -65.795 -35.875 ;
        RECT -66.125 -37.565 -65.795 -37.235 ;
        RECT -66.125 -38.925 -65.795 -38.595 ;
        RECT -66.125 -40.285 -65.795 -39.955 ;
        RECT -66.125 -41.645 -65.795 -41.315 ;
        RECT -66.125 -43.005 -65.795 -42.675 ;
        RECT -66.125 -44.365 -65.795 -44.035 ;
        RECT -66.125 -45.725 -65.795 -45.395 ;
        RECT -66.125 -47.085 -65.795 -46.755 ;
        RECT -66.125 -48.445 -65.795 -48.115 ;
        RECT -66.125 -49.805 -65.795 -49.475 ;
        RECT -66.125 -51.165 -65.795 -50.835 ;
        RECT -66.125 -52.525 -65.795 -52.195 ;
        RECT -66.125 -53.885 -65.795 -53.555 ;
        RECT -66.125 -55.245 -65.795 -54.915 ;
        RECT -66.125 -56.605 -65.795 -56.275 ;
        RECT -66.125 -57.965 -65.795 -57.635 ;
        RECT -66.125 -59.325 -65.795 -58.995 ;
        RECT -66.125 -60.685 -65.795 -60.355 ;
        RECT -66.125 -62.045 -65.795 -61.715 ;
        RECT -66.125 -63.405 -65.795 -63.075 ;
        RECT -66.125 -64.765 -65.795 -64.435 ;
        RECT -66.125 -66.125 -65.795 -65.795 ;
        RECT -66.125 -67.485 -65.795 -67.155 ;
        RECT -66.125 -68.845 -65.795 -68.515 ;
        RECT -66.125 -70.205 -65.795 -69.875 ;
        RECT -66.125 -71.565 -65.795 -71.235 ;
        RECT -66.125 -72.925 -65.795 -72.595 ;
        RECT -66.125 -74.285 -65.795 -73.955 ;
        RECT -66.125 -75.645 -65.795 -75.315 ;
        RECT -66.125 -77.005 -65.795 -76.675 ;
        RECT -66.125 -78.365 -65.795 -78.035 ;
        RECT -66.125 -79.725 -65.795 -79.395 ;
        RECT -66.125 -81.085 -65.795 -80.755 ;
        RECT -66.125 -82.445 -65.795 -82.115 ;
        RECT -66.125 -83.805 -65.795 -83.475 ;
        RECT -66.125 -85.165 -65.795 -84.835 ;
        RECT -66.125 -86.525 -65.795 -86.195 ;
        RECT -66.125 -87.885 -65.795 -87.555 ;
        RECT -66.125 -89.245 -65.795 -88.915 ;
        RECT -66.125 -90.605 -65.795 -90.275 ;
        RECT -66.125 -91.965 -65.795 -91.635 ;
        RECT -66.125 -93.325 -65.795 -92.995 ;
        RECT -66.125 -94.685 -65.795 -94.355 ;
        RECT -66.125 -96.045 -65.795 -95.715 ;
        RECT -66.125 -97.405 -65.795 -97.075 ;
        RECT -66.125 -98.765 -65.795 -98.435 ;
        RECT -66.125 -100.125 -65.795 -99.795 ;
        RECT -66.125 -101.485 -65.795 -101.155 ;
        RECT -66.125 -102.845 -65.795 -102.515 ;
        RECT -66.125 -104.205 -65.795 -103.875 ;
        RECT -66.125 -105.565 -65.795 -105.235 ;
        RECT -66.125 -106.925 -65.795 -106.595 ;
        RECT -66.125 -108.285 -65.795 -107.955 ;
        RECT -66.125 -109.645 -65.795 -109.315 ;
        RECT -66.125 -111.005 -65.795 -110.675 ;
        RECT -66.125 -112.365 -65.795 -112.035 ;
        RECT -66.125 -113.725 -65.795 -113.395 ;
        RECT -66.125 -115.085 -65.795 -114.755 ;
        RECT -66.125 -116.445 -65.795 -116.115 ;
        RECT -66.125 -117.805 -65.795 -117.475 ;
        RECT -66.125 -119.165 -65.795 -118.835 ;
        RECT -66.125 -120.525 -65.795 -120.195 ;
        RECT -66.125 -121.885 -65.795 -121.555 ;
        RECT -66.125 -123.245 -65.795 -122.915 ;
        RECT -66.125 -124.605 -65.795 -124.275 ;
        RECT -66.125 -125.965 -65.795 -125.635 ;
        RECT -66.125 -127.325 -65.795 -126.995 ;
        RECT -66.125 -128.685 -65.795 -128.355 ;
        RECT -66.125 -130.045 -65.795 -129.715 ;
        RECT -66.125 -131.405 -65.795 -131.075 ;
        RECT -66.125 -132.765 -65.795 -132.435 ;
        RECT -66.125 -134.125 -65.795 -133.795 ;
        RECT -66.125 -135.485 -65.795 -135.155 ;
        RECT -66.125 -136.845 -65.795 -136.515 ;
        RECT -66.125 -138.205 -65.795 -137.875 ;
        RECT -66.125 -139.565 -65.795 -139.235 ;
        RECT -66.125 -140.925 -65.795 -140.595 ;
        RECT -66.125 -142.285 -65.795 -141.955 ;
        RECT -66.125 -143.645 -65.795 -143.315 ;
        RECT -66.125 -145.005 -65.795 -144.675 ;
        RECT -66.125 -146.365 -65.795 -146.035 ;
        RECT -66.125 -147.725 -65.795 -147.395 ;
        RECT -66.125 -149.085 -65.795 -148.755 ;
        RECT -66.125 -150.445 -65.795 -150.115 ;
        RECT -66.125 -151.805 -65.795 -151.475 ;
        RECT -66.125 -153.165 -65.795 -152.835 ;
        RECT -66.125 -154.525 -65.795 -154.195 ;
        RECT -66.125 -155.885 -65.795 -155.555 ;
        RECT -66.125 -157.245 -65.795 -156.915 ;
        RECT -66.125 -158.605 -65.795 -158.275 ;
        RECT -66.125 -159.965 -65.795 -159.635 ;
        RECT -66.125 -161.325 -65.795 -160.995 ;
        RECT -66.125 -162.685 -65.795 -162.355 ;
        RECT -66.125 -164.045 -65.795 -163.715 ;
        RECT -66.125 -165.405 -65.795 -165.075 ;
        RECT -66.125 -166.765 -65.795 -166.435 ;
        RECT -66.125 -169.485 -65.795 -169.155 ;
        RECT -66.125 -170.845 -65.795 -170.515 ;
        RECT -66.125 -174.925 -65.795 -174.595 ;
        RECT -66.125 -177.645 -65.795 -177.315 ;
        RECT -66.125 -183.29 -65.795 -182.16 ;
        RECT -66.12 -183.405 -65.8 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -64.765 244.04 -64.435 245.17 ;
        RECT -64.765 239.875 -64.435 240.205 ;
        RECT -64.765 238.515 -64.435 238.845 ;
        RECT -64.765 237.155 -64.435 237.485 ;
        RECT -64.765 235.795 -64.435 236.125 ;
        RECT -64.765 234.435 -64.435 234.765 ;
        RECT -64.765 233.075 -64.435 233.405 ;
        RECT -64.765 231.715 -64.435 232.045 ;
        RECT -64.765 230.355 -64.435 230.685 ;
        RECT -64.765 228.995 -64.435 229.325 ;
        RECT -64.765 227.635 -64.435 227.965 ;
        RECT -64.765 226.275 -64.435 226.605 ;
        RECT -64.765 224.915 -64.435 225.245 ;
        RECT -64.765 223.555 -64.435 223.885 ;
        RECT -64.765 222.195 -64.435 222.525 ;
        RECT -64.765 220.835 -64.435 221.165 ;
        RECT -64.765 219.475 -64.435 219.805 ;
        RECT -64.765 218.115 -64.435 218.445 ;
        RECT -64.765 216.755 -64.435 217.085 ;
        RECT -64.765 215.395 -64.435 215.725 ;
        RECT -64.765 214.035 -64.435 214.365 ;
        RECT -64.765 212.675 -64.435 213.005 ;
        RECT -64.765 211.315 -64.435 211.645 ;
        RECT -64.765 209.955 -64.435 210.285 ;
        RECT -64.765 208.595 -64.435 208.925 ;
        RECT -64.765 207.235 -64.435 207.565 ;
        RECT -64.765 205.875 -64.435 206.205 ;
        RECT -64.765 204.515 -64.435 204.845 ;
        RECT -64.765 203.155 -64.435 203.485 ;
        RECT -64.765 201.795 -64.435 202.125 ;
        RECT -64.765 200.435 -64.435 200.765 ;
        RECT -64.765 199.075 -64.435 199.405 ;
        RECT -64.765 197.715 -64.435 198.045 ;
        RECT -64.765 196.355 -64.435 196.685 ;
        RECT -64.765 194.995 -64.435 195.325 ;
        RECT -64.765 193.635 -64.435 193.965 ;
        RECT -64.765 192.275 -64.435 192.605 ;
        RECT -64.765 190.915 -64.435 191.245 ;
        RECT -64.765 189.555 -64.435 189.885 ;
        RECT -64.765 188.195 -64.435 188.525 ;
        RECT -64.765 186.835 -64.435 187.165 ;
        RECT -64.765 185.475 -64.435 185.805 ;
        RECT -64.765 184.115 -64.435 184.445 ;
        RECT -64.765 182.755 -64.435 183.085 ;
        RECT -64.765 181.395 -64.435 181.725 ;
        RECT -64.765 180.035 -64.435 180.365 ;
        RECT -64.765 178.675 -64.435 179.005 ;
        RECT -64.765 177.315 -64.435 177.645 ;
        RECT -64.765 175.955 -64.435 176.285 ;
        RECT -64.765 174.595 -64.435 174.925 ;
        RECT -64.765 173.235 -64.435 173.565 ;
        RECT -64.765 171.875 -64.435 172.205 ;
        RECT -64.765 170.515 -64.435 170.845 ;
        RECT -64.765 169.155 -64.435 169.485 ;
        RECT -64.765 167.795 -64.435 168.125 ;
        RECT -64.765 166.435 -64.435 166.765 ;
        RECT -64.765 165.075 -64.435 165.405 ;
        RECT -64.765 163.715 -64.435 164.045 ;
        RECT -64.765 162.355 -64.435 162.685 ;
        RECT -64.765 160.995 -64.435 161.325 ;
        RECT -64.765 159.635 -64.435 159.965 ;
        RECT -64.765 158.275 -64.435 158.605 ;
        RECT -64.765 156.915 -64.435 157.245 ;
        RECT -64.765 155.555 -64.435 155.885 ;
        RECT -64.765 154.195 -64.435 154.525 ;
        RECT -64.765 152.835 -64.435 153.165 ;
        RECT -64.765 151.475 -64.435 151.805 ;
        RECT -64.765 150.115 -64.435 150.445 ;
        RECT -64.765 148.755 -64.435 149.085 ;
        RECT -64.765 147.395 -64.435 147.725 ;
        RECT -64.765 146.035 -64.435 146.365 ;
        RECT -64.765 144.675 -64.435 145.005 ;
        RECT -64.765 143.315 -64.435 143.645 ;
        RECT -64.765 141.955 -64.435 142.285 ;
        RECT -64.765 140.595 -64.435 140.925 ;
        RECT -64.765 139.235 -64.435 139.565 ;
        RECT -64.765 97.075 -64.435 97.405 ;
        RECT -64.765 95.715 -64.435 96.045 ;
        RECT -64.765 94.355 -64.435 94.685 ;
        RECT -64.765 92.995 -64.435 93.325 ;
        RECT -64.765 91.635 -64.435 91.965 ;
        RECT -64.765 90.275 -64.435 90.605 ;
        RECT -64.765 88.915 -64.435 89.245 ;
        RECT -64.765 87.555 -64.435 87.885 ;
        RECT -64.765 86.195 -64.435 86.525 ;
        RECT -64.765 84.835 -64.435 85.165 ;
        RECT -64.765 83.475 -64.435 83.805 ;
        RECT -64.765 82.115 -64.435 82.445 ;
        RECT -64.765 80.755 -64.435 81.085 ;
        RECT -64.765 79.395 -64.435 79.725 ;
        RECT -64.765 78.035 -64.435 78.365 ;
        RECT -64.765 76.675 -64.435 77.005 ;
        RECT -64.765 75.315 -64.435 75.645 ;
        RECT -64.765 73.955 -64.435 74.285 ;
        RECT -64.765 72.595 -64.435 72.925 ;
        RECT -64.765 71.235 -64.435 71.565 ;
        RECT -64.765 69.875 -64.435 70.205 ;
        RECT -64.765 68.515 -64.435 68.845 ;
        RECT -64.765 67.155 -64.435 67.485 ;
        RECT -64.765 65.795 -64.435 66.125 ;
        RECT -64.765 64.435 -64.435 64.765 ;
        RECT -64.765 63.075 -64.435 63.405 ;
        RECT -64.765 61.715 -64.435 62.045 ;
        RECT -64.765 60.355 -64.435 60.685 ;
        RECT -64.765 58.995 -64.435 59.325 ;
        RECT -64.765 57.635 -64.435 57.965 ;
        RECT -64.765 56.275 -64.435 56.605 ;
        RECT -64.765 54.915 -64.435 55.245 ;
        RECT -64.765 53.555 -64.435 53.885 ;
        RECT -64.765 52.195 -64.435 52.525 ;
        RECT -64.765 50.835 -64.435 51.165 ;
        RECT -64.765 49.475 -64.435 49.805 ;
        RECT -64.765 48.115 -64.435 48.445 ;
        RECT -64.765 46.755 -64.435 47.085 ;
        RECT -64.765 45.395 -64.435 45.725 ;
        RECT -64.765 44.035 -64.435 44.365 ;
        RECT -64.765 42.675 -64.435 43.005 ;
        RECT -64.765 41.315 -64.435 41.645 ;
        RECT -64.765 39.955 -64.435 40.285 ;
        RECT -64.765 38.595 -64.435 38.925 ;
        RECT -64.765 37.235 -64.435 37.565 ;
        RECT -64.765 35.875 -64.435 36.205 ;
        RECT -64.765 34.515 -64.435 34.845 ;
        RECT -64.765 33.155 -64.435 33.485 ;
        RECT -64.765 31.795 -64.435 32.125 ;
        RECT -64.765 30.435 -64.435 30.765 ;
        RECT -64.765 29.075 -64.435 29.405 ;
        RECT -64.765 27.715 -64.435 28.045 ;
        RECT -64.765 26.355 -64.435 26.685 ;
        RECT -64.765 24.995 -64.435 25.325 ;
        RECT -64.765 23.635 -64.435 23.965 ;
        RECT -64.765 22.275 -64.435 22.605 ;
        RECT -64.765 20.915 -64.435 21.245 ;
        RECT -64.765 19.555 -64.435 19.885 ;
        RECT -64.765 18.195 -64.435 18.525 ;
        RECT -64.765 16.835 -64.435 17.165 ;
        RECT -64.765 15.475 -64.435 15.805 ;
        RECT -64.765 14.115 -64.435 14.445 ;
        RECT -64.765 12.755 -64.435 13.085 ;
        RECT -64.765 11.395 -64.435 11.725 ;
        RECT -64.765 10.035 -64.435 10.365 ;
        RECT -64.765 8.675 -64.435 9.005 ;
        RECT -64.765 7.315 -64.435 7.645 ;
        RECT -64.765 5.955 -64.435 6.285 ;
        RECT -64.765 4.595 -64.435 4.925 ;
        RECT -64.765 3.235 -64.435 3.565 ;
        RECT -64.765 1.875 -64.435 2.205 ;
        RECT -64.765 0.515 -64.435 0.845 ;
        RECT -64.765 -0.845 -64.435 -0.515 ;
        RECT -64.765 -2.205 -64.435 -1.875 ;
        RECT -64.765 -3.565 -64.435 -3.235 ;
        RECT -64.765 -4.925 -64.435 -4.595 ;
        RECT -64.765 -6.285 -64.435 -5.955 ;
        RECT -64.765 -7.645 -64.435 -7.315 ;
        RECT -64.765 -9.005 -64.435 -8.675 ;
        RECT -64.765 -10.365 -64.435 -10.035 ;
        RECT -64.765 -11.725 -64.435 -11.395 ;
        RECT -64.765 -13.085 -64.435 -12.755 ;
        RECT -64.765 -14.445 -64.435 -14.115 ;
        RECT -64.765 -15.805 -64.435 -15.475 ;
        RECT -64.765 -17.165 -64.435 -16.835 ;
        RECT -64.765 -18.525 -64.435 -18.195 ;
        RECT -64.765 -19.885 -64.435 -19.555 ;
        RECT -64.765 -21.245 -64.435 -20.915 ;
        RECT -64.765 -22.605 -64.435 -22.275 ;
        RECT -64.765 -23.965 -64.435 -23.635 ;
        RECT -64.765 -25.325 -64.435 -24.995 ;
        RECT -64.765 -26.685 -64.435 -26.355 ;
        RECT -64.765 -28.045 -64.435 -27.715 ;
        RECT -64.765 -29.405 -64.435 -29.075 ;
        RECT -64.765 -30.765 -64.435 -30.435 ;
        RECT -64.765 -32.125 -64.435 -31.795 ;
        RECT -64.765 -33.485 -64.435 -33.155 ;
        RECT -64.765 -34.845 -64.435 -34.515 ;
        RECT -64.765 -36.205 -64.435 -35.875 ;
        RECT -64.765 -37.565 -64.435 -37.235 ;
        RECT -64.765 -38.925 -64.435 -38.595 ;
        RECT -64.765 -40.285 -64.435 -39.955 ;
        RECT -64.765 -41.645 -64.435 -41.315 ;
        RECT -64.765 -43.005 -64.435 -42.675 ;
        RECT -64.765 -44.365 -64.435 -44.035 ;
        RECT -64.765 -45.725 -64.435 -45.395 ;
        RECT -64.765 -47.085 -64.435 -46.755 ;
        RECT -64.765 -48.445 -64.435 -48.115 ;
        RECT -64.765 -49.805 -64.435 -49.475 ;
        RECT -64.765 -51.165 -64.435 -50.835 ;
        RECT -64.765 -52.525 -64.435 -52.195 ;
        RECT -64.765 -53.885 -64.435 -53.555 ;
        RECT -64.765 -55.245 -64.435 -54.915 ;
        RECT -64.765 -56.605 -64.435 -56.275 ;
        RECT -64.765 -57.965 -64.435 -57.635 ;
        RECT -64.765 -59.325 -64.435 -58.995 ;
        RECT -64.765 -60.685 -64.435 -60.355 ;
        RECT -64.765 -62.045 -64.435 -61.715 ;
        RECT -64.765 -63.405 -64.435 -63.075 ;
        RECT -64.765 -64.765 -64.435 -64.435 ;
        RECT -64.765 -66.125 -64.435 -65.795 ;
        RECT -64.765 -67.485 -64.435 -67.155 ;
        RECT -64.765 -68.845 -64.435 -68.515 ;
        RECT -64.765 -70.205 -64.435 -69.875 ;
        RECT -64.765 -71.565 -64.435 -71.235 ;
        RECT -64.765 -72.925 -64.435 -72.595 ;
        RECT -64.765 -74.285 -64.435 -73.955 ;
        RECT -64.765 -75.645 -64.435 -75.315 ;
        RECT -64.765 -77.005 -64.435 -76.675 ;
        RECT -64.765 -78.365 -64.435 -78.035 ;
        RECT -64.765 -79.725 -64.435 -79.395 ;
        RECT -64.765 -81.085 -64.435 -80.755 ;
        RECT -64.765 -82.445 -64.435 -82.115 ;
        RECT -64.765 -83.805 -64.435 -83.475 ;
        RECT -64.765 -85.165 -64.435 -84.835 ;
        RECT -64.765 -86.525 -64.435 -86.195 ;
        RECT -64.765 -87.885 -64.435 -87.555 ;
        RECT -64.765 -89.245 -64.435 -88.915 ;
        RECT -64.765 -90.605 -64.435 -90.275 ;
        RECT -64.765 -91.965 -64.435 -91.635 ;
        RECT -64.765 -93.325 -64.435 -92.995 ;
        RECT -64.765 -94.685 -64.435 -94.355 ;
        RECT -64.765 -96.045 -64.435 -95.715 ;
        RECT -64.765 -97.405 -64.435 -97.075 ;
        RECT -64.765 -98.765 -64.435 -98.435 ;
        RECT -64.765 -100.125 -64.435 -99.795 ;
        RECT -64.765 -101.485 -64.435 -101.155 ;
        RECT -64.765 -102.845 -64.435 -102.515 ;
        RECT -64.765 -104.205 -64.435 -103.875 ;
        RECT -64.765 -105.565 -64.435 -105.235 ;
        RECT -64.765 -106.925 -64.435 -106.595 ;
        RECT -64.765 -108.285 -64.435 -107.955 ;
        RECT -64.765 -109.645 -64.435 -109.315 ;
        RECT -64.765 -111.005 -64.435 -110.675 ;
        RECT -64.76 -111.68 -64.44 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -63.405 244.04 -63.075 245.17 ;
        RECT -63.405 239.875 -63.075 240.205 ;
        RECT -63.405 238.515 -63.075 238.845 ;
        RECT -63.405 237.155 -63.075 237.485 ;
        RECT -63.405 235.795 -63.075 236.125 ;
        RECT -63.405 234.435 -63.075 234.765 ;
        RECT -63.405 233.075 -63.075 233.405 ;
        RECT -63.405 231.715 -63.075 232.045 ;
        RECT -63.405 230.355 -63.075 230.685 ;
        RECT -63.405 228.995 -63.075 229.325 ;
        RECT -63.405 227.635 -63.075 227.965 ;
        RECT -63.405 226.275 -63.075 226.605 ;
        RECT -63.405 224.915 -63.075 225.245 ;
        RECT -63.405 223.555 -63.075 223.885 ;
        RECT -63.405 222.195 -63.075 222.525 ;
        RECT -63.405 220.835 -63.075 221.165 ;
        RECT -63.405 219.475 -63.075 219.805 ;
        RECT -63.405 218.115 -63.075 218.445 ;
        RECT -63.405 216.755 -63.075 217.085 ;
        RECT -63.405 215.395 -63.075 215.725 ;
        RECT -63.405 214.035 -63.075 214.365 ;
        RECT -63.405 212.675 -63.075 213.005 ;
        RECT -63.405 211.315 -63.075 211.645 ;
        RECT -63.405 209.955 -63.075 210.285 ;
        RECT -63.405 208.595 -63.075 208.925 ;
        RECT -63.405 207.235 -63.075 207.565 ;
        RECT -63.405 205.875 -63.075 206.205 ;
        RECT -63.405 204.515 -63.075 204.845 ;
        RECT -63.405 203.155 -63.075 203.485 ;
        RECT -63.405 201.795 -63.075 202.125 ;
        RECT -63.405 200.435 -63.075 200.765 ;
        RECT -63.405 199.075 -63.075 199.405 ;
        RECT -63.405 197.715 -63.075 198.045 ;
        RECT -63.405 196.355 -63.075 196.685 ;
        RECT -63.405 194.995 -63.075 195.325 ;
        RECT -63.405 193.635 -63.075 193.965 ;
        RECT -63.405 192.275 -63.075 192.605 ;
        RECT -63.405 190.915 -63.075 191.245 ;
        RECT -63.405 189.555 -63.075 189.885 ;
        RECT -63.405 188.195 -63.075 188.525 ;
        RECT -63.405 186.835 -63.075 187.165 ;
        RECT -63.405 185.475 -63.075 185.805 ;
        RECT -63.405 184.115 -63.075 184.445 ;
        RECT -63.405 182.755 -63.075 183.085 ;
        RECT -63.405 181.395 -63.075 181.725 ;
        RECT -63.405 180.035 -63.075 180.365 ;
        RECT -63.405 178.675 -63.075 179.005 ;
        RECT -63.405 177.315 -63.075 177.645 ;
        RECT -63.405 175.955 -63.075 176.285 ;
        RECT -63.405 174.595 -63.075 174.925 ;
        RECT -63.405 173.235 -63.075 173.565 ;
        RECT -63.405 171.875 -63.075 172.205 ;
        RECT -63.405 170.515 -63.075 170.845 ;
        RECT -63.405 169.155 -63.075 169.485 ;
        RECT -63.405 167.795 -63.075 168.125 ;
        RECT -63.405 166.435 -63.075 166.765 ;
        RECT -63.405 165.075 -63.075 165.405 ;
        RECT -63.405 163.715 -63.075 164.045 ;
        RECT -63.405 162.355 -63.075 162.685 ;
        RECT -63.405 160.995 -63.075 161.325 ;
        RECT -63.405 159.635 -63.075 159.965 ;
        RECT -63.405 158.275 -63.075 158.605 ;
        RECT -63.405 156.915 -63.075 157.245 ;
        RECT -63.405 155.555 -63.075 155.885 ;
        RECT -63.405 154.195 -63.075 154.525 ;
        RECT -63.405 152.835 -63.075 153.165 ;
        RECT -63.405 151.475 -63.075 151.805 ;
        RECT -63.405 150.115 -63.075 150.445 ;
        RECT -63.405 148.755 -63.075 149.085 ;
        RECT -63.405 147.395 -63.075 147.725 ;
        RECT -63.405 146.035 -63.075 146.365 ;
        RECT -63.405 144.675 -63.075 145.005 ;
        RECT -63.405 143.315 -63.075 143.645 ;
        RECT -63.405 141.955 -63.075 142.285 ;
        RECT -63.405 140.595 -63.075 140.925 ;
        RECT -63.405 139.235 -63.075 139.565 ;
        RECT -63.405 136.42 -63.075 136.75 ;
        RECT -63.405 134.245 -63.075 134.575 ;
        RECT -63.405 133.395 -63.075 133.725 ;
        RECT -63.405 131.085 -63.075 131.415 ;
        RECT -63.405 130.235 -63.075 130.565 ;
        RECT -63.405 127.925 -63.075 128.255 ;
        RECT -63.405 127.075 -63.075 127.405 ;
        RECT -63.405 124.765 -63.075 125.095 ;
        RECT -63.405 123.915 -63.075 124.245 ;
        RECT -63.405 121.605 -63.075 121.935 ;
        RECT -63.405 120.755 -63.075 121.085 ;
        RECT -63.405 118.445 -63.075 118.775 ;
        RECT -63.405 117.595 -63.075 117.925 ;
        RECT -63.405 115.285 -63.075 115.615 ;
        RECT -63.405 114.435 -63.075 114.765 ;
        RECT -63.405 112.125 -63.075 112.455 ;
        RECT -63.405 111.275 -63.075 111.605 ;
        RECT -63.405 108.965 -63.075 109.295 ;
        RECT -63.405 108.115 -63.075 108.445 ;
        RECT -63.405 105.805 -63.075 106.135 ;
        RECT -63.405 104.955 -63.075 105.285 ;
        RECT -63.405 102.645 -63.075 102.975 ;
        RECT -63.405 101.795 -63.075 102.125 ;
        RECT -63.405 99.62 -63.075 99.95 ;
        RECT -63.405 97.075 -63.075 97.405 ;
        RECT -63.405 95.715 -63.075 96.045 ;
        RECT -63.405 94.355 -63.075 94.685 ;
        RECT -63.405 92.995 -63.075 93.325 ;
        RECT -63.405 91.635 -63.075 91.965 ;
        RECT -63.405 90.275 -63.075 90.605 ;
        RECT -63.405 88.915 -63.075 89.245 ;
        RECT -63.405 87.555 -63.075 87.885 ;
        RECT -63.405 86.195 -63.075 86.525 ;
        RECT -63.405 84.835 -63.075 85.165 ;
        RECT -63.405 83.475 -63.075 83.805 ;
        RECT -63.405 82.115 -63.075 82.445 ;
        RECT -63.405 80.755 -63.075 81.085 ;
        RECT -63.405 79.395 -63.075 79.725 ;
        RECT -63.405 78.035 -63.075 78.365 ;
        RECT -63.405 76.675 -63.075 77.005 ;
        RECT -63.405 75.315 -63.075 75.645 ;
        RECT -63.405 73.955 -63.075 74.285 ;
        RECT -63.405 72.595 -63.075 72.925 ;
        RECT -63.405 71.235 -63.075 71.565 ;
        RECT -63.405 69.875 -63.075 70.205 ;
        RECT -63.405 68.515 -63.075 68.845 ;
        RECT -63.405 67.155 -63.075 67.485 ;
        RECT -63.405 65.795 -63.075 66.125 ;
        RECT -63.405 64.435 -63.075 64.765 ;
        RECT -63.405 63.075 -63.075 63.405 ;
        RECT -63.405 61.715 -63.075 62.045 ;
        RECT -63.405 60.355 -63.075 60.685 ;
        RECT -63.405 58.995 -63.075 59.325 ;
        RECT -63.405 57.635 -63.075 57.965 ;
        RECT -63.405 56.275 -63.075 56.605 ;
        RECT -63.405 54.915 -63.075 55.245 ;
        RECT -63.405 53.555 -63.075 53.885 ;
        RECT -63.405 52.195 -63.075 52.525 ;
        RECT -63.405 50.835 -63.075 51.165 ;
        RECT -63.405 49.475 -63.075 49.805 ;
        RECT -63.405 48.115 -63.075 48.445 ;
        RECT -63.405 46.755 -63.075 47.085 ;
        RECT -63.405 45.395 -63.075 45.725 ;
        RECT -63.405 44.035 -63.075 44.365 ;
        RECT -63.405 42.675 -63.075 43.005 ;
        RECT -63.405 41.315 -63.075 41.645 ;
        RECT -63.405 39.955 -63.075 40.285 ;
        RECT -63.405 38.595 -63.075 38.925 ;
        RECT -63.405 37.235 -63.075 37.565 ;
        RECT -63.405 35.875 -63.075 36.205 ;
        RECT -63.405 34.515 -63.075 34.845 ;
        RECT -63.405 33.155 -63.075 33.485 ;
        RECT -63.405 31.795 -63.075 32.125 ;
        RECT -63.405 30.435 -63.075 30.765 ;
        RECT -63.405 29.075 -63.075 29.405 ;
        RECT -63.405 27.715 -63.075 28.045 ;
        RECT -63.405 26.355 -63.075 26.685 ;
        RECT -63.405 24.995 -63.075 25.325 ;
        RECT -63.405 23.635 -63.075 23.965 ;
        RECT -63.405 22.275 -63.075 22.605 ;
        RECT -63.405 20.915 -63.075 21.245 ;
        RECT -63.405 19.555 -63.075 19.885 ;
        RECT -63.405 18.195 -63.075 18.525 ;
        RECT -63.405 16.835 -63.075 17.165 ;
        RECT -63.405 15.475 -63.075 15.805 ;
        RECT -63.405 14.115 -63.075 14.445 ;
        RECT -63.405 12.755 -63.075 13.085 ;
        RECT -63.405 11.395 -63.075 11.725 ;
        RECT -63.405 10.035 -63.075 10.365 ;
        RECT -63.405 8.675 -63.075 9.005 ;
        RECT -63.405 7.315 -63.075 7.645 ;
        RECT -63.405 5.955 -63.075 6.285 ;
        RECT -63.405 4.595 -63.075 4.925 ;
        RECT -63.405 3.235 -63.075 3.565 ;
        RECT -63.405 1.875 -63.075 2.205 ;
        RECT -63.405 0.515 -63.075 0.845 ;
        RECT -63.405 -0.845 -63.075 -0.515 ;
        RECT -63.405 -2.205 -63.075 -1.875 ;
        RECT -63.405 -3.565 -63.075 -3.235 ;
        RECT -63.405 -4.925 -63.075 -4.595 ;
        RECT -63.405 -6.285 -63.075 -5.955 ;
        RECT -63.405 -7.645 -63.075 -7.315 ;
        RECT -63.405 -9.005 -63.075 -8.675 ;
        RECT -63.405 -10.365 -63.075 -10.035 ;
        RECT -63.405 -11.725 -63.075 -11.395 ;
        RECT -63.405 -13.085 -63.075 -12.755 ;
        RECT -63.405 -14.445 -63.075 -14.115 ;
        RECT -63.405 -15.805 -63.075 -15.475 ;
        RECT -63.405 -17.165 -63.075 -16.835 ;
        RECT -63.405 -18.525 -63.075 -18.195 ;
        RECT -63.405 -19.885 -63.075 -19.555 ;
        RECT -63.405 -21.245 -63.075 -20.915 ;
        RECT -63.405 -22.605 -63.075 -22.275 ;
        RECT -63.405 -23.965 -63.075 -23.635 ;
        RECT -63.405 -25.325 -63.075 -24.995 ;
        RECT -63.405 -26.685 -63.075 -26.355 ;
        RECT -63.405 -28.045 -63.075 -27.715 ;
        RECT -63.405 -29.405 -63.075 -29.075 ;
        RECT -63.405 -30.765 -63.075 -30.435 ;
        RECT -63.405 -32.125 -63.075 -31.795 ;
        RECT -63.405 -33.485 -63.075 -33.155 ;
        RECT -63.405 -34.845 -63.075 -34.515 ;
        RECT -63.405 -36.205 -63.075 -35.875 ;
        RECT -63.405 -37.565 -63.075 -37.235 ;
        RECT -63.405 -38.925 -63.075 -38.595 ;
        RECT -63.405 -40.285 -63.075 -39.955 ;
        RECT -63.405 -41.645 -63.075 -41.315 ;
        RECT -63.405 -43.005 -63.075 -42.675 ;
        RECT -63.405 -44.365 -63.075 -44.035 ;
        RECT -63.405 -45.725 -63.075 -45.395 ;
        RECT -63.405 -47.085 -63.075 -46.755 ;
        RECT -63.405 -48.445 -63.075 -48.115 ;
        RECT -63.405 -49.805 -63.075 -49.475 ;
        RECT -63.405 -51.165 -63.075 -50.835 ;
        RECT -63.405 -52.525 -63.075 -52.195 ;
        RECT -63.405 -53.885 -63.075 -53.555 ;
        RECT -63.405 -55.245 -63.075 -54.915 ;
        RECT -63.405 -56.605 -63.075 -56.275 ;
        RECT -63.405 -57.965 -63.075 -57.635 ;
        RECT -63.405 -59.325 -63.075 -58.995 ;
        RECT -63.405 -60.685 -63.075 -60.355 ;
        RECT -63.405 -62.045 -63.075 -61.715 ;
        RECT -63.405 -63.405 -63.075 -63.075 ;
        RECT -63.405 -64.765 -63.075 -64.435 ;
        RECT -63.405 -66.125 -63.075 -65.795 ;
        RECT -63.405 -67.485 -63.075 -67.155 ;
        RECT -63.405 -68.845 -63.075 -68.515 ;
        RECT -63.405 -70.205 -63.075 -69.875 ;
        RECT -63.405 -71.565 -63.075 -71.235 ;
        RECT -63.405 -72.925 -63.075 -72.595 ;
        RECT -63.405 -74.285 -63.075 -73.955 ;
        RECT -63.405 -75.645 -63.075 -75.315 ;
        RECT -63.405 -77.005 -63.075 -76.675 ;
        RECT -63.405 -78.365 -63.075 -78.035 ;
        RECT -63.405 -79.725 -63.075 -79.395 ;
        RECT -63.405 -81.085 -63.075 -80.755 ;
        RECT -63.405 -82.445 -63.075 -82.115 ;
        RECT -63.405 -83.805 -63.075 -83.475 ;
        RECT -63.405 -85.165 -63.075 -84.835 ;
        RECT -63.405 -86.525 -63.075 -86.195 ;
        RECT -63.405 -87.885 -63.075 -87.555 ;
        RECT -63.405 -89.245 -63.075 -88.915 ;
        RECT -63.405 -90.605 -63.075 -90.275 ;
        RECT -63.405 -91.965 -63.075 -91.635 ;
        RECT -63.405 -93.325 -63.075 -92.995 ;
        RECT -63.405 -94.685 -63.075 -94.355 ;
        RECT -63.405 -96.045 -63.075 -95.715 ;
        RECT -63.405 -97.405 -63.075 -97.075 ;
        RECT -63.405 -98.765 -63.075 -98.435 ;
        RECT -63.405 -100.125 -63.075 -99.795 ;
        RECT -63.405 -101.485 -63.075 -101.155 ;
        RECT -63.405 -102.845 -63.075 -102.515 ;
        RECT -63.405 -104.205 -63.075 -103.875 ;
        RECT -63.405 -105.565 -63.075 -105.235 ;
        RECT -63.405 -106.925 -63.075 -106.595 ;
        RECT -63.405 -108.285 -63.075 -107.955 ;
        RECT -63.405 -109.645 -63.075 -109.315 ;
        RECT -63.405 -111.005 -63.075 -110.675 ;
        RECT -63.405 -113.725 -63.075 -113.395 ;
        RECT -63.405 -115.085 -63.075 -114.755 ;
        RECT -63.405 -116.445 -63.075 -116.115 ;
        RECT -63.405 -117.805 -63.075 -117.475 ;
        RECT -63.405 -119.165 -63.075 -118.835 ;
        RECT -63.405 -120.525 -63.075 -120.195 ;
        RECT -63.405 -121.885 -63.075 -121.555 ;
        RECT -63.405 -123.245 -63.075 -122.915 ;
        RECT -63.405 -124.605 -63.075 -124.275 ;
        RECT -63.405 -125.965 -63.075 -125.635 ;
        RECT -63.405 -127.325 -63.075 -126.995 ;
        RECT -63.405 -128.685 -63.075 -128.355 ;
        RECT -63.405 -130.045 -63.075 -129.715 ;
        RECT -63.405 -131.405 -63.075 -131.075 ;
        RECT -63.405 -132.765 -63.075 -132.435 ;
        RECT -63.405 -134.125 -63.075 -133.795 ;
        RECT -63.405 -135.485 -63.075 -135.155 ;
        RECT -63.405 -136.845 -63.075 -136.515 ;
        RECT -63.405 -138.205 -63.075 -137.875 ;
        RECT -63.405 -139.565 -63.075 -139.235 ;
        RECT -63.405 -140.925 -63.075 -140.595 ;
        RECT -63.405 -142.285 -63.075 -141.955 ;
        RECT -63.405 -143.645 -63.075 -143.315 ;
        RECT -63.405 -145.005 -63.075 -144.675 ;
        RECT -63.405 -146.365 -63.075 -146.035 ;
        RECT -63.405 -147.725 -63.075 -147.395 ;
        RECT -63.405 -149.085 -63.075 -148.755 ;
        RECT -63.405 -150.445 -63.075 -150.115 ;
        RECT -63.405 -151.805 -63.075 -151.475 ;
        RECT -63.405 -153.165 -63.075 -152.835 ;
        RECT -63.405 -154.525 -63.075 -154.195 ;
        RECT -63.405 -155.885 -63.075 -155.555 ;
        RECT -63.405 -157.245 -63.075 -156.915 ;
        RECT -63.405 -158.605 -63.075 -158.275 ;
        RECT -63.405 -159.965 -63.075 -159.635 ;
        RECT -63.405 -161.325 -63.075 -160.995 ;
        RECT -63.405 -162.685 -63.075 -162.355 ;
        RECT -63.405 -164.045 -63.075 -163.715 ;
        RECT -63.405 -165.405 -63.075 -165.075 ;
        RECT -63.405 -166.765 -63.075 -166.435 ;
        RECT -63.405 -168.655 -63.075 -168.325 ;
        RECT -63.405 -169.485 -63.075 -169.155 ;
        RECT -63.405 -170.845 -63.075 -170.515 ;
        RECT -63.405 -174.925 -63.075 -174.595 ;
        RECT -63.405 -177.645 -63.075 -177.315 ;
        RECT -63.405 -183.29 -63.075 -182.16 ;
        RECT -63.4 -183.405 -63.08 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -62.045 -55.245 -61.715 -54.915 ;
        RECT -62.045 -56.605 -61.715 -56.275 ;
        RECT -62.045 -57.965 -61.715 -57.635 ;
        RECT -62.045 -59.325 -61.715 -58.995 ;
        RECT -62.045 -60.685 -61.715 -60.355 ;
        RECT -62.045 -62.045 -61.715 -61.715 ;
        RECT -62.045 -63.405 -61.715 -63.075 ;
        RECT -62.045 -64.765 -61.715 -64.435 ;
        RECT -62.045 -66.125 -61.715 -65.795 ;
        RECT -62.045 -67.485 -61.715 -67.155 ;
        RECT -62.045 -68.845 -61.715 -68.515 ;
        RECT -62.045 -70.205 -61.715 -69.875 ;
        RECT -62.045 -71.565 -61.715 -71.235 ;
        RECT -62.045 -72.925 -61.715 -72.595 ;
        RECT -62.045 -74.285 -61.715 -73.955 ;
        RECT -62.045 -75.645 -61.715 -75.315 ;
        RECT -62.045 -77.005 -61.715 -76.675 ;
        RECT -62.045 -78.365 -61.715 -78.035 ;
        RECT -62.045 -79.725 -61.715 -79.395 ;
        RECT -62.045 -81.085 -61.715 -80.755 ;
        RECT -62.045 -82.445 -61.715 -82.115 ;
        RECT -62.045 -83.805 -61.715 -83.475 ;
        RECT -62.045 -85.165 -61.715 -84.835 ;
        RECT -62.045 -86.525 -61.715 -86.195 ;
        RECT -62.045 -87.885 -61.715 -87.555 ;
        RECT -62.045 -89.245 -61.715 -88.915 ;
        RECT -62.045 -90.605 -61.715 -90.275 ;
        RECT -62.045 -91.965 -61.715 -91.635 ;
        RECT -62.045 -93.325 -61.715 -92.995 ;
        RECT -62.045 -94.685 -61.715 -94.355 ;
        RECT -62.045 -96.045 -61.715 -95.715 ;
        RECT -62.045 -97.405 -61.715 -97.075 ;
        RECT -62.045 -98.765 -61.715 -98.435 ;
        RECT -62.045 -100.125 -61.715 -99.795 ;
        RECT -62.045 -101.485 -61.715 -101.155 ;
        RECT -62.045 -102.845 -61.715 -102.515 ;
        RECT -62.045 -104.205 -61.715 -103.875 ;
        RECT -62.045 -105.565 -61.715 -105.235 ;
        RECT -62.045 -106.925 -61.715 -106.595 ;
        RECT -62.045 -108.285 -61.715 -107.955 ;
        RECT -62.045 -109.645 -61.715 -109.315 ;
        RECT -62.04 -111 -61.72 245.285 ;
        RECT -62.045 244.04 -61.715 245.17 ;
        RECT -62.045 239.875 -61.715 240.205 ;
        RECT -62.045 238.515 -61.715 238.845 ;
        RECT -62.045 237.155 -61.715 237.485 ;
        RECT -62.045 235.795 -61.715 236.125 ;
        RECT -62.045 234.435 -61.715 234.765 ;
        RECT -62.045 233.075 -61.715 233.405 ;
        RECT -62.045 231.715 -61.715 232.045 ;
        RECT -62.045 230.355 -61.715 230.685 ;
        RECT -62.045 228.995 -61.715 229.325 ;
        RECT -62.045 227.635 -61.715 227.965 ;
        RECT -62.045 226.275 -61.715 226.605 ;
        RECT -62.045 224.915 -61.715 225.245 ;
        RECT -62.045 223.555 -61.715 223.885 ;
        RECT -62.045 222.195 -61.715 222.525 ;
        RECT -62.045 220.835 -61.715 221.165 ;
        RECT -62.045 219.475 -61.715 219.805 ;
        RECT -62.045 218.115 -61.715 218.445 ;
        RECT -62.045 216.755 -61.715 217.085 ;
        RECT -62.045 215.395 -61.715 215.725 ;
        RECT -62.045 214.035 -61.715 214.365 ;
        RECT -62.045 212.675 -61.715 213.005 ;
        RECT -62.045 211.315 -61.715 211.645 ;
        RECT -62.045 209.955 -61.715 210.285 ;
        RECT -62.045 208.595 -61.715 208.925 ;
        RECT -62.045 207.235 -61.715 207.565 ;
        RECT -62.045 205.875 -61.715 206.205 ;
        RECT -62.045 204.515 -61.715 204.845 ;
        RECT -62.045 203.155 -61.715 203.485 ;
        RECT -62.045 201.795 -61.715 202.125 ;
        RECT -62.045 200.435 -61.715 200.765 ;
        RECT -62.045 199.075 -61.715 199.405 ;
        RECT -62.045 197.715 -61.715 198.045 ;
        RECT -62.045 196.355 -61.715 196.685 ;
        RECT -62.045 194.995 -61.715 195.325 ;
        RECT -62.045 193.635 -61.715 193.965 ;
        RECT -62.045 192.275 -61.715 192.605 ;
        RECT -62.045 190.915 -61.715 191.245 ;
        RECT -62.045 189.555 -61.715 189.885 ;
        RECT -62.045 188.195 -61.715 188.525 ;
        RECT -62.045 186.835 -61.715 187.165 ;
        RECT -62.045 185.475 -61.715 185.805 ;
        RECT -62.045 184.115 -61.715 184.445 ;
        RECT -62.045 182.755 -61.715 183.085 ;
        RECT -62.045 181.395 -61.715 181.725 ;
        RECT -62.045 180.035 -61.715 180.365 ;
        RECT -62.045 178.675 -61.715 179.005 ;
        RECT -62.045 177.315 -61.715 177.645 ;
        RECT -62.045 175.955 -61.715 176.285 ;
        RECT -62.045 174.595 -61.715 174.925 ;
        RECT -62.045 173.235 -61.715 173.565 ;
        RECT -62.045 171.875 -61.715 172.205 ;
        RECT -62.045 170.515 -61.715 170.845 ;
        RECT -62.045 169.155 -61.715 169.485 ;
        RECT -62.045 167.795 -61.715 168.125 ;
        RECT -62.045 166.435 -61.715 166.765 ;
        RECT -62.045 165.075 -61.715 165.405 ;
        RECT -62.045 163.715 -61.715 164.045 ;
        RECT -62.045 162.355 -61.715 162.685 ;
        RECT -62.045 160.995 -61.715 161.325 ;
        RECT -62.045 159.635 -61.715 159.965 ;
        RECT -62.045 158.275 -61.715 158.605 ;
        RECT -62.045 156.915 -61.715 157.245 ;
        RECT -62.045 155.555 -61.715 155.885 ;
        RECT -62.045 154.195 -61.715 154.525 ;
        RECT -62.045 152.835 -61.715 153.165 ;
        RECT -62.045 151.475 -61.715 151.805 ;
        RECT -62.045 150.115 -61.715 150.445 ;
        RECT -62.045 148.755 -61.715 149.085 ;
        RECT -62.045 147.395 -61.715 147.725 ;
        RECT -62.045 146.035 -61.715 146.365 ;
        RECT -62.045 144.675 -61.715 145.005 ;
        RECT -62.045 143.315 -61.715 143.645 ;
        RECT -62.045 141.955 -61.715 142.285 ;
        RECT -62.045 140.595 -61.715 140.925 ;
        RECT -62.045 139.235 -61.715 139.565 ;
        RECT -62.045 136.42 -61.715 136.75 ;
        RECT -62.045 134.245 -61.715 134.575 ;
        RECT -62.045 133.395 -61.715 133.725 ;
        RECT -62.045 131.085 -61.715 131.415 ;
        RECT -62.045 130.235 -61.715 130.565 ;
        RECT -62.045 127.925 -61.715 128.255 ;
        RECT -62.045 127.075 -61.715 127.405 ;
        RECT -62.045 124.765 -61.715 125.095 ;
        RECT -62.045 123.915 -61.715 124.245 ;
        RECT -62.045 121.605 -61.715 121.935 ;
        RECT -62.045 120.755 -61.715 121.085 ;
        RECT -62.045 118.445 -61.715 118.775 ;
        RECT -62.045 117.595 -61.715 117.925 ;
        RECT -62.045 115.285 -61.715 115.615 ;
        RECT -62.045 114.435 -61.715 114.765 ;
        RECT -62.045 112.125 -61.715 112.455 ;
        RECT -62.045 111.275 -61.715 111.605 ;
        RECT -62.045 108.965 -61.715 109.295 ;
        RECT -62.045 108.115 -61.715 108.445 ;
        RECT -62.045 105.805 -61.715 106.135 ;
        RECT -62.045 104.955 -61.715 105.285 ;
        RECT -62.045 102.645 -61.715 102.975 ;
        RECT -62.045 101.795 -61.715 102.125 ;
        RECT -62.045 99.62 -61.715 99.95 ;
        RECT -62.045 97.075 -61.715 97.405 ;
        RECT -62.045 95.715 -61.715 96.045 ;
        RECT -62.045 94.355 -61.715 94.685 ;
        RECT -62.045 92.995 -61.715 93.325 ;
        RECT -62.045 91.635 -61.715 91.965 ;
        RECT -62.045 90.275 -61.715 90.605 ;
        RECT -62.045 88.915 -61.715 89.245 ;
        RECT -62.045 87.555 -61.715 87.885 ;
        RECT -62.045 86.195 -61.715 86.525 ;
        RECT -62.045 84.835 -61.715 85.165 ;
        RECT -62.045 83.475 -61.715 83.805 ;
        RECT -62.045 82.115 -61.715 82.445 ;
        RECT -62.045 80.755 -61.715 81.085 ;
        RECT -62.045 79.395 -61.715 79.725 ;
        RECT -62.045 78.035 -61.715 78.365 ;
        RECT -62.045 76.675 -61.715 77.005 ;
        RECT -62.045 75.315 -61.715 75.645 ;
        RECT -62.045 73.955 -61.715 74.285 ;
        RECT -62.045 72.595 -61.715 72.925 ;
        RECT -62.045 71.235 -61.715 71.565 ;
        RECT -62.045 69.875 -61.715 70.205 ;
        RECT -62.045 68.515 -61.715 68.845 ;
        RECT -62.045 67.155 -61.715 67.485 ;
        RECT -62.045 65.795 -61.715 66.125 ;
        RECT -62.045 64.435 -61.715 64.765 ;
        RECT -62.045 63.075 -61.715 63.405 ;
        RECT -62.045 61.715 -61.715 62.045 ;
        RECT -62.045 60.355 -61.715 60.685 ;
        RECT -62.045 58.995 -61.715 59.325 ;
        RECT -62.045 57.635 -61.715 57.965 ;
        RECT -62.045 56.275 -61.715 56.605 ;
        RECT -62.045 54.915 -61.715 55.245 ;
        RECT -62.045 53.555 -61.715 53.885 ;
        RECT -62.045 52.195 -61.715 52.525 ;
        RECT -62.045 50.835 -61.715 51.165 ;
        RECT -62.045 49.475 -61.715 49.805 ;
        RECT -62.045 48.115 -61.715 48.445 ;
        RECT -62.045 46.755 -61.715 47.085 ;
        RECT -62.045 45.395 -61.715 45.725 ;
        RECT -62.045 44.035 -61.715 44.365 ;
        RECT -62.045 42.675 -61.715 43.005 ;
        RECT -62.045 41.315 -61.715 41.645 ;
        RECT -62.045 39.955 -61.715 40.285 ;
        RECT -62.045 38.595 -61.715 38.925 ;
        RECT -62.045 37.235 -61.715 37.565 ;
        RECT -62.045 35.875 -61.715 36.205 ;
        RECT -62.045 34.515 -61.715 34.845 ;
        RECT -62.045 33.155 -61.715 33.485 ;
        RECT -62.045 31.795 -61.715 32.125 ;
        RECT -62.045 30.435 -61.715 30.765 ;
        RECT -62.045 29.075 -61.715 29.405 ;
        RECT -62.045 27.715 -61.715 28.045 ;
        RECT -62.045 26.355 -61.715 26.685 ;
        RECT -62.045 24.995 -61.715 25.325 ;
        RECT -62.045 23.635 -61.715 23.965 ;
        RECT -62.045 22.275 -61.715 22.605 ;
        RECT -62.045 20.915 -61.715 21.245 ;
        RECT -62.045 19.555 -61.715 19.885 ;
        RECT -62.045 18.195 -61.715 18.525 ;
        RECT -62.045 16.835 -61.715 17.165 ;
        RECT -62.045 15.475 -61.715 15.805 ;
        RECT -62.045 14.115 -61.715 14.445 ;
        RECT -62.045 12.755 -61.715 13.085 ;
        RECT -62.045 11.395 -61.715 11.725 ;
        RECT -62.045 10.035 -61.715 10.365 ;
        RECT -62.045 8.675 -61.715 9.005 ;
        RECT -62.045 7.315 -61.715 7.645 ;
        RECT -62.045 5.955 -61.715 6.285 ;
        RECT -62.045 4.595 -61.715 4.925 ;
        RECT -62.045 3.235 -61.715 3.565 ;
        RECT -62.045 1.875 -61.715 2.205 ;
        RECT -62.045 0.515 -61.715 0.845 ;
        RECT -62.045 -0.845 -61.715 -0.515 ;
        RECT -62.045 -2.205 -61.715 -1.875 ;
        RECT -62.045 -3.565 -61.715 -3.235 ;
        RECT -62.045 -4.925 -61.715 -4.595 ;
        RECT -62.045 -6.285 -61.715 -5.955 ;
        RECT -62.045 -7.645 -61.715 -7.315 ;
        RECT -62.045 -9.005 -61.715 -8.675 ;
        RECT -62.045 -10.365 -61.715 -10.035 ;
        RECT -62.045 -11.725 -61.715 -11.395 ;
        RECT -62.045 -13.085 -61.715 -12.755 ;
        RECT -62.045 -14.445 -61.715 -14.115 ;
        RECT -62.045 -15.805 -61.715 -15.475 ;
        RECT -62.045 -17.165 -61.715 -16.835 ;
        RECT -62.045 -18.525 -61.715 -18.195 ;
        RECT -62.045 -19.885 -61.715 -19.555 ;
        RECT -62.045 -21.245 -61.715 -20.915 ;
        RECT -62.045 -22.605 -61.715 -22.275 ;
        RECT -62.045 -23.965 -61.715 -23.635 ;
        RECT -62.045 -25.325 -61.715 -24.995 ;
        RECT -62.045 -26.685 -61.715 -26.355 ;
        RECT -62.045 -28.045 -61.715 -27.715 ;
        RECT -62.045 -29.405 -61.715 -29.075 ;
        RECT -62.045 -30.765 -61.715 -30.435 ;
        RECT -62.045 -32.125 -61.715 -31.795 ;
        RECT -62.045 -33.485 -61.715 -33.155 ;
        RECT -62.045 -34.845 -61.715 -34.515 ;
        RECT -62.045 -36.205 -61.715 -35.875 ;
        RECT -62.045 -37.565 -61.715 -37.235 ;
        RECT -62.045 -38.925 -61.715 -38.595 ;
        RECT -62.045 -40.285 -61.715 -39.955 ;
        RECT -62.045 -41.645 -61.715 -41.315 ;
        RECT -62.045 -43.005 -61.715 -42.675 ;
        RECT -62.045 -44.365 -61.715 -44.035 ;
        RECT -62.045 -45.725 -61.715 -45.395 ;
        RECT -62.045 -47.085 -61.715 -46.755 ;
        RECT -62.045 -48.445 -61.715 -48.115 ;
        RECT -62.045 -49.805 -61.715 -49.475 ;
        RECT -62.045 -51.165 -61.715 -50.835 ;
        RECT -62.045 -52.525 -61.715 -52.195 ;
        RECT -62.045 -53.885 -61.715 -53.555 ;
    END
    PORT
      LAYER met3 ;
        RECT -70.205 244.04 -69.875 245.17 ;
        RECT -70.205 239.875 -69.875 240.205 ;
        RECT -70.205 238.515 -69.875 238.845 ;
        RECT -70.205 237.155 -69.875 237.485 ;
        RECT -70.205 235.795 -69.875 236.125 ;
        RECT -70.205 234.435 -69.875 234.765 ;
        RECT -70.205 233.075 -69.875 233.405 ;
        RECT -70.205 231.715 -69.875 232.045 ;
        RECT -70.205 230.355 -69.875 230.685 ;
        RECT -70.205 228.995 -69.875 229.325 ;
        RECT -70.205 227.635 -69.875 227.965 ;
        RECT -70.205 226.275 -69.875 226.605 ;
        RECT -70.205 224.915 -69.875 225.245 ;
        RECT -70.205 223.555 -69.875 223.885 ;
        RECT -70.205 222.195 -69.875 222.525 ;
        RECT -70.205 220.835 -69.875 221.165 ;
        RECT -70.205 219.475 -69.875 219.805 ;
        RECT -70.205 218.115 -69.875 218.445 ;
        RECT -70.205 216.755 -69.875 217.085 ;
        RECT -70.205 215.395 -69.875 215.725 ;
        RECT -70.205 214.035 -69.875 214.365 ;
        RECT -70.205 212.675 -69.875 213.005 ;
        RECT -70.205 211.315 -69.875 211.645 ;
        RECT -70.205 209.955 -69.875 210.285 ;
        RECT -70.205 208.595 -69.875 208.925 ;
        RECT -70.205 207.235 -69.875 207.565 ;
        RECT -70.205 205.875 -69.875 206.205 ;
        RECT -70.205 204.515 -69.875 204.845 ;
        RECT -70.205 203.155 -69.875 203.485 ;
        RECT -70.205 201.795 -69.875 202.125 ;
        RECT -70.205 200.435 -69.875 200.765 ;
        RECT -70.205 199.075 -69.875 199.405 ;
        RECT -70.205 197.715 -69.875 198.045 ;
        RECT -70.205 196.355 -69.875 196.685 ;
        RECT -70.205 194.995 -69.875 195.325 ;
        RECT -70.205 193.635 -69.875 193.965 ;
        RECT -70.205 192.275 -69.875 192.605 ;
        RECT -70.205 190.915 -69.875 191.245 ;
        RECT -70.205 189.555 -69.875 189.885 ;
        RECT -70.205 188.195 -69.875 188.525 ;
        RECT -70.205 186.835 -69.875 187.165 ;
        RECT -70.205 185.475 -69.875 185.805 ;
        RECT -70.205 184.115 -69.875 184.445 ;
        RECT -70.205 182.755 -69.875 183.085 ;
        RECT -70.205 181.395 -69.875 181.725 ;
        RECT -70.205 180.035 -69.875 180.365 ;
        RECT -70.205 178.675 -69.875 179.005 ;
        RECT -70.205 177.315 -69.875 177.645 ;
        RECT -70.205 175.955 -69.875 176.285 ;
        RECT -70.205 174.595 -69.875 174.925 ;
        RECT -70.205 173.235 -69.875 173.565 ;
        RECT -70.205 171.875 -69.875 172.205 ;
        RECT -70.205 170.515 -69.875 170.845 ;
        RECT -70.205 169.155 -69.875 169.485 ;
        RECT -70.205 167.795 -69.875 168.125 ;
        RECT -70.205 166.435 -69.875 166.765 ;
        RECT -70.205 165.075 -69.875 165.405 ;
        RECT -70.205 163.715 -69.875 164.045 ;
        RECT -70.205 162.355 -69.875 162.685 ;
        RECT -70.205 160.995 -69.875 161.325 ;
        RECT -70.205 159.635 -69.875 159.965 ;
        RECT -70.205 158.275 -69.875 158.605 ;
        RECT -70.205 156.915 -69.875 157.245 ;
        RECT -70.205 155.555 -69.875 155.885 ;
        RECT -70.205 154.195 -69.875 154.525 ;
        RECT -70.205 152.835 -69.875 153.165 ;
        RECT -70.205 151.475 -69.875 151.805 ;
        RECT -70.205 150.115 -69.875 150.445 ;
        RECT -70.205 148.755 -69.875 149.085 ;
        RECT -70.205 147.395 -69.875 147.725 ;
        RECT -70.205 146.035 -69.875 146.365 ;
        RECT -70.205 144.675 -69.875 145.005 ;
        RECT -70.205 143.315 -69.875 143.645 ;
        RECT -70.205 141.955 -69.875 142.285 ;
        RECT -70.205 140.595 -69.875 140.925 ;
        RECT -70.205 139.235 -69.875 139.565 ;
        RECT -70.205 137.875 -69.875 138.205 ;
        RECT -70.205 136.515 -69.875 136.845 ;
        RECT -70.205 135.155 -69.875 135.485 ;
        RECT -70.205 133.795 -69.875 134.125 ;
        RECT -70.205 132.435 -69.875 132.765 ;
        RECT -70.205 131.075 -69.875 131.405 ;
        RECT -70.205 129.715 -69.875 130.045 ;
        RECT -70.205 128.355 -69.875 128.685 ;
        RECT -70.205 126.995 -69.875 127.325 ;
        RECT -70.205 125.635 -69.875 125.965 ;
        RECT -70.205 124.275 -69.875 124.605 ;
        RECT -70.205 122.915 -69.875 123.245 ;
        RECT -70.205 121.555 -69.875 121.885 ;
        RECT -70.205 120.195 -69.875 120.525 ;
        RECT -70.205 118.835 -69.875 119.165 ;
        RECT -70.205 117.475 -69.875 117.805 ;
        RECT -70.205 116.115 -69.875 116.445 ;
        RECT -70.205 114.755 -69.875 115.085 ;
        RECT -70.205 113.395 -69.875 113.725 ;
        RECT -70.205 112.035 -69.875 112.365 ;
        RECT -70.205 110.675 -69.875 111.005 ;
        RECT -70.205 109.315 -69.875 109.645 ;
        RECT -70.205 107.955 -69.875 108.285 ;
        RECT -70.205 106.595 -69.875 106.925 ;
        RECT -70.205 105.235 -69.875 105.565 ;
        RECT -70.205 103.875 -69.875 104.205 ;
        RECT -70.205 102.515 -69.875 102.845 ;
        RECT -70.205 101.155 -69.875 101.485 ;
        RECT -70.205 99.795 -69.875 100.125 ;
        RECT -70.205 98.435 -69.875 98.765 ;
        RECT -70.205 97.075 -69.875 97.405 ;
        RECT -70.205 95.715 -69.875 96.045 ;
        RECT -70.205 94.355 -69.875 94.685 ;
        RECT -70.205 92.995 -69.875 93.325 ;
        RECT -70.205 91.635 -69.875 91.965 ;
        RECT -70.205 90.275 -69.875 90.605 ;
        RECT -70.205 88.915 -69.875 89.245 ;
        RECT -70.205 87.555 -69.875 87.885 ;
        RECT -70.205 86.195 -69.875 86.525 ;
        RECT -70.205 84.835 -69.875 85.165 ;
        RECT -70.205 83.475 -69.875 83.805 ;
        RECT -70.205 82.115 -69.875 82.445 ;
        RECT -70.205 80.755 -69.875 81.085 ;
        RECT -70.205 79.395 -69.875 79.725 ;
        RECT -70.205 78.035 -69.875 78.365 ;
        RECT -70.205 76.675 -69.875 77.005 ;
        RECT -70.205 75.315 -69.875 75.645 ;
        RECT -70.205 73.955 -69.875 74.285 ;
        RECT -70.205 72.595 -69.875 72.925 ;
        RECT -70.205 71.235 -69.875 71.565 ;
        RECT -70.205 69.875 -69.875 70.205 ;
        RECT -70.205 68.515 -69.875 68.845 ;
        RECT -70.205 67.155 -69.875 67.485 ;
        RECT -70.205 65.795 -69.875 66.125 ;
        RECT -70.205 64.435 -69.875 64.765 ;
        RECT -70.205 63.075 -69.875 63.405 ;
        RECT -70.205 61.715 -69.875 62.045 ;
        RECT -70.205 60.355 -69.875 60.685 ;
        RECT -70.205 58.995 -69.875 59.325 ;
        RECT -70.205 57.635 -69.875 57.965 ;
        RECT -70.205 56.275 -69.875 56.605 ;
        RECT -70.205 54.915 -69.875 55.245 ;
        RECT -70.205 53.555 -69.875 53.885 ;
        RECT -70.205 52.195 -69.875 52.525 ;
        RECT -70.205 50.835 -69.875 51.165 ;
        RECT -70.205 49.475 -69.875 49.805 ;
        RECT -70.205 48.115 -69.875 48.445 ;
        RECT -70.205 46.755 -69.875 47.085 ;
        RECT -70.205 45.395 -69.875 45.725 ;
        RECT -70.205 44.035 -69.875 44.365 ;
        RECT -70.205 42.675 -69.875 43.005 ;
        RECT -70.205 41.315 -69.875 41.645 ;
        RECT -70.205 39.955 -69.875 40.285 ;
        RECT -70.205 38.595 -69.875 38.925 ;
        RECT -70.205 37.235 -69.875 37.565 ;
        RECT -70.205 35.875 -69.875 36.205 ;
        RECT -70.205 34.515 -69.875 34.845 ;
        RECT -70.205 33.155 -69.875 33.485 ;
        RECT -70.205 31.795 -69.875 32.125 ;
        RECT -70.205 30.435 -69.875 30.765 ;
        RECT -70.205 29.075 -69.875 29.405 ;
        RECT -70.205 27.715 -69.875 28.045 ;
        RECT -70.205 26.355 -69.875 26.685 ;
        RECT -70.205 24.995 -69.875 25.325 ;
        RECT -70.205 23.635 -69.875 23.965 ;
        RECT -70.205 22.275 -69.875 22.605 ;
        RECT -70.205 20.915 -69.875 21.245 ;
        RECT -70.205 19.555 -69.875 19.885 ;
        RECT -70.205 18.195 -69.875 18.525 ;
        RECT -70.205 16.835 -69.875 17.165 ;
        RECT -70.205 15.475 -69.875 15.805 ;
        RECT -70.205 14.115 -69.875 14.445 ;
        RECT -70.205 12.755 -69.875 13.085 ;
        RECT -70.205 11.395 -69.875 11.725 ;
        RECT -70.205 10.035 -69.875 10.365 ;
        RECT -70.205 8.675 -69.875 9.005 ;
        RECT -70.205 7.315 -69.875 7.645 ;
        RECT -70.205 5.955 -69.875 6.285 ;
        RECT -70.205 4.595 -69.875 4.925 ;
        RECT -70.205 3.235 -69.875 3.565 ;
        RECT -70.205 1.875 -69.875 2.205 ;
        RECT -70.205 0.515 -69.875 0.845 ;
        RECT -70.205 -0.845 -69.875 -0.515 ;
        RECT -70.205 -2.205 -69.875 -1.875 ;
        RECT -70.205 -3.565 -69.875 -3.235 ;
        RECT -70.205 -4.925 -69.875 -4.595 ;
        RECT -70.205 -6.285 -69.875 -5.955 ;
        RECT -70.205 -7.645 -69.875 -7.315 ;
        RECT -70.205 -9.005 -69.875 -8.675 ;
        RECT -70.205 -10.365 -69.875 -10.035 ;
        RECT -70.205 -11.725 -69.875 -11.395 ;
        RECT -70.205 -13.085 -69.875 -12.755 ;
        RECT -70.205 -14.445 -69.875 -14.115 ;
        RECT -70.205 -15.805 -69.875 -15.475 ;
        RECT -70.205 -17.165 -69.875 -16.835 ;
        RECT -70.205 -18.525 -69.875 -18.195 ;
        RECT -70.205 -19.885 -69.875 -19.555 ;
        RECT -70.205 -21.245 -69.875 -20.915 ;
        RECT -70.205 -22.605 -69.875 -22.275 ;
        RECT -70.205 -23.965 -69.875 -23.635 ;
        RECT -70.205 -25.325 -69.875 -24.995 ;
        RECT -70.205 -26.685 -69.875 -26.355 ;
        RECT -70.205 -28.045 -69.875 -27.715 ;
        RECT -70.205 -29.405 -69.875 -29.075 ;
        RECT -70.205 -30.765 -69.875 -30.435 ;
        RECT -70.205 -32.125 -69.875 -31.795 ;
        RECT -70.205 -33.485 -69.875 -33.155 ;
        RECT -70.205 -34.845 -69.875 -34.515 ;
        RECT -70.205 -36.205 -69.875 -35.875 ;
        RECT -70.205 -37.565 -69.875 -37.235 ;
        RECT -70.205 -38.925 -69.875 -38.595 ;
        RECT -70.205 -40.285 -69.875 -39.955 ;
        RECT -70.205 -41.645 -69.875 -41.315 ;
        RECT -70.205 -43.005 -69.875 -42.675 ;
        RECT -70.205 -44.365 -69.875 -44.035 ;
        RECT -70.205 -45.725 -69.875 -45.395 ;
        RECT -70.205 -47.085 -69.875 -46.755 ;
        RECT -70.205 -48.445 -69.875 -48.115 ;
        RECT -70.205 -49.805 -69.875 -49.475 ;
        RECT -70.205 -51.165 -69.875 -50.835 ;
        RECT -70.205 -52.525 -69.875 -52.195 ;
        RECT -70.205 -53.885 -69.875 -53.555 ;
        RECT -70.205 -55.245 -69.875 -54.915 ;
        RECT -70.205 -56.605 -69.875 -56.275 ;
        RECT -70.205 -57.965 -69.875 -57.635 ;
        RECT -70.205 -59.325 -69.875 -58.995 ;
        RECT -70.205 -60.685 -69.875 -60.355 ;
        RECT -70.205 -62.045 -69.875 -61.715 ;
        RECT -70.205 -63.405 -69.875 -63.075 ;
        RECT -70.205 -64.765 -69.875 -64.435 ;
        RECT -70.205 -66.125 -69.875 -65.795 ;
        RECT -70.205 -67.485 -69.875 -67.155 ;
        RECT -70.205 -68.845 -69.875 -68.515 ;
        RECT -70.205 -70.205 -69.875 -69.875 ;
        RECT -70.205 -71.565 -69.875 -71.235 ;
        RECT -70.205 -72.925 -69.875 -72.595 ;
        RECT -70.205 -74.285 -69.875 -73.955 ;
        RECT -70.205 -75.645 -69.875 -75.315 ;
        RECT -70.205 -77.005 -69.875 -76.675 ;
        RECT -70.205 -78.365 -69.875 -78.035 ;
        RECT -70.205 -79.725 -69.875 -79.395 ;
        RECT -70.205 -81.085 -69.875 -80.755 ;
        RECT -70.205 -82.445 -69.875 -82.115 ;
        RECT -70.205 -83.805 -69.875 -83.475 ;
        RECT -70.205 -85.165 -69.875 -84.835 ;
        RECT -70.205 -86.525 -69.875 -86.195 ;
        RECT -70.205 -87.885 -69.875 -87.555 ;
        RECT -70.205 -89.245 -69.875 -88.915 ;
        RECT -70.205 -90.605 -69.875 -90.275 ;
        RECT -70.205 -91.965 -69.875 -91.635 ;
        RECT -70.205 -93.325 -69.875 -92.995 ;
        RECT -70.205 -94.685 -69.875 -94.355 ;
        RECT -70.205 -96.045 -69.875 -95.715 ;
        RECT -70.205 -97.405 -69.875 -97.075 ;
        RECT -70.205 -98.765 -69.875 -98.435 ;
        RECT -70.205 -100.125 -69.875 -99.795 ;
        RECT -70.205 -101.485 -69.875 -101.155 ;
        RECT -70.205 -102.845 -69.875 -102.515 ;
        RECT -70.205 -104.205 -69.875 -103.875 ;
        RECT -70.205 -105.565 -69.875 -105.235 ;
        RECT -70.205 -106.925 -69.875 -106.595 ;
        RECT -70.205 -108.285 -69.875 -107.955 ;
        RECT -70.205 -109.645 -69.875 -109.315 ;
        RECT -70.205 -111.005 -69.875 -110.675 ;
        RECT -70.205 -112.365 -69.875 -112.035 ;
        RECT -70.205 -113.725 -69.875 -113.395 ;
        RECT -70.205 -115.085 -69.875 -114.755 ;
        RECT -70.205 -116.445 -69.875 -116.115 ;
        RECT -70.205 -117.805 -69.875 -117.475 ;
        RECT -70.205 -119.165 -69.875 -118.835 ;
        RECT -70.205 -120.525 -69.875 -120.195 ;
        RECT -70.205 -121.885 -69.875 -121.555 ;
        RECT -70.205 -123.245 -69.875 -122.915 ;
        RECT -70.205 -124.605 -69.875 -124.275 ;
        RECT -70.205 -125.965 -69.875 -125.635 ;
        RECT -70.205 -127.325 -69.875 -126.995 ;
        RECT -70.205 -128.685 -69.875 -128.355 ;
        RECT -70.205 -130.045 -69.875 -129.715 ;
        RECT -70.205 -131.405 -69.875 -131.075 ;
        RECT -70.205 -132.765 -69.875 -132.435 ;
        RECT -70.205 -134.125 -69.875 -133.795 ;
        RECT -70.205 -135.485 -69.875 -135.155 ;
        RECT -70.205 -136.845 -69.875 -136.515 ;
        RECT -70.205 -138.205 -69.875 -137.875 ;
        RECT -70.205 -139.565 -69.875 -139.235 ;
        RECT -70.205 -140.925 -69.875 -140.595 ;
        RECT -70.205 -142.285 -69.875 -141.955 ;
        RECT -70.205 -143.645 -69.875 -143.315 ;
        RECT -70.205 -145.005 -69.875 -144.675 ;
        RECT -70.205 -146.365 -69.875 -146.035 ;
        RECT -70.205 -147.725 -69.875 -147.395 ;
        RECT -70.205 -149.085 -69.875 -148.755 ;
        RECT -70.205 -150.445 -69.875 -150.115 ;
        RECT -70.205 -151.805 -69.875 -151.475 ;
        RECT -70.205 -153.165 -69.875 -152.835 ;
        RECT -70.205 -154.525 -69.875 -154.195 ;
        RECT -70.205 -155.885 -69.875 -155.555 ;
        RECT -70.205 -157.245 -69.875 -156.915 ;
        RECT -70.205 -158.605 -69.875 -158.275 ;
        RECT -70.205 -159.965 -69.875 -159.635 ;
        RECT -70.205 -161.325 -69.875 -160.995 ;
        RECT -70.205 -162.685 -69.875 -162.355 ;
        RECT -70.205 -164.045 -69.875 -163.715 ;
        RECT -70.205 -165.405 -69.875 -165.075 ;
        RECT -70.205 -166.765 -69.875 -166.435 ;
        RECT -70.205 -168.655 -69.875 -168.325 ;
        RECT -70.205 -169.485 -69.875 -169.155 ;
        RECT -70.205 -170.845 -69.875 -170.515 ;
        RECT -70.205 -173.565 -69.875 -173.235 ;
        RECT -70.205 -174.925 -69.875 -174.595 ;
        RECT -70.205 -177.645 -69.875 -177.315 ;
        RECT -70.205 -183.29 -69.875 -182.16 ;
        RECT -70.2 -183.405 -69.88 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -68.845 244.04 -68.515 245.17 ;
        RECT -68.845 239.875 -68.515 240.205 ;
        RECT -68.845 238.515 -68.515 238.845 ;
        RECT -68.845 237.155 -68.515 237.485 ;
        RECT -68.845 235.795 -68.515 236.125 ;
        RECT -68.845 234.435 -68.515 234.765 ;
        RECT -68.845 233.075 -68.515 233.405 ;
        RECT -68.845 231.715 -68.515 232.045 ;
        RECT -68.845 230.355 -68.515 230.685 ;
        RECT -68.845 228.995 -68.515 229.325 ;
        RECT -68.845 227.635 -68.515 227.965 ;
        RECT -68.845 226.275 -68.515 226.605 ;
        RECT -68.845 224.915 -68.515 225.245 ;
        RECT -68.845 223.555 -68.515 223.885 ;
        RECT -68.845 222.195 -68.515 222.525 ;
        RECT -68.845 220.835 -68.515 221.165 ;
        RECT -68.845 219.475 -68.515 219.805 ;
        RECT -68.845 218.115 -68.515 218.445 ;
        RECT -68.845 216.755 -68.515 217.085 ;
        RECT -68.845 215.395 -68.515 215.725 ;
        RECT -68.845 214.035 -68.515 214.365 ;
        RECT -68.845 212.675 -68.515 213.005 ;
        RECT -68.845 211.315 -68.515 211.645 ;
        RECT -68.845 209.955 -68.515 210.285 ;
        RECT -68.845 208.595 -68.515 208.925 ;
        RECT -68.845 207.235 -68.515 207.565 ;
        RECT -68.845 205.875 -68.515 206.205 ;
        RECT -68.845 204.515 -68.515 204.845 ;
        RECT -68.845 203.155 -68.515 203.485 ;
        RECT -68.845 201.795 -68.515 202.125 ;
        RECT -68.845 200.435 -68.515 200.765 ;
        RECT -68.845 199.075 -68.515 199.405 ;
        RECT -68.845 197.715 -68.515 198.045 ;
        RECT -68.845 196.355 -68.515 196.685 ;
        RECT -68.845 194.995 -68.515 195.325 ;
        RECT -68.845 193.635 -68.515 193.965 ;
        RECT -68.845 192.275 -68.515 192.605 ;
        RECT -68.845 190.915 -68.515 191.245 ;
        RECT -68.845 189.555 -68.515 189.885 ;
        RECT -68.845 188.195 -68.515 188.525 ;
        RECT -68.845 186.835 -68.515 187.165 ;
        RECT -68.845 185.475 -68.515 185.805 ;
        RECT -68.845 184.115 -68.515 184.445 ;
        RECT -68.845 182.755 -68.515 183.085 ;
        RECT -68.845 181.395 -68.515 181.725 ;
        RECT -68.845 180.035 -68.515 180.365 ;
        RECT -68.845 178.675 -68.515 179.005 ;
        RECT -68.845 177.315 -68.515 177.645 ;
        RECT -68.845 175.955 -68.515 176.285 ;
        RECT -68.845 174.595 -68.515 174.925 ;
        RECT -68.845 173.235 -68.515 173.565 ;
        RECT -68.845 171.875 -68.515 172.205 ;
        RECT -68.845 170.515 -68.515 170.845 ;
        RECT -68.845 169.155 -68.515 169.485 ;
        RECT -68.845 167.795 -68.515 168.125 ;
        RECT -68.845 166.435 -68.515 166.765 ;
        RECT -68.845 165.075 -68.515 165.405 ;
        RECT -68.845 163.715 -68.515 164.045 ;
        RECT -68.845 162.355 -68.515 162.685 ;
        RECT -68.845 160.995 -68.515 161.325 ;
        RECT -68.845 159.635 -68.515 159.965 ;
        RECT -68.845 158.275 -68.515 158.605 ;
        RECT -68.845 156.915 -68.515 157.245 ;
        RECT -68.845 155.555 -68.515 155.885 ;
        RECT -68.845 154.195 -68.515 154.525 ;
        RECT -68.845 152.835 -68.515 153.165 ;
        RECT -68.845 151.475 -68.515 151.805 ;
        RECT -68.845 150.115 -68.515 150.445 ;
        RECT -68.845 148.755 -68.515 149.085 ;
        RECT -68.845 147.395 -68.515 147.725 ;
        RECT -68.845 146.035 -68.515 146.365 ;
        RECT -68.845 144.675 -68.515 145.005 ;
        RECT -68.845 143.315 -68.515 143.645 ;
        RECT -68.845 141.955 -68.515 142.285 ;
        RECT -68.845 140.595 -68.515 140.925 ;
        RECT -68.845 139.235 -68.515 139.565 ;
        RECT -68.845 137.875 -68.515 138.205 ;
        RECT -68.845 136.515 -68.515 136.845 ;
        RECT -68.845 135.155 -68.515 135.485 ;
        RECT -68.845 133.795 -68.515 134.125 ;
        RECT -68.845 132.435 -68.515 132.765 ;
        RECT -68.845 131.075 -68.515 131.405 ;
        RECT -68.845 129.715 -68.515 130.045 ;
        RECT -68.845 128.355 -68.515 128.685 ;
        RECT -68.845 126.995 -68.515 127.325 ;
        RECT -68.845 125.635 -68.515 125.965 ;
        RECT -68.845 124.275 -68.515 124.605 ;
        RECT -68.845 122.915 -68.515 123.245 ;
        RECT -68.845 121.555 -68.515 121.885 ;
        RECT -68.845 120.195 -68.515 120.525 ;
        RECT -68.845 118.835 -68.515 119.165 ;
        RECT -68.845 117.475 -68.515 117.805 ;
        RECT -68.845 116.115 -68.515 116.445 ;
        RECT -68.845 114.755 -68.515 115.085 ;
        RECT -68.845 113.395 -68.515 113.725 ;
        RECT -68.845 112.035 -68.515 112.365 ;
        RECT -68.845 110.675 -68.515 111.005 ;
        RECT -68.845 109.315 -68.515 109.645 ;
        RECT -68.845 107.955 -68.515 108.285 ;
        RECT -68.845 106.595 -68.515 106.925 ;
        RECT -68.845 105.235 -68.515 105.565 ;
        RECT -68.845 103.875 -68.515 104.205 ;
        RECT -68.845 102.515 -68.515 102.845 ;
        RECT -68.845 101.155 -68.515 101.485 ;
        RECT -68.845 99.795 -68.515 100.125 ;
        RECT -68.845 98.435 -68.515 98.765 ;
        RECT -68.845 97.075 -68.515 97.405 ;
        RECT -68.845 95.715 -68.515 96.045 ;
        RECT -68.845 94.355 -68.515 94.685 ;
        RECT -68.845 92.995 -68.515 93.325 ;
        RECT -68.845 91.635 -68.515 91.965 ;
        RECT -68.845 90.275 -68.515 90.605 ;
        RECT -68.845 88.915 -68.515 89.245 ;
        RECT -68.845 87.555 -68.515 87.885 ;
        RECT -68.845 86.195 -68.515 86.525 ;
        RECT -68.845 84.835 -68.515 85.165 ;
        RECT -68.845 83.475 -68.515 83.805 ;
        RECT -68.845 82.115 -68.515 82.445 ;
        RECT -68.845 80.755 -68.515 81.085 ;
        RECT -68.845 79.395 -68.515 79.725 ;
        RECT -68.845 78.035 -68.515 78.365 ;
        RECT -68.845 76.675 -68.515 77.005 ;
        RECT -68.845 75.315 -68.515 75.645 ;
        RECT -68.845 73.955 -68.515 74.285 ;
        RECT -68.845 72.595 -68.515 72.925 ;
        RECT -68.845 71.235 -68.515 71.565 ;
        RECT -68.845 69.875 -68.515 70.205 ;
        RECT -68.845 68.515 -68.515 68.845 ;
        RECT -68.845 67.155 -68.515 67.485 ;
        RECT -68.845 65.795 -68.515 66.125 ;
        RECT -68.845 64.435 -68.515 64.765 ;
        RECT -68.845 63.075 -68.515 63.405 ;
        RECT -68.845 61.715 -68.515 62.045 ;
        RECT -68.845 60.355 -68.515 60.685 ;
        RECT -68.845 58.995 -68.515 59.325 ;
        RECT -68.845 57.635 -68.515 57.965 ;
        RECT -68.845 56.275 -68.515 56.605 ;
        RECT -68.845 54.915 -68.515 55.245 ;
        RECT -68.845 53.555 -68.515 53.885 ;
        RECT -68.845 52.195 -68.515 52.525 ;
        RECT -68.845 50.835 -68.515 51.165 ;
        RECT -68.845 49.475 -68.515 49.805 ;
        RECT -68.845 48.115 -68.515 48.445 ;
        RECT -68.845 46.755 -68.515 47.085 ;
        RECT -68.845 45.395 -68.515 45.725 ;
        RECT -68.845 44.035 -68.515 44.365 ;
        RECT -68.845 42.675 -68.515 43.005 ;
        RECT -68.845 41.315 -68.515 41.645 ;
        RECT -68.845 39.955 -68.515 40.285 ;
        RECT -68.845 38.595 -68.515 38.925 ;
        RECT -68.845 37.235 -68.515 37.565 ;
        RECT -68.845 35.875 -68.515 36.205 ;
        RECT -68.845 34.515 -68.515 34.845 ;
        RECT -68.845 33.155 -68.515 33.485 ;
        RECT -68.845 31.795 -68.515 32.125 ;
        RECT -68.845 30.435 -68.515 30.765 ;
        RECT -68.845 29.075 -68.515 29.405 ;
        RECT -68.845 27.715 -68.515 28.045 ;
        RECT -68.845 26.355 -68.515 26.685 ;
        RECT -68.845 24.995 -68.515 25.325 ;
        RECT -68.845 23.635 -68.515 23.965 ;
        RECT -68.845 22.275 -68.515 22.605 ;
        RECT -68.845 20.915 -68.515 21.245 ;
        RECT -68.845 19.555 -68.515 19.885 ;
        RECT -68.845 18.195 -68.515 18.525 ;
        RECT -68.845 16.835 -68.515 17.165 ;
        RECT -68.845 15.475 -68.515 15.805 ;
        RECT -68.845 14.115 -68.515 14.445 ;
        RECT -68.845 12.755 -68.515 13.085 ;
        RECT -68.845 11.395 -68.515 11.725 ;
        RECT -68.845 10.035 -68.515 10.365 ;
        RECT -68.845 8.675 -68.515 9.005 ;
        RECT -68.845 7.315 -68.515 7.645 ;
        RECT -68.845 5.955 -68.515 6.285 ;
        RECT -68.845 4.595 -68.515 4.925 ;
        RECT -68.845 3.235 -68.515 3.565 ;
        RECT -68.845 1.875 -68.515 2.205 ;
        RECT -68.845 0.515 -68.515 0.845 ;
        RECT -68.845 -0.845 -68.515 -0.515 ;
        RECT -68.845 -2.205 -68.515 -1.875 ;
        RECT -68.845 -3.565 -68.515 -3.235 ;
        RECT -68.845 -4.925 -68.515 -4.595 ;
        RECT -68.845 -6.285 -68.515 -5.955 ;
        RECT -68.845 -7.645 -68.515 -7.315 ;
        RECT -68.845 -9.005 -68.515 -8.675 ;
        RECT -68.845 -10.365 -68.515 -10.035 ;
        RECT -68.845 -11.725 -68.515 -11.395 ;
        RECT -68.845 -13.085 -68.515 -12.755 ;
        RECT -68.845 -14.445 -68.515 -14.115 ;
        RECT -68.845 -15.805 -68.515 -15.475 ;
        RECT -68.845 -17.165 -68.515 -16.835 ;
        RECT -68.845 -18.525 -68.515 -18.195 ;
        RECT -68.845 -19.885 -68.515 -19.555 ;
        RECT -68.845 -21.245 -68.515 -20.915 ;
        RECT -68.845 -22.605 -68.515 -22.275 ;
        RECT -68.845 -23.965 -68.515 -23.635 ;
        RECT -68.845 -25.325 -68.515 -24.995 ;
        RECT -68.845 -26.685 -68.515 -26.355 ;
        RECT -68.845 -28.045 -68.515 -27.715 ;
        RECT -68.845 -29.405 -68.515 -29.075 ;
        RECT -68.845 -30.765 -68.515 -30.435 ;
        RECT -68.845 -32.125 -68.515 -31.795 ;
        RECT -68.845 -33.485 -68.515 -33.155 ;
        RECT -68.845 -34.845 -68.515 -34.515 ;
        RECT -68.845 -36.205 -68.515 -35.875 ;
        RECT -68.845 -37.565 -68.515 -37.235 ;
        RECT -68.845 -38.925 -68.515 -38.595 ;
        RECT -68.845 -40.285 -68.515 -39.955 ;
        RECT -68.845 -41.645 -68.515 -41.315 ;
        RECT -68.845 -43.005 -68.515 -42.675 ;
        RECT -68.845 -44.365 -68.515 -44.035 ;
        RECT -68.845 -45.725 -68.515 -45.395 ;
        RECT -68.845 -47.085 -68.515 -46.755 ;
        RECT -68.845 -48.445 -68.515 -48.115 ;
        RECT -68.845 -49.805 -68.515 -49.475 ;
        RECT -68.845 -51.165 -68.515 -50.835 ;
        RECT -68.845 -52.525 -68.515 -52.195 ;
        RECT -68.845 -53.885 -68.515 -53.555 ;
        RECT -68.845 -55.245 -68.515 -54.915 ;
        RECT -68.845 -56.605 -68.515 -56.275 ;
        RECT -68.845 -57.965 -68.515 -57.635 ;
        RECT -68.845 -59.325 -68.515 -58.995 ;
        RECT -68.845 -60.685 -68.515 -60.355 ;
        RECT -68.845 -62.045 -68.515 -61.715 ;
        RECT -68.845 -63.405 -68.515 -63.075 ;
        RECT -68.845 -64.765 -68.515 -64.435 ;
        RECT -68.845 -66.125 -68.515 -65.795 ;
        RECT -68.845 -67.485 -68.515 -67.155 ;
        RECT -68.845 -68.845 -68.515 -68.515 ;
        RECT -68.845 -70.205 -68.515 -69.875 ;
        RECT -68.845 -71.565 -68.515 -71.235 ;
        RECT -68.845 -72.925 -68.515 -72.595 ;
        RECT -68.845 -74.285 -68.515 -73.955 ;
        RECT -68.845 -75.645 -68.515 -75.315 ;
        RECT -68.845 -77.005 -68.515 -76.675 ;
        RECT -68.845 -78.365 -68.515 -78.035 ;
        RECT -68.845 -79.725 -68.515 -79.395 ;
        RECT -68.845 -81.085 -68.515 -80.755 ;
        RECT -68.845 -82.445 -68.515 -82.115 ;
        RECT -68.845 -83.805 -68.515 -83.475 ;
        RECT -68.845 -85.165 -68.515 -84.835 ;
        RECT -68.845 -86.525 -68.515 -86.195 ;
        RECT -68.845 -87.885 -68.515 -87.555 ;
        RECT -68.845 -89.245 -68.515 -88.915 ;
        RECT -68.845 -90.605 -68.515 -90.275 ;
        RECT -68.845 -91.965 -68.515 -91.635 ;
        RECT -68.845 -93.325 -68.515 -92.995 ;
        RECT -68.845 -94.685 -68.515 -94.355 ;
        RECT -68.845 -96.045 -68.515 -95.715 ;
        RECT -68.845 -97.405 -68.515 -97.075 ;
        RECT -68.845 -98.765 -68.515 -98.435 ;
        RECT -68.845 -100.125 -68.515 -99.795 ;
        RECT -68.845 -101.485 -68.515 -101.155 ;
        RECT -68.845 -102.845 -68.515 -102.515 ;
        RECT -68.845 -104.205 -68.515 -103.875 ;
        RECT -68.845 -105.565 -68.515 -105.235 ;
        RECT -68.845 -106.925 -68.515 -106.595 ;
        RECT -68.845 -108.285 -68.515 -107.955 ;
        RECT -68.845 -109.645 -68.515 -109.315 ;
        RECT -68.845 -111.005 -68.515 -110.675 ;
        RECT -68.845 -112.365 -68.515 -112.035 ;
        RECT -68.845 -113.725 -68.515 -113.395 ;
        RECT -68.845 -115.085 -68.515 -114.755 ;
        RECT -68.845 -116.445 -68.515 -116.115 ;
        RECT -68.845 -117.805 -68.515 -117.475 ;
        RECT -68.845 -119.165 -68.515 -118.835 ;
        RECT -68.845 -120.525 -68.515 -120.195 ;
        RECT -68.845 -121.885 -68.515 -121.555 ;
        RECT -68.845 -123.245 -68.515 -122.915 ;
        RECT -68.845 -124.605 -68.515 -124.275 ;
        RECT -68.845 -125.965 -68.515 -125.635 ;
        RECT -68.845 -127.325 -68.515 -126.995 ;
        RECT -68.845 -128.685 -68.515 -128.355 ;
        RECT -68.845 -130.045 -68.515 -129.715 ;
        RECT -68.845 -131.405 -68.515 -131.075 ;
        RECT -68.845 -132.765 -68.515 -132.435 ;
        RECT -68.845 -134.125 -68.515 -133.795 ;
        RECT -68.845 -135.485 -68.515 -135.155 ;
        RECT -68.845 -136.845 -68.515 -136.515 ;
        RECT -68.845 -138.205 -68.515 -137.875 ;
        RECT -68.845 -139.565 -68.515 -139.235 ;
        RECT -68.845 -140.925 -68.515 -140.595 ;
        RECT -68.845 -142.285 -68.515 -141.955 ;
        RECT -68.845 -143.645 -68.515 -143.315 ;
        RECT -68.845 -145.005 -68.515 -144.675 ;
        RECT -68.845 -146.365 -68.515 -146.035 ;
        RECT -68.845 -147.725 -68.515 -147.395 ;
        RECT -68.845 -149.085 -68.515 -148.755 ;
        RECT -68.845 -150.445 -68.515 -150.115 ;
        RECT -68.845 -151.805 -68.515 -151.475 ;
        RECT -68.845 -153.165 -68.515 -152.835 ;
        RECT -68.845 -154.525 -68.515 -154.195 ;
        RECT -68.845 -155.885 -68.515 -155.555 ;
        RECT -68.845 -157.245 -68.515 -156.915 ;
        RECT -68.845 -158.605 -68.515 -158.275 ;
        RECT -68.845 -159.965 -68.515 -159.635 ;
        RECT -68.845 -161.325 -68.515 -160.995 ;
        RECT -68.845 -162.685 -68.515 -162.355 ;
        RECT -68.845 -164.045 -68.515 -163.715 ;
        RECT -68.845 -165.405 -68.515 -165.075 ;
        RECT -68.845 -166.765 -68.515 -166.435 ;
        RECT -68.845 -168.655 -68.515 -168.325 ;
        RECT -68.845 -169.485 -68.515 -169.155 ;
        RECT -68.845 -170.845 -68.515 -170.515 ;
        RECT -68.845 -172.205 -68.515 -171.875 ;
        RECT -68.845 -173.565 -68.515 -173.235 ;
        RECT -68.845 -174.925 -68.515 -174.595 ;
        RECT -68.845 -177.645 -68.515 -177.315 ;
        RECT -68.845 -183.29 -68.515 -182.16 ;
        RECT -68.84 -183.405 -68.52 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -67.485 79.395 -67.155 79.725 ;
        RECT -67.485 78.035 -67.155 78.365 ;
        RECT -67.485 76.675 -67.155 77.005 ;
        RECT -67.485 75.315 -67.155 75.645 ;
        RECT -67.485 73.955 -67.155 74.285 ;
        RECT -67.485 72.595 -67.155 72.925 ;
        RECT -67.485 71.235 -67.155 71.565 ;
        RECT -67.485 69.875 -67.155 70.205 ;
        RECT -67.485 68.515 -67.155 68.845 ;
        RECT -67.485 67.155 -67.155 67.485 ;
        RECT -67.485 65.795 -67.155 66.125 ;
        RECT -67.485 64.435 -67.155 64.765 ;
        RECT -67.485 63.075 -67.155 63.405 ;
        RECT -67.485 61.715 -67.155 62.045 ;
        RECT -67.485 60.355 -67.155 60.685 ;
        RECT -67.485 58.995 -67.155 59.325 ;
        RECT -67.485 57.635 -67.155 57.965 ;
        RECT -67.485 56.275 -67.155 56.605 ;
        RECT -67.485 54.915 -67.155 55.245 ;
        RECT -67.485 53.555 -67.155 53.885 ;
        RECT -67.485 52.195 -67.155 52.525 ;
        RECT -67.485 50.835 -67.155 51.165 ;
        RECT -67.485 49.475 -67.155 49.805 ;
        RECT -67.485 48.115 -67.155 48.445 ;
        RECT -67.485 46.755 -67.155 47.085 ;
        RECT -67.485 45.395 -67.155 45.725 ;
        RECT -67.485 44.035 -67.155 44.365 ;
        RECT -67.485 42.675 -67.155 43.005 ;
        RECT -67.485 41.315 -67.155 41.645 ;
        RECT -67.485 39.955 -67.155 40.285 ;
        RECT -67.485 38.595 -67.155 38.925 ;
        RECT -67.485 37.235 -67.155 37.565 ;
        RECT -67.485 35.875 -67.155 36.205 ;
        RECT -67.485 34.515 -67.155 34.845 ;
        RECT -67.485 33.155 -67.155 33.485 ;
        RECT -67.485 31.795 -67.155 32.125 ;
        RECT -67.485 30.435 -67.155 30.765 ;
        RECT -67.485 29.075 -67.155 29.405 ;
        RECT -67.485 27.715 -67.155 28.045 ;
        RECT -67.485 26.355 -67.155 26.685 ;
        RECT -67.485 24.995 -67.155 25.325 ;
        RECT -67.485 23.635 -67.155 23.965 ;
        RECT -67.485 22.275 -67.155 22.605 ;
        RECT -67.485 20.915 -67.155 21.245 ;
        RECT -67.485 19.555 -67.155 19.885 ;
        RECT -67.485 18.195 -67.155 18.525 ;
        RECT -67.485 16.835 -67.155 17.165 ;
        RECT -67.485 15.475 -67.155 15.805 ;
        RECT -67.485 14.115 -67.155 14.445 ;
        RECT -67.485 12.755 -67.155 13.085 ;
        RECT -67.485 11.395 -67.155 11.725 ;
        RECT -67.485 10.035 -67.155 10.365 ;
        RECT -67.485 8.675 -67.155 9.005 ;
        RECT -67.485 7.315 -67.155 7.645 ;
        RECT -67.485 5.955 -67.155 6.285 ;
        RECT -67.485 4.595 -67.155 4.925 ;
        RECT -67.485 3.235 -67.155 3.565 ;
        RECT -67.485 1.875 -67.155 2.205 ;
        RECT -67.485 0.515 -67.155 0.845 ;
        RECT -67.485 -0.845 -67.155 -0.515 ;
        RECT -67.485 -2.205 -67.155 -1.875 ;
        RECT -67.485 -3.565 -67.155 -3.235 ;
        RECT -67.485 -4.925 -67.155 -4.595 ;
        RECT -67.485 -6.285 -67.155 -5.955 ;
        RECT -67.485 -7.645 -67.155 -7.315 ;
        RECT -67.485 -9.005 -67.155 -8.675 ;
        RECT -67.485 -10.365 -67.155 -10.035 ;
        RECT -67.485 -11.725 -67.155 -11.395 ;
        RECT -67.485 -13.085 -67.155 -12.755 ;
        RECT -67.485 -14.445 -67.155 -14.115 ;
        RECT -67.485 -15.805 -67.155 -15.475 ;
        RECT -67.485 -17.165 -67.155 -16.835 ;
        RECT -67.485 -18.525 -67.155 -18.195 ;
        RECT -67.485 -19.885 -67.155 -19.555 ;
        RECT -67.485 -21.245 -67.155 -20.915 ;
        RECT -67.485 -22.605 -67.155 -22.275 ;
        RECT -67.485 -23.965 -67.155 -23.635 ;
        RECT -67.485 -25.325 -67.155 -24.995 ;
        RECT -67.485 -26.685 -67.155 -26.355 ;
        RECT -67.485 -28.045 -67.155 -27.715 ;
        RECT -67.485 -29.405 -67.155 -29.075 ;
        RECT -67.485 -30.765 -67.155 -30.435 ;
        RECT -67.485 -32.125 -67.155 -31.795 ;
        RECT -67.485 -33.485 -67.155 -33.155 ;
        RECT -67.485 -34.845 -67.155 -34.515 ;
        RECT -67.485 -36.205 -67.155 -35.875 ;
        RECT -67.485 -37.565 -67.155 -37.235 ;
        RECT -67.485 -38.925 -67.155 -38.595 ;
        RECT -67.485 -40.285 -67.155 -39.955 ;
        RECT -67.485 -41.645 -67.155 -41.315 ;
        RECT -67.485 -43.005 -67.155 -42.675 ;
        RECT -67.485 -44.365 -67.155 -44.035 ;
        RECT -67.485 -45.725 -67.155 -45.395 ;
        RECT -67.485 -47.085 -67.155 -46.755 ;
        RECT -67.485 -48.445 -67.155 -48.115 ;
        RECT -67.485 -49.805 -67.155 -49.475 ;
        RECT -67.485 -51.165 -67.155 -50.835 ;
        RECT -67.485 -52.525 -67.155 -52.195 ;
        RECT -67.485 -53.885 -67.155 -53.555 ;
        RECT -67.485 -55.245 -67.155 -54.915 ;
        RECT -67.485 -56.605 -67.155 -56.275 ;
        RECT -67.485 -57.965 -67.155 -57.635 ;
        RECT -67.485 -59.325 -67.155 -58.995 ;
        RECT -67.485 -60.685 -67.155 -60.355 ;
        RECT -67.485 -62.045 -67.155 -61.715 ;
        RECT -67.485 -63.405 -67.155 -63.075 ;
        RECT -67.485 -64.765 -67.155 -64.435 ;
        RECT -67.485 -66.125 -67.155 -65.795 ;
        RECT -67.485 -67.485 -67.155 -67.155 ;
        RECT -67.485 -68.845 -67.155 -68.515 ;
        RECT -67.485 -70.205 -67.155 -69.875 ;
        RECT -67.485 -71.565 -67.155 -71.235 ;
        RECT -67.485 -72.925 -67.155 -72.595 ;
        RECT -67.485 -74.285 -67.155 -73.955 ;
        RECT -67.485 -75.645 -67.155 -75.315 ;
        RECT -67.485 -77.005 -67.155 -76.675 ;
        RECT -67.485 -78.365 -67.155 -78.035 ;
        RECT -67.485 -79.725 -67.155 -79.395 ;
        RECT -67.485 -81.085 -67.155 -80.755 ;
        RECT -67.485 -82.445 -67.155 -82.115 ;
        RECT -67.485 -83.805 -67.155 -83.475 ;
        RECT -67.485 -85.165 -67.155 -84.835 ;
        RECT -67.485 -86.525 -67.155 -86.195 ;
        RECT -67.485 -87.885 -67.155 -87.555 ;
        RECT -67.485 -89.245 -67.155 -88.915 ;
        RECT -67.485 -90.605 -67.155 -90.275 ;
        RECT -67.485 -91.965 -67.155 -91.635 ;
        RECT -67.485 -93.325 -67.155 -92.995 ;
        RECT -67.485 -94.685 -67.155 -94.355 ;
        RECT -67.485 -96.045 -67.155 -95.715 ;
        RECT -67.485 -97.405 -67.155 -97.075 ;
        RECT -67.485 -98.765 -67.155 -98.435 ;
        RECT -67.485 -100.125 -67.155 -99.795 ;
        RECT -67.485 -101.485 -67.155 -101.155 ;
        RECT -67.485 -102.845 -67.155 -102.515 ;
        RECT -67.485 -104.205 -67.155 -103.875 ;
        RECT -67.485 -105.565 -67.155 -105.235 ;
        RECT -67.485 -106.925 -67.155 -106.595 ;
        RECT -67.485 -108.285 -67.155 -107.955 ;
        RECT -67.485 -109.645 -67.155 -109.315 ;
        RECT -67.485 -111.005 -67.155 -110.675 ;
        RECT -67.485 -112.365 -67.155 -112.035 ;
        RECT -67.485 -113.725 -67.155 -113.395 ;
        RECT -67.485 -115.085 -67.155 -114.755 ;
        RECT -67.485 -116.445 -67.155 -116.115 ;
        RECT -67.485 -117.805 -67.155 -117.475 ;
        RECT -67.485 -119.165 -67.155 -118.835 ;
        RECT -67.485 -120.525 -67.155 -120.195 ;
        RECT -67.485 -121.885 -67.155 -121.555 ;
        RECT -67.485 -123.245 -67.155 -122.915 ;
        RECT -67.485 -124.605 -67.155 -124.275 ;
        RECT -67.485 -125.965 -67.155 -125.635 ;
        RECT -67.485 -127.325 -67.155 -126.995 ;
        RECT -67.485 -128.685 -67.155 -128.355 ;
        RECT -67.485 -130.045 -67.155 -129.715 ;
        RECT -67.485 -131.405 -67.155 -131.075 ;
        RECT -67.485 -132.765 -67.155 -132.435 ;
        RECT -67.485 -134.125 -67.155 -133.795 ;
        RECT -67.485 -135.485 -67.155 -135.155 ;
        RECT -67.485 -136.845 -67.155 -136.515 ;
        RECT -67.485 -138.205 -67.155 -137.875 ;
        RECT -67.485 -139.565 -67.155 -139.235 ;
        RECT -67.485 -140.925 -67.155 -140.595 ;
        RECT -67.485 -142.285 -67.155 -141.955 ;
        RECT -67.485 -143.645 -67.155 -143.315 ;
        RECT -67.485 -145.005 -67.155 -144.675 ;
        RECT -67.485 -146.365 -67.155 -146.035 ;
        RECT -67.485 -147.725 -67.155 -147.395 ;
        RECT -67.485 -149.085 -67.155 -148.755 ;
        RECT -67.485 -150.445 -67.155 -150.115 ;
        RECT -67.485 -151.805 -67.155 -151.475 ;
        RECT -67.485 -153.165 -67.155 -152.835 ;
        RECT -67.485 -154.525 -67.155 -154.195 ;
        RECT -67.485 -155.885 -67.155 -155.555 ;
        RECT -67.485 -157.245 -67.155 -156.915 ;
        RECT -67.485 -158.605 -67.155 -158.275 ;
        RECT -67.485 -159.965 -67.155 -159.635 ;
        RECT -67.485 -161.325 -67.155 -160.995 ;
        RECT -67.485 -162.685 -67.155 -162.355 ;
        RECT -67.485 -164.045 -67.155 -163.715 ;
        RECT -67.485 -165.405 -67.155 -165.075 ;
        RECT -67.485 -166.765 -67.155 -166.435 ;
        RECT -67.485 -168.655 -67.155 -168.325 ;
        RECT -67.485 -169.485 -67.155 -169.155 ;
        RECT -67.485 -170.845 -67.155 -170.515 ;
        RECT -67.485 -172.205 -67.155 -171.875 ;
        RECT -67.485 -174.925 -67.155 -174.595 ;
        RECT -67.485 -177.645 -67.155 -177.315 ;
        RECT -67.485 -183.29 -67.155 -182.16 ;
        RECT -67.48 -183.405 -67.16 245.285 ;
        RECT -67.485 244.04 -67.155 245.17 ;
        RECT -67.485 239.875 -67.155 240.205 ;
        RECT -67.485 238.515 -67.155 238.845 ;
        RECT -67.485 237.155 -67.155 237.485 ;
        RECT -67.485 235.795 -67.155 236.125 ;
        RECT -67.485 234.435 -67.155 234.765 ;
        RECT -67.485 233.075 -67.155 233.405 ;
        RECT -67.485 231.715 -67.155 232.045 ;
        RECT -67.485 230.355 -67.155 230.685 ;
        RECT -67.485 228.995 -67.155 229.325 ;
        RECT -67.485 227.635 -67.155 227.965 ;
        RECT -67.485 226.275 -67.155 226.605 ;
        RECT -67.485 224.915 -67.155 225.245 ;
        RECT -67.485 223.555 -67.155 223.885 ;
        RECT -67.485 222.195 -67.155 222.525 ;
        RECT -67.485 220.835 -67.155 221.165 ;
        RECT -67.485 219.475 -67.155 219.805 ;
        RECT -67.485 218.115 -67.155 218.445 ;
        RECT -67.485 216.755 -67.155 217.085 ;
        RECT -67.485 215.395 -67.155 215.725 ;
        RECT -67.485 214.035 -67.155 214.365 ;
        RECT -67.485 212.675 -67.155 213.005 ;
        RECT -67.485 211.315 -67.155 211.645 ;
        RECT -67.485 209.955 -67.155 210.285 ;
        RECT -67.485 208.595 -67.155 208.925 ;
        RECT -67.485 207.235 -67.155 207.565 ;
        RECT -67.485 205.875 -67.155 206.205 ;
        RECT -67.485 204.515 -67.155 204.845 ;
        RECT -67.485 203.155 -67.155 203.485 ;
        RECT -67.485 201.795 -67.155 202.125 ;
        RECT -67.485 200.435 -67.155 200.765 ;
        RECT -67.485 199.075 -67.155 199.405 ;
        RECT -67.485 197.715 -67.155 198.045 ;
        RECT -67.485 196.355 -67.155 196.685 ;
        RECT -67.485 194.995 -67.155 195.325 ;
        RECT -67.485 193.635 -67.155 193.965 ;
        RECT -67.485 192.275 -67.155 192.605 ;
        RECT -67.485 190.915 -67.155 191.245 ;
        RECT -67.485 189.555 -67.155 189.885 ;
        RECT -67.485 188.195 -67.155 188.525 ;
        RECT -67.485 186.835 -67.155 187.165 ;
        RECT -67.485 185.475 -67.155 185.805 ;
        RECT -67.485 184.115 -67.155 184.445 ;
        RECT -67.485 182.755 -67.155 183.085 ;
        RECT -67.485 181.395 -67.155 181.725 ;
        RECT -67.485 180.035 -67.155 180.365 ;
        RECT -67.485 178.675 -67.155 179.005 ;
        RECT -67.485 177.315 -67.155 177.645 ;
        RECT -67.485 175.955 -67.155 176.285 ;
        RECT -67.485 174.595 -67.155 174.925 ;
        RECT -67.485 173.235 -67.155 173.565 ;
        RECT -67.485 171.875 -67.155 172.205 ;
        RECT -67.485 170.515 -67.155 170.845 ;
        RECT -67.485 169.155 -67.155 169.485 ;
        RECT -67.485 167.795 -67.155 168.125 ;
        RECT -67.485 166.435 -67.155 166.765 ;
        RECT -67.485 165.075 -67.155 165.405 ;
        RECT -67.485 163.715 -67.155 164.045 ;
        RECT -67.485 162.355 -67.155 162.685 ;
        RECT -67.485 160.995 -67.155 161.325 ;
        RECT -67.485 159.635 -67.155 159.965 ;
        RECT -67.485 158.275 -67.155 158.605 ;
        RECT -67.485 156.915 -67.155 157.245 ;
        RECT -67.485 155.555 -67.155 155.885 ;
        RECT -67.485 154.195 -67.155 154.525 ;
        RECT -67.485 152.835 -67.155 153.165 ;
        RECT -67.485 151.475 -67.155 151.805 ;
        RECT -67.485 150.115 -67.155 150.445 ;
        RECT -67.485 148.755 -67.155 149.085 ;
        RECT -67.485 147.395 -67.155 147.725 ;
        RECT -67.485 146.035 -67.155 146.365 ;
        RECT -67.485 144.675 -67.155 145.005 ;
        RECT -67.485 143.315 -67.155 143.645 ;
        RECT -67.485 141.955 -67.155 142.285 ;
        RECT -67.485 140.595 -67.155 140.925 ;
        RECT -67.485 139.235 -67.155 139.565 ;
        RECT -67.485 137.875 -67.155 138.205 ;
        RECT -67.485 136.515 -67.155 136.845 ;
        RECT -67.485 135.155 -67.155 135.485 ;
        RECT -67.485 133.795 -67.155 134.125 ;
        RECT -67.485 132.435 -67.155 132.765 ;
        RECT -67.485 131.075 -67.155 131.405 ;
        RECT -67.485 129.715 -67.155 130.045 ;
        RECT -67.485 128.355 -67.155 128.685 ;
        RECT -67.485 126.995 -67.155 127.325 ;
        RECT -67.485 125.635 -67.155 125.965 ;
        RECT -67.485 124.275 -67.155 124.605 ;
        RECT -67.485 122.915 -67.155 123.245 ;
        RECT -67.485 121.555 -67.155 121.885 ;
        RECT -67.485 120.195 -67.155 120.525 ;
        RECT -67.485 118.835 -67.155 119.165 ;
        RECT -67.485 117.475 -67.155 117.805 ;
        RECT -67.485 116.115 -67.155 116.445 ;
        RECT -67.485 114.755 -67.155 115.085 ;
        RECT -67.485 113.395 -67.155 113.725 ;
        RECT -67.485 112.035 -67.155 112.365 ;
        RECT -67.485 110.675 -67.155 111.005 ;
        RECT -67.485 109.315 -67.155 109.645 ;
        RECT -67.485 107.955 -67.155 108.285 ;
        RECT -67.485 106.595 -67.155 106.925 ;
        RECT -67.485 105.235 -67.155 105.565 ;
        RECT -67.485 103.875 -67.155 104.205 ;
        RECT -67.485 102.515 -67.155 102.845 ;
        RECT -67.485 101.155 -67.155 101.485 ;
        RECT -67.485 99.795 -67.155 100.125 ;
        RECT -67.485 98.435 -67.155 98.765 ;
        RECT -67.485 97.075 -67.155 97.405 ;
        RECT -67.485 95.715 -67.155 96.045 ;
        RECT -67.485 94.355 -67.155 94.685 ;
        RECT -67.485 92.995 -67.155 93.325 ;
        RECT -67.485 91.635 -67.155 91.965 ;
        RECT -67.485 90.275 -67.155 90.605 ;
        RECT -67.485 88.915 -67.155 89.245 ;
        RECT -67.485 87.555 -67.155 87.885 ;
        RECT -67.485 86.195 -67.155 86.525 ;
        RECT -67.485 84.835 -67.155 85.165 ;
        RECT -67.485 83.475 -67.155 83.805 ;
        RECT -67.485 82.115 -67.155 82.445 ;
        RECT -67.485 80.755 -67.155 81.085 ;
    END
    PORT
      LAYER met3 ;
        RECT -74.285 244.04 -73.955 245.17 ;
        RECT -74.285 239.875 -73.955 240.205 ;
        RECT -74.285 238.515 -73.955 238.845 ;
        RECT -74.285 237.155 -73.955 237.485 ;
        RECT -74.285 235.795 -73.955 236.125 ;
        RECT -74.285 234.435 -73.955 234.765 ;
        RECT -74.285 233.075 -73.955 233.405 ;
        RECT -74.285 231.715 -73.955 232.045 ;
        RECT -74.285 230.355 -73.955 230.685 ;
        RECT -74.285 228.995 -73.955 229.325 ;
        RECT -74.285 227.635 -73.955 227.965 ;
        RECT -74.285 226.275 -73.955 226.605 ;
        RECT -74.285 224.915 -73.955 225.245 ;
        RECT -74.285 223.555 -73.955 223.885 ;
        RECT -74.285 222.195 -73.955 222.525 ;
        RECT -74.285 220.835 -73.955 221.165 ;
        RECT -74.285 219.475 -73.955 219.805 ;
        RECT -74.285 218.115 -73.955 218.445 ;
        RECT -74.285 216.755 -73.955 217.085 ;
        RECT -74.285 215.395 -73.955 215.725 ;
        RECT -74.285 214.035 -73.955 214.365 ;
        RECT -74.285 212.675 -73.955 213.005 ;
        RECT -74.285 211.315 -73.955 211.645 ;
        RECT -74.285 209.955 -73.955 210.285 ;
        RECT -74.285 208.595 -73.955 208.925 ;
        RECT -74.285 207.235 -73.955 207.565 ;
        RECT -74.285 205.875 -73.955 206.205 ;
        RECT -74.285 204.515 -73.955 204.845 ;
        RECT -74.285 203.155 -73.955 203.485 ;
        RECT -74.285 201.795 -73.955 202.125 ;
        RECT -74.285 200.435 -73.955 200.765 ;
        RECT -74.285 199.075 -73.955 199.405 ;
        RECT -74.285 197.715 -73.955 198.045 ;
        RECT -74.285 196.355 -73.955 196.685 ;
        RECT -74.285 194.995 -73.955 195.325 ;
        RECT -74.285 193.635 -73.955 193.965 ;
        RECT -74.285 192.275 -73.955 192.605 ;
        RECT -74.285 190.915 -73.955 191.245 ;
        RECT -74.285 189.555 -73.955 189.885 ;
        RECT -74.285 188.195 -73.955 188.525 ;
        RECT -74.285 186.835 -73.955 187.165 ;
        RECT -74.285 185.475 -73.955 185.805 ;
        RECT -74.285 184.115 -73.955 184.445 ;
        RECT -74.285 182.755 -73.955 183.085 ;
        RECT -74.285 181.395 -73.955 181.725 ;
        RECT -74.285 180.035 -73.955 180.365 ;
        RECT -74.285 178.675 -73.955 179.005 ;
        RECT -74.285 177.315 -73.955 177.645 ;
        RECT -74.285 175.955 -73.955 176.285 ;
        RECT -74.285 174.595 -73.955 174.925 ;
        RECT -74.285 173.235 -73.955 173.565 ;
        RECT -74.285 171.875 -73.955 172.205 ;
        RECT -74.285 170.515 -73.955 170.845 ;
        RECT -74.285 169.155 -73.955 169.485 ;
        RECT -74.285 167.795 -73.955 168.125 ;
        RECT -74.285 166.435 -73.955 166.765 ;
        RECT -74.285 165.075 -73.955 165.405 ;
        RECT -74.285 163.715 -73.955 164.045 ;
        RECT -74.285 162.355 -73.955 162.685 ;
        RECT -74.285 160.995 -73.955 161.325 ;
        RECT -74.285 159.635 -73.955 159.965 ;
        RECT -74.285 158.275 -73.955 158.605 ;
        RECT -74.285 156.915 -73.955 157.245 ;
        RECT -74.285 155.555 -73.955 155.885 ;
        RECT -74.285 154.195 -73.955 154.525 ;
        RECT -74.285 152.835 -73.955 153.165 ;
        RECT -74.285 151.475 -73.955 151.805 ;
        RECT -74.285 150.115 -73.955 150.445 ;
        RECT -74.285 148.755 -73.955 149.085 ;
        RECT -74.285 147.395 -73.955 147.725 ;
        RECT -74.285 146.035 -73.955 146.365 ;
        RECT -74.285 144.675 -73.955 145.005 ;
        RECT -74.285 143.315 -73.955 143.645 ;
        RECT -74.285 141.955 -73.955 142.285 ;
        RECT -74.285 140.595 -73.955 140.925 ;
        RECT -74.285 139.235 -73.955 139.565 ;
        RECT -74.285 137.875 -73.955 138.205 ;
        RECT -74.285 136.515 -73.955 136.845 ;
        RECT -74.285 135.155 -73.955 135.485 ;
        RECT -74.285 133.795 -73.955 134.125 ;
        RECT -74.285 132.435 -73.955 132.765 ;
        RECT -74.285 131.075 -73.955 131.405 ;
        RECT -74.285 129.715 -73.955 130.045 ;
        RECT -74.285 128.355 -73.955 128.685 ;
        RECT -74.285 126.995 -73.955 127.325 ;
        RECT -74.285 125.635 -73.955 125.965 ;
        RECT -74.285 124.275 -73.955 124.605 ;
        RECT -74.285 122.915 -73.955 123.245 ;
        RECT -74.285 121.555 -73.955 121.885 ;
        RECT -74.285 120.195 -73.955 120.525 ;
        RECT -74.285 118.835 -73.955 119.165 ;
        RECT -74.285 117.475 -73.955 117.805 ;
        RECT -74.285 116.115 -73.955 116.445 ;
        RECT -74.285 114.755 -73.955 115.085 ;
        RECT -74.285 113.395 -73.955 113.725 ;
        RECT -74.285 112.035 -73.955 112.365 ;
        RECT -74.285 110.675 -73.955 111.005 ;
        RECT -74.285 109.315 -73.955 109.645 ;
        RECT -74.285 107.955 -73.955 108.285 ;
        RECT -74.285 106.595 -73.955 106.925 ;
        RECT -74.285 105.235 -73.955 105.565 ;
        RECT -74.285 103.875 -73.955 104.205 ;
        RECT -74.285 102.515 -73.955 102.845 ;
        RECT -74.285 101.155 -73.955 101.485 ;
        RECT -74.285 99.795 -73.955 100.125 ;
        RECT -74.285 98.435 -73.955 98.765 ;
        RECT -74.285 97.075 -73.955 97.405 ;
        RECT -74.285 95.715 -73.955 96.045 ;
        RECT -74.285 94.355 -73.955 94.685 ;
        RECT -74.285 92.995 -73.955 93.325 ;
        RECT -74.285 91.635 -73.955 91.965 ;
        RECT -74.285 90.275 -73.955 90.605 ;
        RECT -74.285 88.915 -73.955 89.245 ;
        RECT -74.285 87.555 -73.955 87.885 ;
        RECT -74.285 86.195 -73.955 86.525 ;
        RECT -74.285 84.835 -73.955 85.165 ;
        RECT -74.285 83.475 -73.955 83.805 ;
        RECT -74.285 82.115 -73.955 82.445 ;
        RECT -74.285 80.755 -73.955 81.085 ;
        RECT -74.285 79.395 -73.955 79.725 ;
        RECT -74.285 78.035 -73.955 78.365 ;
        RECT -74.285 76.675 -73.955 77.005 ;
        RECT -74.285 75.315 -73.955 75.645 ;
        RECT -74.285 73.955 -73.955 74.285 ;
        RECT -74.285 72.595 -73.955 72.925 ;
        RECT -74.285 71.235 -73.955 71.565 ;
        RECT -74.285 69.875 -73.955 70.205 ;
        RECT -74.285 68.515 -73.955 68.845 ;
        RECT -74.285 67.155 -73.955 67.485 ;
        RECT -74.285 65.795 -73.955 66.125 ;
        RECT -74.285 64.435 -73.955 64.765 ;
        RECT -74.285 63.075 -73.955 63.405 ;
        RECT -74.285 61.715 -73.955 62.045 ;
        RECT -74.285 60.355 -73.955 60.685 ;
        RECT -74.285 58.995 -73.955 59.325 ;
        RECT -74.285 57.635 -73.955 57.965 ;
        RECT -74.285 56.275 -73.955 56.605 ;
        RECT -74.285 54.915 -73.955 55.245 ;
        RECT -74.285 53.555 -73.955 53.885 ;
        RECT -74.285 52.195 -73.955 52.525 ;
        RECT -74.285 50.835 -73.955 51.165 ;
        RECT -74.285 49.475 -73.955 49.805 ;
        RECT -74.285 48.115 -73.955 48.445 ;
        RECT -74.285 46.755 -73.955 47.085 ;
        RECT -74.285 45.395 -73.955 45.725 ;
        RECT -74.285 44.035 -73.955 44.365 ;
        RECT -74.285 42.675 -73.955 43.005 ;
        RECT -74.285 41.315 -73.955 41.645 ;
        RECT -74.285 39.955 -73.955 40.285 ;
        RECT -74.285 38.595 -73.955 38.925 ;
        RECT -74.285 37.235 -73.955 37.565 ;
        RECT -74.285 35.875 -73.955 36.205 ;
        RECT -74.285 34.515 -73.955 34.845 ;
        RECT -74.285 33.155 -73.955 33.485 ;
        RECT -74.285 31.795 -73.955 32.125 ;
        RECT -74.285 30.435 -73.955 30.765 ;
        RECT -74.285 29.075 -73.955 29.405 ;
        RECT -74.285 27.715 -73.955 28.045 ;
        RECT -74.285 26.355 -73.955 26.685 ;
        RECT -74.285 24.995 -73.955 25.325 ;
        RECT -74.285 23.635 -73.955 23.965 ;
        RECT -74.285 22.275 -73.955 22.605 ;
        RECT -74.285 20.915 -73.955 21.245 ;
        RECT -74.285 19.555 -73.955 19.885 ;
        RECT -74.285 18.195 -73.955 18.525 ;
        RECT -74.285 16.835 -73.955 17.165 ;
        RECT -74.285 15.475 -73.955 15.805 ;
        RECT -74.285 14.115 -73.955 14.445 ;
        RECT -74.285 12.755 -73.955 13.085 ;
        RECT -74.285 11.395 -73.955 11.725 ;
        RECT -74.285 10.035 -73.955 10.365 ;
        RECT -74.285 8.675 -73.955 9.005 ;
        RECT -74.285 7.315 -73.955 7.645 ;
        RECT -74.285 5.955 -73.955 6.285 ;
        RECT -74.285 4.595 -73.955 4.925 ;
        RECT -74.285 3.235 -73.955 3.565 ;
        RECT -74.285 1.875 -73.955 2.205 ;
        RECT -74.285 0.515 -73.955 0.845 ;
        RECT -74.285 -0.845 -73.955 -0.515 ;
        RECT -74.285 -2.205 -73.955 -1.875 ;
        RECT -74.285 -3.565 -73.955 -3.235 ;
        RECT -74.285 -4.925 -73.955 -4.595 ;
        RECT -74.285 -6.285 -73.955 -5.955 ;
        RECT -74.285 -7.645 -73.955 -7.315 ;
        RECT -74.285 -9.005 -73.955 -8.675 ;
        RECT -74.285 -10.365 -73.955 -10.035 ;
        RECT -74.285 -11.725 -73.955 -11.395 ;
        RECT -74.285 -13.085 -73.955 -12.755 ;
        RECT -74.285 -14.445 -73.955 -14.115 ;
        RECT -74.285 -15.805 -73.955 -15.475 ;
        RECT -74.285 -17.165 -73.955 -16.835 ;
        RECT -74.285 -18.525 -73.955 -18.195 ;
        RECT -74.285 -19.885 -73.955 -19.555 ;
        RECT -74.285 -21.245 -73.955 -20.915 ;
        RECT -74.285 -22.605 -73.955 -22.275 ;
        RECT -74.285 -23.965 -73.955 -23.635 ;
        RECT -74.285 -25.325 -73.955 -24.995 ;
        RECT -74.285 -26.685 -73.955 -26.355 ;
        RECT -74.285 -28.045 -73.955 -27.715 ;
        RECT -74.285 -29.405 -73.955 -29.075 ;
        RECT -74.285 -30.765 -73.955 -30.435 ;
        RECT -74.285 -32.125 -73.955 -31.795 ;
        RECT -74.285 -33.485 -73.955 -33.155 ;
        RECT -74.285 -34.845 -73.955 -34.515 ;
        RECT -74.285 -36.205 -73.955 -35.875 ;
        RECT -74.285 -37.565 -73.955 -37.235 ;
        RECT -74.285 -38.925 -73.955 -38.595 ;
        RECT -74.285 -40.285 -73.955 -39.955 ;
        RECT -74.285 -41.645 -73.955 -41.315 ;
        RECT -74.285 -43.005 -73.955 -42.675 ;
        RECT -74.285 -44.365 -73.955 -44.035 ;
        RECT -74.285 -45.725 -73.955 -45.395 ;
        RECT -74.285 -47.085 -73.955 -46.755 ;
        RECT -74.285 -48.445 -73.955 -48.115 ;
        RECT -74.285 -49.805 -73.955 -49.475 ;
        RECT -74.285 -51.165 -73.955 -50.835 ;
        RECT -74.285 -52.525 -73.955 -52.195 ;
        RECT -74.285 -53.885 -73.955 -53.555 ;
        RECT -74.285 -55.245 -73.955 -54.915 ;
        RECT -74.285 -56.605 -73.955 -56.275 ;
        RECT -74.285 -57.965 -73.955 -57.635 ;
        RECT -74.285 -59.325 -73.955 -58.995 ;
        RECT -74.285 -60.685 -73.955 -60.355 ;
        RECT -74.285 -62.045 -73.955 -61.715 ;
        RECT -74.285 -63.405 -73.955 -63.075 ;
        RECT -74.285 -64.765 -73.955 -64.435 ;
        RECT -74.285 -66.125 -73.955 -65.795 ;
        RECT -74.285 -67.485 -73.955 -67.155 ;
        RECT -74.285 -68.845 -73.955 -68.515 ;
        RECT -74.285 -70.205 -73.955 -69.875 ;
        RECT -74.285 -71.565 -73.955 -71.235 ;
        RECT -74.285 -72.925 -73.955 -72.595 ;
        RECT -74.285 -74.285 -73.955 -73.955 ;
        RECT -74.285 -75.645 -73.955 -75.315 ;
        RECT -74.285 -77.005 -73.955 -76.675 ;
        RECT -74.285 -78.365 -73.955 -78.035 ;
        RECT -74.285 -79.725 -73.955 -79.395 ;
        RECT -74.285 -81.085 -73.955 -80.755 ;
        RECT -74.285 -82.445 -73.955 -82.115 ;
        RECT -74.285 -83.805 -73.955 -83.475 ;
        RECT -74.285 -85.165 -73.955 -84.835 ;
        RECT -74.285 -86.525 -73.955 -86.195 ;
        RECT -74.285 -87.885 -73.955 -87.555 ;
        RECT -74.285 -89.245 -73.955 -88.915 ;
        RECT -74.285 -90.605 -73.955 -90.275 ;
        RECT -74.285 -91.965 -73.955 -91.635 ;
        RECT -74.285 -93.325 -73.955 -92.995 ;
        RECT -74.285 -94.685 -73.955 -94.355 ;
        RECT -74.285 -96.045 -73.955 -95.715 ;
        RECT -74.285 -97.405 -73.955 -97.075 ;
        RECT -74.285 -98.765 -73.955 -98.435 ;
        RECT -74.285 -100.125 -73.955 -99.795 ;
        RECT -74.285 -101.485 -73.955 -101.155 ;
        RECT -74.285 -102.845 -73.955 -102.515 ;
        RECT -74.285 -104.205 -73.955 -103.875 ;
        RECT -74.285 -105.565 -73.955 -105.235 ;
        RECT -74.285 -106.925 -73.955 -106.595 ;
        RECT -74.285 -108.285 -73.955 -107.955 ;
        RECT -74.285 -109.645 -73.955 -109.315 ;
        RECT -74.285 -111.005 -73.955 -110.675 ;
        RECT -74.285 -112.365 -73.955 -112.035 ;
        RECT -74.285 -113.725 -73.955 -113.395 ;
        RECT -74.285 -115.085 -73.955 -114.755 ;
        RECT -74.285 -116.445 -73.955 -116.115 ;
        RECT -74.285 -117.805 -73.955 -117.475 ;
        RECT -74.285 -119.165 -73.955 -118.835 ;
        RECT -74.285 -120.525 -73.955 -120.195 ;
        RECT -74.285 -121.885 -73.955 -121.555 ;
        RECT -74.285 -123.245 -73.955 -122.915 ;
        RECT -74.285 -124.605 -73.955 -124.275 ;
        RECT -74.285 -125.965 -73.955 -125.635 ;
        RECT -74.285 -127.325 -73.955 -126.995 ;
        RECT -74.285 -128.685 -73.955 -128.355 ;
        RECT -74.285 -130.045 -73.955 -129.715 ;
        RECT -74.285 -131.405 -73.955 -131.075 ;
        RECT -74.285 -132.765 -73.955 -132.435 ;
        RECT -74.285 -134.125 -73.955 -133.795 ;
        RECT -74.285 -135.485 -73.955 -135.155 ;
        RECT -74.285 -136.845 -73.955 -136.515 ;
        RECT -74.285 -138.205 -73.955 -137.875 ;
        RECT -74.285 -139.565 -73.955 -139.235 ;
        RECT -74.285 -140.925 -73.955 -140.595 ;
        RECT -74.285 -142.285 -73.955 -141.955 ;
        RECT -74.285 -143.645 -73.955 -143.315 ;
        RECT -74.285 -145.005 -73.955 -144.675 ;
        RECT -74.285 -146.365 -73.955 -146.035 ;
        RECT -74.285 -147.725 -73.955 -147.395 ;
        RECT -74.285 -149.085 -73.955 -148.755 ;
        RECT -74.285 -150.445 -73.955 -150.115 ;
        RECT -74.285 -151.805 -73.955 -151.475 ;
        RECT -74.285 -153.165 -73.955 -152.835 ;
        RECT -74.285 -154.525 -73.955 -154.195 ;
        RECT -74.285 -155.885 -73.955 -155.555 ;
        RECT -74.285 -157.245 -73.955 -156.915 ;
        RECT -74.285 -158.605 -73.955 -158.275 ;
        RECT -74.285 -159.965 -73.955 -159.635 ;
        RECT -74.285 -161.325 -73.955 -160.995 ;
        RECT -74.285 -162.685 -73.955 -162.355 ;
        RECT -74.285 -164.045 -73.955 -163.715 ;
        RECT -74.285 -165.405 -73.955 -165.075 ;
        RECT -74.285 -166.765 -73.955 -166.435 ;
        RECT -74.285 -168.125 -73.955 -167.795 ;
        RECT -74.285 -169.485 -73.955 -169.155 ;
        RECT -74.285 -170.845 -73.955 -170.515 ;
        RECT -74.285 -172.205 -73.955 -171.875 ;
        RECT -74.285 -173.565 -73.955 -173.235 ;
        RECT -74.285 -174.925 -73.955 -174.595 ;
        RECT -74.285 -176.285 -73.955 -175.955 ;
        RECT -74.285 -177.645 -73.955 -177.315 ;
        RECT -74.285 -183.29 -73.955 -182.16 ;
        RECT -74.28 -183.405 -73.96 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -72.925 244.04 -72.595 245.17 ;
        RECT -72.925 239.875 -72.595 240.205 ;
        RECT -72.925 238.515 -72.595 238.845 ;
        RECT -72.925 237.155 -72.595 237.485 ;
        RECT -72.925 235.795 -72.595 236.125 ;
        RECT -72.925 234.435 -72.595 234.765 ;
        RECT -72.925 233.075 -72.595 233.405 ;
        RECT -72.925 231.715 -72.595 232.045 ;
        RECT -72.925 230.355 -72.595 230.685 ;
        RECT -72.925 228.995 -72.595 229.325 ;
        RECT -72.925 227.635 -72.595 227.965 ;
        RECT -72.925 226.275 -72.595 226.605 ;
        RECT -72.925 224.915 -72.595 225.245 ;
        RECT -72.925 223.555 -72.595 223.885 ;
        RECT -72.925 222.195 -72.595 222.525 ;
        RECT -72.925 220.835 -72.595 221.165 ;
        RECT -72.925 219.475 -72.595 219.805 ;
        RECT -72.925 218.115 -72.595 218.445 ;
        RECT -72.925 216.755 -72.595 217.085 ;
        RECT -72.925 215.395 -72.595 215.725 ;
        RECT -72.925 214.035 -72.595 214.365 ;
        RECT -72.925 212.675 -72.595 213.005 ;
        RECT -72.925 211.315 -72.595 211.645 ;
        RECT -72.925 209.955 -72.595 210.285 ;
        RECT -72.925 208.595 -72.595 208.925 ;
        RECT -72.925 207.235 -72.595 207.565 ;
        RECT -72.925 205.875 -72.595 206.205 ;
        RECT -72.925 204.515 -72.595 204.845 ;
        RECT -72.925 203.155 -72.595 203.485 ;
        RECT -72.925 201.795 -72.595 202.125 ;
        RECT -72.925 200.435 -72.595 200.765 ;
        RECT -72.925 199.075 -72.595 199.405 ;
        RECT -72.925 197.715 -72.595 198.045 ;
        RECT -72.925 196.355 -72.595 196.685 ;
        RECT -72.925 194.995 -72.595 195.325 ;
        RECT -72.925 193.635 -72.595 193.965 ;
        RECT -72.925 192.275 -72.595 192.605 ;
        RECT -72.925 190.915 -72.595 191.245 ;
        RECT -72.925 189.555 -72.595 189.885 ;
        RECT -72.925 188.195 -72.595 188.525 ;
        RECT -72.925 186.835 -72.595 187.165 ;
        RECT -72.925 185.475 -72.595 185.805 ;
        RECT -72.925 184.115 -72.595 184.445 ;
        RECT -72.925 182.755 -72.595 183.085 ;
        RECT -72.925 181.395 -72.595 181.725 ;
        RECT -72.925 180.035 -72.595 180.365 ;
        RECT -72.925 178.675 -72.595 179.005 ;
        RECT -72.925 177.315 -72.595 177.645 ;
        RECT -72.925 175.955 -72.595 176.285 ;
        RECT -72.925 174.595 -72.595 174.925 ;
        RECT -72.925 173.235 -72.595 173.565 ;
        RECT -72.925 171.875 -72.595 172.205 ;
        RECT -72.925 170.515 -72.595 170.845 ;
        RECT -72.925 169.155 -72.595 169.485 ;
        RECT -72.925 167.795 -72.595 168.125 ;
        RECT -72.925 166.435 -72.595 166.765 ;
        RECT -72.925 165.075 -72.595 165.405 ;
        RECT -72.925 163.715 -72.595 164.045 ;
        RECT -72.925 162.355 -72.595 162.685 ;
        RECT -72.925 160.995 -72.595 161.325 ;
        RECT -72.925 159.635 -72.595 159.965 ;
        RECT -72.925 158.275 -72.595 158.605 ;
        RECT -72.925 156.915 -72.595 157.245 ;
        RECT -72.925 155.555 -72.595 155.885 ;
        RECT -72.925 154.195 -72.595 154.525 ;
        RECT -72.925 152.835 -72.595 153.165 ;
        RECT -72.925 151.475 -72.595 151.805 ;
        RECT -72.925 150.115 -72.595 150.445 ;
        RECT -72.925 148.755 -72.595 149.085 ;
        RECT -72.925 147.395 -72.595 147.725 ;
        RECT -72.925 146.035 -72.595 146.365 ;
        RECT -72.925 144.675 -72.595 145.005 ;
        RECT -72.925 143.315 -72.595 143.645 ;
        RECT -72.925 141.955 -72.595 142.285 ;
        RECT -72.925 140.595 -72.595 140.925 ;
        RECT -72.925 139.235 -72.595 139.565 ;
        RECT -72.925 137.875 -72.595 138.205 ;
        RECT -72.925 136.515 -72.595 136.845 ;
        RECT -72.925 135.155 -72.595 135.485 ;
        RECT -72.925 133.795 -72.595 134.125 ;
        RECT -72.925 132.435 -72.595 132.765 ;
        RECT -72.925 131.075 -72.595 131.405 ;
        RECT -72.925 129.715 -72.595 130.045 ;
        RECT -72.925 128.355 -72.595 128.685 ;
        RECT -72.925 126.995 -72.595 127.325 ;
        RECT -72.925 125.635 -72.595 125.965 ;
        RECT -72.925 124.275 -72.595 124.605 ;
        RECT -72.925 122.915 -72.595 123.245 ;
        RECT -72.925 121.555 -72.595 121.885 ;
        RECT -72.925 120.195 -72.595 120.525 ;
        RECT -72.925 118.835 -72.595 119.165 ;
        RECT -72.925 117.475 -72.595 117.805 ;
        RECT -72.925 116.115 -72.595 116.445 ;
        RECT -72.925 114.755 -72.595 115.085 ;
        RECT -72.925 113.395 -72.595 113.725 ;
        RECT -72.925 112.035 -72.595 112.365 ;
        RECT -72.925 110.675 -72.595 111.005 ;
        RECT -72.925 109.315 -72.595 109.645 ;
        RECT -72.925 107.955 -72.595 108.285 ;
        RECT -72.925 106.595 -72.595 106.925 ;
        RECT -72.925 105.235 -72.595 105.565 ;
        RECT -72.925 103.875 -72.595 104.205 ;
        RECT -72.925 102.515 -72.595 102.845 ;
        RECT -72.925 101.155 -72.595 101.485 ;
        RECT -72.925 99.795 -72.595 100.125 ;
        RECT -72.925 98.435 -72.595 98.765 ;
        RECT -72.925 97.075 -72.595 97.405 ;
        RECT -72.925 95.715 -72.595 96.045 ;
        RECT -72.925 94.355 -72.595 94.685 ;
        RECT -72.925 92.995 -72.595 93.325 ;
        RECT -72.925 91.635 -72.595 91.965 ;
        RECT -72.925 90.275 -72.595 90.605 ;
        RECT -72.925 88.915 -72.595 89.245 ;
        RECT -72.925 87.555 -72.595 87.885 ;
        RECT -72.925 86.195 -72.595 86.525 ;
        RECT -72.925 84.835 -72.595 85.165 ;
        RECT -72.925 83.475 -72.595 83.805 ;
        RECT -72.925 82.115 -72.595 82.445 ;
        RECT -72.925 80.755 -72.595 81.085 ;
        RECT -72.925 79.395 -72.595 79.725 ;
        RECT -72.925 78.035 -72.595 78.365 ;
        RECT -72.925 76.675 -72.595 77.005 ;
        RECT -72.925 75.315 -72.595 75.645 ;
        RECT -72.925 73.955 -72.595 74.285 ;
        RECT -72.925 72.595 -72.595 72.925 ;
        RECT -72.925 71.235 -72.595 71.565 ;
        RECT -72.925 69.875 -72.595 70.205 ;
        RECT -72.925 68.515 -72.595 68.845 ;
        RECT -72.925 67.155 -72.595 67.485 ;
        RECT -72.925 65.795 -72.595 66.125 ;
        RECT -72.925 64.435 -72.595 64.765 ;
        RECT -72.925 63.075 -72.595 63.405 ;
        RECT -72.925 61.715 -72.595 62.045 ;
        RECT -72.925 60.355 -72.595 60.685 ;
        RECT -72.925 58.995 -72.595 59.325 ;
        RECT -72.925 57.635 -72.595 57.965 ;
        RECT -72.925 56.275 -72.595 56.605 ;
        RECT -72.925 54.915 -72.595 55.245 ;
        RECT -72.925 53.555 -72.595 53.885 ;
        RECT -72.925 52.195 -72.595 52.525 ;
        RECT -72.925 50.835 -72.595 51.165 ;
        RECT -72.925 49.475 -72.595 49.805 ;
        RECT -72.925 48.115 -72.595 48.445 ;
        RECT -72.925 46.755 -72.595 47.085 ;
        RECT -72.925 45.395 -72.595 45.725 ;
        RECT -72.925 44.035 -72.595 44.365 ;
        RECT -72.925 42.675 -72.595 43.005 ;
        RECT -72.925 41.315 -72.595 41.645 ;
        RECT -72.925 39.955 -72.595 40.285 ;
        RECT -72.925 38.595 -72.595 38.925 ;
        RECT -72.925 37.235 -72.595 37.565 ;
        RECT -72.925 35.875 -72.595 36.205 ;
        RECT -72.925 34.515 -72.595 34.845 ;
        RECT -72.925 33.155 -72.595 33.485 ;
        RECT -72.925 31.795 -72.595 32.125 ;
        RECT -72.925 30.435 -72.595 30.765 ;
        RECT -72.925 29.075 -72.595 29.405 ;
        RECT -72.925 27.715 -72.595 28.045 ;
        RECT -72.925 26.355 -72.595 26.685 ;
        RECT -72.925 24.995 -72.595 25.325 ;
        RECT -72.925 23.635 -72.595 23.965 ;
        RECT -72.925 22.275 -72.595 22.605 ;
        RECT -72.925 20.915 -72.595 21.245 ;
        RECT -72.925 19.555 -72.595 19.885 ;
        RECT -72.925 18.195 -72.595 18.525 ;
        RECT -72.925 16.835 -72.595 17.165 ;
        RECT -72.925 15.475 -72.595 15.805 ;
        RECT -72.925 14.115 -72.595 14.445 ;
        RECT -72.925 12.755 -72.595 13.085 ;
        RECT -72.925 11.395 -72.595 11.725 ;
        RECT -72.925 10.035 -72.595 10.365 ;
        RECT -72.925 8.675 -72.595 9.005 ;
        RECT -72.925 7.315 -72.595 7.645 ;
        RECT -72.925 5.955 -72.595 6.285 ;
        RECT -72.925 4.595 -72.595 4.925 ;
        RECT -72.925 3.235 -72.595 3.565 ;
        RECT -72.925 1.875 -72.595 2.205 ;
        RECT -72.925 0.515 -72.595 0.845 ;
        RECT -72.925 -0.845 -72.595 -0.515 ;
        RECT -72.925 -2.205 -72.595 -1.875 ;
        RECT -72.925 -3.565 -72.595 -3.235 ;
        RECT -72.925 -4.925 -72.595 -4.595 ;
        RECT -72.925 -6.285 -72.595 -5.955 ;
        RECT -72.925 -7.645 -72.595 -7.315 ;
        RECT -72.925 -9.005 -72.595 -8.675 ;
        RECT -72.925 -10.365 -72.595 -10.035 ;
        RECT -72.925 -11.725 -72.595 -11.395 ;
        RECT -72.925 -13.085 -72.595 -12.755 ;
        RECT -72.925 -14.445 -72.595 -14.115 ;
        RECT -72.925 -15.805 -72.595 -15.475 ;
        RECT -72.925 -17.165 -72.595 -16.835 ;
        RECT -72.925 -18.525 -72.595 -18.195 ;
        RECT -72.925 -19.885 -72.595 -19.555 ;
        RECT -72.925 -21.245 -72.595 -20.915 ;
        RECT -72.925 -22.605 -72.595 -22.275 ;
        RECT -72.925 -23.965 -72.595 -23.635 ;
        RECT -72.925 -25.325 -72.595 -24.995 ;
        RECT -72.925 -26.685 -72.595 -26.355 ;
        RECT -72.925 -28.045 -72.595 -27.715 ;
        RECT -72.925 -29.405 -72.595 -29.075 ;
        RECT -72.925 -30.765 -72.595 -30.435 ;
        RECT -72.925 -32.125 -72.595 -31.795 ;
        RECT -72.925 -33.485 -72.595 -33.155 ;
        RECT -72.925 -34.845 -72.595 -34.515 ;
        RECT -72.925 -36.205 -72.595 -35.875 ;
        RECT -72.925 -37.565 -72.595 -37.235 ;
        RECT -72.925 -38.925 -72.595 -38.595 ;
        RECT -72.925 -40.285 -72.595 -39.955 ;
        RECT -72.925 -41.645 -72.595 -41.315 ;
        RECT -72.925 -43.005 -72.595 -42.675 ;
        RECT -72.925 -44.365 -72.595 -44.035 ;
        RECT -72.925 -45.725 -72.595 -45.395 ;
        RECT -72.925 -47.085 -72.595 -46.755 ;
        RECT -72.925 -48.445 -72.595 -48.115 ;
        RECT -72.925 -49.805 -72.595 -49.475 ;
        RECT -72.925 -51.165 -72.595 -50.835 ;
        RECT -72.925 -52.525 -72.595 -52.195 ;
        RECT -72.925 -53.885 -72.595 -53.555 ;
        RECT -72.925 -55.245 -72.595 -54.915 ;
        RECT -72.925 -56.605 -72.595 -56.275 ;
        RECT -72.925 -57.965 -72.595 -57.635 ;
        RECT -72.925 -59.325 -72.595 -58.995 ;
        RECT -72.925 -60.685 -72.595 -60.355 ;
        RECT -72.925 -62.045 -72.595 -61.715 ;
        RECT -72.925 -63.405 -72.595 -63.075 ;
        RECT -72.925 -64.765 -72.595 -64.435 ;
        RECT -72.925 -66.125 -72.595 -65.795 ;
        RECT -72.925 -67.485 -72.595 -67.155 ;
        RECT -72.925 -68.845 -72.595 -68.515 ;
        RECT -72.925 -70.205 -72.595 -69.875 ;
        RECT -72.925 -71.565 -72.595 -71.235 ;
        RECT -72.925 -72.925 -72.595 -72.595 ;
        RECT -72.925 -74.285 -72.595 -73.955 ;
        RECT -72.925 -75.645 -72.595 -75.315 ;
        RECT -72.925 -77.005 -72.595 -76.675 ;
        RECT -72.925 -78.365 -72.595 -78.035 ;
        RECT -72.925 -79.725 -72.595 -79.395 ;
        RECT -72.925 -81.085 -72.595 -80.755 ;
        RECT -72.925 -82.445 -72.595 -82.115 ;
        RECT -72.925 -83.805 -72.595 -83.475 ;
        RECT -72.925 -85.165 -72.595 -84.835 ;
        RECT -72.925 -86.525 -72.595 -86.195 ;
        RECT -72.925 -87.885 -72.595 -87.555 ;
        RECT -72.925 -89.245 -72.595 -88.915 ;
        RECT -72.925 -90.605 -72.595 -90.275 ;
        RECT -72.925 -91.965 -72.595 -91.635 ;
        RECT -72.925 -93.325 -72.595 -92.995 ;
        RECT -72.925 -94.685 -72.595 -94.355 ;
        RECT -72.925 -96.045 -72.595 -95.715 ;
        RECT -72.925 -97.405 -72.595 -97.075 ;
        RECT -72.925 -98.765 -72.595 -98.435 ;
        RECT -72.925 -100.125 -72.595 -99.795 ;
        RECT -72.925 -101.485 -72.595 -101.155 ;
        RECT -72.925 -102.845 -72.595 -102.515 ;
        RECT -72.925 -104.205 -72.595 -103.875 ;
        RECT -72.925 -105.565 -72.595 -105.235 ;
        RECT -72.925 -106.925 -72.595 -106.595 ;
        RECT -72.925 -108.285 -72.595 -107.955 ;
        RECT -72.925 -109.645 -72.595 -109.315 ;
        RECT -72.925 -111.005 -72.595 -110.675 ;
        RECT -72.925 -112.365 -72.595 -112.035 ;
        RECT -72.925 -113.725 -72.595 -113.395 ;
        RECT -72.925 -115.085 -72.595 -114.755 ;
        RECT -72.925 -116.445 -72.595 -116.115 ;
        RECT -72.925 -117.805 -72.595 -117.475 ;
        RECT -72.925 -119.165 -72.595 -118.835 ;
        RECT -72.925 -120.525 -72.595 -120.195 ;
        RECT -72.925 -121.885 -72.595 -121.555 ;
        RECT -72.925 -123.245 -72.595 -122.915 ;
        RECT -72.925 -124.605 -72.595 -124.275 ;
        RECT -72.925 -125.965 -72.595 -125.635 ;
        RECT -72.925 -127.325 -72.595 -126.995 ;
        RECT -72.925 -128.685 -72.595 -128.355 ;
        RECT -72.925 -130.045 -72.595 -129.715 ;
        RECT -72.925 -131.405 -72.595 -131.075 ;
        RECT -72.925 -132.765 -72.595 -132.435 ;
        RECT -72.925 -134.125 -72.595 -133.795 ;
        RECT -72.925 -135.485 -72.595 -135.155 ;
        RECT -72.925 -136.845 -72.595 -136.515 ;
        RECT -72.925 -138.205 -72.595 -137.875 ;
        RECT -72.925 -139.565 -72.595 -139.235 ;
        RECT -72.925 -140.925 -72.595 -140.595 ;
        RECT -72.925 -142.285 -72.595 -141.955 ;
        RECT -72.925 -143.645 -72.595 -143.315 ;
        RECT -72.925 -145.005 -72.595 -144.675 ;
        RECT -72.925 -146.365 -72.595 -146.035 ;
        RECT -72.925 -147.725 -72.595 -147.395 ;
        RECT -72.925 -149.085 -72.595 -148.755 ;
        RECT -72.925 -150.445 -72.595 -150.115 ;
        RECT -72.925 -151.805 -72.595 -151.475 ;
        RECT -72.925 -153.165 -72.595 -152.835 ;
        RECT -72.925 -154.525 -72.595 -154.195 ;
        RECT -72.925 -155.885 -72.595 -155.555 ;
        RECT -72.925 -157.245 -72.595 -156.915 ;
        RECT -72.925 -158.605 -72.595 -158.275 ;
        RECT -72.925 -159.965 -72.595 -159.635 ;
        RECT -72.925 -161.325 -72.595 -160.995 ;
        RECT -72.925 -162.685 -72.595 -162.355 ;
        RECT -72.925 -164.045 -72.595 -163.715 ;
        RECT -72.925 -165.405 -72.595 -165.075 ;
        RECT -72.925 -166.765 -72.595 -166.435 ;
        RECT -72.925 -168.125 -72.595 -167.795 ;
        RECT -72.925 -169.485 -72.595 -169.155 ;
        RECT -72.925 -170.845 -72.595 -170.515 ;
        RECT -72.925 -172.205 -72.595 -171.875 ;
        RECT -72.925 -173.565 -72.595 -173.235 ;
        RECT -72.925 -174.925 -72.595 -174.595 ;
        RECT -72.925 -176.285 -72.595 -175.955 ;
        RECT -72.925 -177.645 -72.595 -177.315 ;
        RECT -72.925 -183.29 -72.595 -182.16 ;
        RECT -72.92 -183.405 -72.6 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -71.565 -18.525 -71.235 -18.195 ;
        RECT -71.565 -19.885 -71.235 -19.555 ;
        RECT -71.565 -21.245 -71.235 -20.915 ;
        RECT -71.565 -22.605 -71.235 -22.275 ;
        RECT -71.565 -23.965 -71.235 -23.635 ;
        RECT -71.565 -25.325 -71.235 -24.995 ;
        RECT -71.565 -26.685 -71.235 -26.355 ;
        RECT -71.565 -28.045 -71.235 -27.715 ;
        RECT -71.565 -29.405 -71.235 -29.075 ;
        RECT -71.565 -30.765 -71.235 -30.435 ;
        RECT -71.565 -32.125 -71.235 -31.795 ;
        RECT -71.565 -33.485 -71.235 -33.155 ;
        RECT -71.565 -34.845 -71.235 -34.515 ;
        RECT -71.565 -36.205 -71.235 -35.875 ;
        RECT -71.565 -37.565 -71.235 -37.235 ;
        RECT -71.565 -38.925 -71.235 -38.595 ;
        RECT -71.565 -40.285 -71.235 -39.955 ;
        RECT -71.565 -41.645 -71.235 -41.315 ;
        RECT -71.565 -43.005 -71.235 -42.675 ;
        RECT -71.565 -44.365 -71.235 -44.035 ;
        RECT -71.565 -45.725 -71.235 -45.395 ;
        RECT -71.565 -47.085 -71.235 -46.755 ;
        RECT -71.565 -48.445 -71.235 -48.115 ;
        RECT -71.565 -49.805 -71.235 -49.475 ;
        RECT -71.565 -51.165 -71.235 -50.835 ;
        RECT -71.565 -52.525 -71.235 -52.195 ;
        RECT -71.565 -53.885 -71.235 -53.555 ;
        RECT -71.565 -55.245 -71.235 -54.915 ;
        RECT -71.565 -56.605 -71.235 -56.275 ;
        RECT -71.565 -57.965 -71.235 -57.635 ;
        RECT -71.565 -59.325 -71.235 -58.995 ;
        RECT -71.565 -60.685 -71.235 -60.355 ;
        RECT -71.565 -62.045 -71.235 -61.715 ;
        RECT -71.565 -63.405 -71.235 -63.075 ;
        RECT -71.565 -64.765 -71.235 -64.435 ;
        RECT -71.565 -66.125 -71.235 -65.795 ;
        RECT -71.565 -67.485 -71.235 -67.155 ;
        RECT -71.565 -68.845 -71.235 -68.515 ;
        RECT -71.565 -70.205 -71.235 -69.875 ;
        RECT -71.565 -71.565 -71.235 -71.235 ;
        RECT -71.565 -72.925 -71.235 -72.595 ;
        RECT -71.565 -74.285 -71.235 -73.955 ;
        RECT -71.565 -75.645 -71.235 -75.315 ;
        RECT -71.565 -77.005 -71.235 -76.675 ;
        RECT -71.565 -78.365 -71.235 -78.035 ;
        RECT -71.565 -79.725 -71.235 -79.395 ;
        RECT -71.565 -81.085 -71.235 -80.755 ;
        RECT -71.565 -82.445 -71.235 -82.115 ;
        RECT -71.565 -83.805 -71.235 -83.475 ;
        RECT -71.565 -85.165 -71.235 -84.835 ;
        RECT -71.565 -86.525 -71.235 -86.195 ;
        RECT -71.565 -87.885 -71.235 -87.555 ;
        RECT -71.565 -89.245 -71.235 -88.915 ;
        RECT -71.565 -90.605 -71.235 -90.275 ;
        RECT -71.565 -91.965 -71.235 -91.635 ;
        RECT -71.565 -93.325 -71.235 -92.995 ;
        RECT -71.565 -94.685 -71.235 -94.355 ;
        RECT -71.565 -96.045 -71.235 -95.715 ;
        RECT -71.565 -97.405 -71.235 -97.075 ;
        RECT -71.565 -98.765 -71.235 -98.435 ;
        RECT -71.565 -100.125 -71.235 -99.795 ;
        RECT -71.565 -101.485 -71.235 -101.155 ;
        RECT -71.565 -102.845 -71.235 -102.515 ;
        RECT -71.565 -104.205 -71.235 -103.875 ;
        RECT -71.565 -105.565 -71.235 -105.235 ;
        RECT -71.565 -106.925 -71.235 -106.595 ;
        RECT -71.565 -108.285 -71.235 -107.955 ;
        RECT -71.565 -109.645 -71.235 -109.315 ;
        RECT -71.565 -111.005 -71.235 -110.675 ;
        RECT -71.565 -112.365 -71.235 -112.035 ;
        RECT -71.565 -113.725 -71.235 -113.395 ;
        RECT -71.565 -115.085 -71.235 -114.755 ;
        RECT -71.565 -116.445 -71.235 -116.115 ;
        RECT -71.565 -117.805 -71.235 -117.475 ;
        RECT -71.565 -119.165 -71.235 -118.835 ;
        RECT -71.565 -120.525 -71.235 -120.195 ;
        RECT -71.565 -121.885 -71.235 -121.555 ;
        RECT -71.565 -123.245 -71.235 -122.915 ;
        RECT -71.565 -124.605 -71.235 -124.275 ;
        RECT -71.565 -125.965 -71.235 -125.635 ;
        RECT -71.565 -127.325 -71.235 -126.995 ;
        RECT -71.565 -128.685 -71.235 -128.355 ;
        RECT -71.565 -130.045 -71.235 -129.715 ;
        RECT -71.565 -131.405 -71.235 -131.075 ;
        RECT -71.565 -132.765 -71.235 -132.435 ;
        RECT -71.565 -134.125 -71.235 -133.795 ;
        RECT -71.565 -135.485 -71.235 -135.155 ;
        RECT -71.565 -136.845 -71.235 -136.515 ;
        RECT -71.565 -138.205 -71.235 -137.875 ;
        RECT -71.565 -139.565 -71.235 -139.235 ;
        RECT -71.565 -140.925 -71.235 -140.595 ;
        RECT -71.565 -142.285 -71.235 -141.955 ;
        RECT -71.565 -143.645 -71.235 -143.315 ;
        RECT -71.565 -145.005 -71.235 -144.675 ;
        RECT -71.565 -146.365 -71.235 -146.035 ;
        RECT -71.565 -147.725 -71.235 -147.395 ;
        RECT -71.565 -149.085 -71.235 -148.755 ;
        RECT -71.565 -150.445 -71.235 -150.115 ;
        RECT -71.565 -151.805 -71.235 -151.475 ;
        RECT -71.565 -153.165 -71.235 -152.835 ;
        RECT -71.565 -154.525 -71.235 -154.195 ;
        RECT -71.565 -155.885 -71.235 -155.555 ;
        RECT -71.565 -157.245 -71.235 -156.915 ;
        RECT -71.565 -158.605 -71.235 -158.275 ;
        RECT -71.565 -159.965 -71.235 -159.635 ;
        RECT -71.565 -161.325 -71.235 -160.995 ;
        RECT -71.565 -162.685 -71.235 -162.355 ;
        RECT -71.565 -164.045 -71.235 -163.715 ;
        RECT -71.565 -165.405 -71.235 -165.075 ;
        RECT -71.565 -166.765 -71.235 -166.435 ;
        RECT -71.565 -168.655 -71.235 -168.325 ;
        RECT -71.565 -169.485 -71.235 -169.155 ;
        RECT -71.565 -170.845 -71.235 -170.515 ;
        RECT -71.565 -172.205 -71.235 -171.875 ;
        RECT -71.565 -173.565 -71.235 -173.235 ;
        RECT -71.565 -174.925 -71.235 -174.595 ;
        RECT -71.565 -177.645 -71.235 -177.315 ;
        RECT -71.565 -183.29 -71.235 -182.16 ;
        RECT -71.56 -183.405 -71.24 245.285 ;
        RECT -71.565 244.04 -71.235 245.17 ;
        RECT -71.565 239.875 -71.235 240.205 ;
        RECT -71.565 238.515 -71.235 238.845 ;
        RECT -71.565 237.155 -71.235 237.485 ;
        RECT -71.565 235.795 -71.235 236.125 ;
        RECT -71.565 234.435 -71.235 234.765 ;
        RECT -71.565 233.075 -71.235 233.405 ;
        RECT -71.565 231.715 -71.235 232.045 ;
        RECT -71.565 230.355 -71.235 230.685 ;
        RECT -71.565 228.995 -71.235 229.325 ;
        RECT -71.565 227.635 -71.235 227.965 ;
        RECT -71.565 226.275 -71.235 226.605 ;
        RECT -71.565 224.915 -71.235 225.245 ;
        RECT -71.565 223.555 -71.235 223.885 ;
        RECT -71.565 222.195 -71.235 222.525 ;
        RECT -71.565 220.835 -71.235 221.165 ;
        RECT -71.565 219.475 -71.235 219.805 ;
        RECT -71.565 218.115 -71.235 218.445 ;
        RECT -71.565 216.755 -71.235 217.085 ;
        RECT -71.565 215.395 -71.235 215.725 ;
        RECT -71.565 214.035 -71.235 214.365 ;
        RECT -71.565 212.675 -71.235 213.005 ;
        RECT -71.565 211.315 -71.235 211.645 ;
        RECT -71.565 209.955 -71.235 210.285 ;
        RECT -71.565 208.595 -71.235 208.925 ;
        RECT -71.565 207.235 -71.235 207.565 ;
        RECT -71.565 205.875 -71.235 206.205 ;
        RECT -71.565 204.515 -71.235 204.845 ;
        RECT -71.565 203.155 -71.235 203.485 ;
        RECT -71.565 201.795 -71.235 202.125 ;
        RECT -71.565 200.435 -71.235 200.765 ;
        RECT -71.565 199.075 -71.235 199.405 ;
        RECT -71.565 197.715 -71.235 198.045 ;
        RECT -71.565 196.355 -71.235 196.685 ;
        RECT -71.565 194.995 -71.235 195.325 ;
        RECT -71.565 193.635 -71.235 193.965 ;
        RECT -71.565 192.275 -71.235 192.605 ;
        RECT -71.565 190.915 -71.235 191.245 ;
        RECT -71.565 189.555 -71.235 189.885 ;
        RECT -71.565 188.195 -71.235 188.525 ;
        RECT -71.565 186.835 -71.235 187.165 ;
        RECT -71.565 185.475 -71.235 185.805 ;
        RECT -71.565 184.115 -71.235 184.445 ;
        RECT -71.565 182.755 -71.235 183.085 ;
        RECT -71.565 181.395 -71.235 181.725 ;
        RECT -71.565 180.035 -71.235 180.365 ;
        RECT -71.565 178.675 -71.235 179.005 ;
        RECT -71.565 177.315 -71.235 177.645 ;
        RECT -71.565 175.955 -71.235 176.285 ;
        RECT -71.565 174.595 -71.235 174.925 ;
        RECT -71.565 173.235 -71.235 173.565 ;
        RECT -71.565 171.875 -71.235 172.205 ;
        RECT -71.565 170.515 -71.235 170.845 ;
        RECT -71.565 169.155 -71.235 169.485 ;
        RECT -71.565 167.795 -71.235 168.125 ;
        RECT -71.565 166.435 -71.235 166.765 ;
        RECT -71.565 165.075 -71.235 165.405 ;
        RECT -71.565 163.715 -71.235 164.045 ;
        RECT -71.565 162.355 -71.235 162.685 ;
        RECT -71.565 160.995 -71.235 161.325 ;
        RECT -71.565 159.635 -71.235 159.965 ;
        RECT -71.565 158.275 -71.235 158.605 ;
        RECT -71.565 156.915 -71.235 157.245 ;
        RECT -71.565 155.555 -71.235 155.885 ;
        RECT -71.565 154.195 -71.235 154.525 ;
        RECT -71.565 152.835 -71.235 153.165 ;
        RECT -71.565 151.475 -71.235 151.805 ;
        RECT -71.565 150.115 -71.235 150.445 ;
        RECT -71.565 148.755 -71.235 149.085 ;
        RECT -71.565 147.395 -71.235 147.725 ;
        RECT -71.565 146.035 -71.235 146.365 ;
        RECT -71.565 144.675 -71.235 145.005 ;
        RECT -71.565 143.315 -71.235 143.645 ;
        RECT -71.565 141.955 -71.235 142.285 ;
        RECT -71.565 140.595 -71.235 140.925 ;
        RECT -71.565 139.235 -71.235 139.565 ;
        RECT -71.565 137.875 -71.235 138.205 ;
        RECT -71.565 136.515 -71.235 136.845 ;
        RECT -71.565 135.155 -71.235 135.485 ;
        RECT -71.565 133.795 -71.235 134.125 ;
        RECT -71.565 132.435 -71.235 132.765 ;
        RECT -71.565 131.075 -71.235 131.405 ;
        RECT -71.565 129.715 -71.235 130.045 ;
        RECT -71.565 128.355 -71.235 128.685 ;
        RECT -71.565 126.995 -71.235 127.325 ;
        RECT -71.565 125.635 -71.235 125.965 ;
        RECT -71.565 124.275 -71.235 124.605 ;
        RECT -71.565 122.915 -71.235 123.245 ;
        RECT -71.565 121.555 -71.235 121.885 ;
        RECT -71.565 120.195 -71.235 120.525 ;
        RECT -71.565 118.835 -71.235 119.165 ;
        RECT -71.565 117.475 -71.235 117.805 ;
        RECT -71.565 116.115 -71.235 116.445 ;
        RECT -71.565 114.755 -71.235 115.085 ;
        RECT -71.565 113.395 -71.235 113.725 ;
        RECT -71.565 112.035 -71.235 112.365 ;
        RECT -71.565 110.675 -71.235 111.005 ;
        RECT -71.565 109.315 -71.235 109.645 ;
        RECT -71.565 107.955 -71.235 108.285 ;
        RECT -71.565 106.595 -71.235 106.925 ;
        RECT -71.565 105.235 -71.235 105.565 ;
        RECT -71.565 103.875 -71.235 104.205 ;
        RECT -71.565 102.515 -71.235 102.845 ;
        RECT -71.565 101.155 -71.235 101.485 ;
        RECT -71.565 99.795 -71.235 100.125 ;
        RECT -71.565 98.435 -71.235 98.765 ;
        RECT -71.565 97.075 -71.235 97.405 ;
        RECT -71.565 95.715 -71.235 96.045 ;
        RECT -71.565 94.355 -71.235 94.685 ;
        RECT -71.565 92.995 -71.235 93.325 ;
        RECT -71.565 91.635 -71.235 91.965 ;
        RECT -71.565 90.275 -71.235 90.605 ;
        RECT -71.565 88.915 -71.235 89.245 ;
        RECT -71.565 87.555 -71.235 87.885 ;
        RECT -71.565 86.195 -71.235 86.525 ;
        RECT -71.565 84.835 -71.235 85.165 ;
        RECT -71.565 83.475 -71.235 83.805 ;
        RECT -71.565 82.115 -71.235 82.445 ;
        RECT -71.565 80.755 -71.235 81.085 ;
        RECT -71.565 79.395 -71.235 79.725 ;
        RECT -71.565 78.035 -71.235 78.365 ;
        RECT -71.565 76.675 -71.235 77.005 ;
        RECT -71.565 75.315 -71.235 75.645 ;
        RECT -71.565 73.955 -71.235 74.285 ;
        RECT -71.565 72.595 -71.235 72.925 ;
        RECT -71.565 71.235 -71.235 71.565 ;
        RECT -71.565 69.875 -71.235 70.205 ;
        RECT -71.565 68.515 -71.235 68.845 ;
        RECT -71.565 67.155 -71.235 67.485 ;
        RECT -71.565 65.795 -71.235 66.125 ;
        RECT -71.565 64.435 -71.235 64.765 ;
        RECT -71.565 63.075 -71.235 63.405 ;
        RECT -71.565 61.715 -71.235 62.045 ;
        RECT -71.565 60.355 -71.235 60.685 ;
        RECT -71.565 58.995 -71.235 59.325 ;
        RECT -71.565 57.635 -71.235 57.965 ;
        RECT -71.565 56.275 -71.235 56.605 ;
        RECT -71.565 54.915 -71.235 55.245 ;
        RECT -71.565 53.555 -71.235 53.885 ;
        RECT -71.565 52.195 -71.235 52.525 ;
        RECT -71.565 50.835 -71.235 51.165 ;
        RECT -71.565 49.475 -71.235 49.805 ;
        RECT -71.565 48.115 -71.235 48.445 ;
        RECT -71.565 46.755 -71.235 47.085 ;
        RECT -71.565 45.395 -71.235 45.725 ;
        RECT -71.565 44.035 -71.235 44.365 ;
        RECT -71.565 42.675 -71.235 43.005 ;
        RECT -71.565 41.315 -71.235 41.645 ;
        RECT -71.565 39.955 -71.235 40.285 ;
        RECT -71.565 38.595 -71.235 38.925 ;
        RECT -71.565 37.235 -71.235 37.565 ;
        RECT -71.565 35.875 -71.235 36.205 ;
        RECT -71.565 34.515 -71.235 34.845 ;
        RECT -71.565 33.155 -71.235 33.485 ;
        RECT -71.565 31.795 -71.235 32.125 ;
        RECT -71.565 30.435 -71.235 30.765 ;
        RECT -71.565 29.075 -71.235 29.405 ;
        RECT -71.565 27.715 -71.235 28.045 ;
        RECT -71.565 26.355 -71.235 26.685 ;
        RECT -71.565 24.995 -71.235 25.325 ;
        RECT -71.565 23.635 -71.235 23.965 ;
        RECT -71.565 22.275 -71.235 22.605 ;
        RECT -71.565 20.915 -71.235 21.245 ;
        RECT -71.565 19.555 -71.235 19.885 ;
        RECT -71.565 18.195 -71.235 18.525 ;
        RECT -71.565 16.835 -71.235 17.165 ;
        RECT -71.565 15.475 -71.235 15.805 ;
        RECT -71.565 14.115 -71.235 14.445 ;
        RECT -71.565 12.755 -71.235 13.085 ;
        RECT -71.565 11.395 -71.235 11.725 ;
        RECT -71.565 10.035 -71.235 10.365 ;
        RECT -71.565 8.675 -71.235 9.005 ;
        RECT -71.565 7.315 -71.235 7.645 ;
        RECT -71.565 5.955 -71.235 6.285 ;
        RECT -71.565 4.595 -71.235 4.925 ;
        RECT -71.565 3.235 -71.235 3.565 ;
        RECT -71.565 1.875 -71.235 2.205 ;
        RECT -71.565 0.515 -71.235 0.845 ;
        RECT -71.565 -0.845 -71.235 -0.515 ;
        RECT -71.565 -2.205 -71.235 -1.875 ;
        RECT -71.565 -3.565 -71.235 -3.235 ;
        RECT -71.565 -4.925 -71.235 -4.595 ;
        RECT -71.565 -6.285 -71.235 -5.955 ;
        RECT -71.565 -7.645 -71.235 -7.315 ;
        RECT -71.565 -9.005 -71.235 -8.675 ;
        RECT -71.565 -10.365 -71.235 -10.035 ;
        RECT -71.565 -11.725 -71.235 -11.395 ;
        RECT -71.565 -13.085 -71.235 -12.755 ;
        RECT -71.565 -14.445 -71.235 -14.115 ;
        RECT -71.565 -15.805 -71.235 -15.475 ;
        RECT -71.565 -17.165 -71.235 -16.835 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 398.315 241.32 398.645 242.45 ;
        RECT 398.315 239.195 398.645 239.525 ;
        RECT 398.315 237.835 398.645 238.165 ;
        RECT 398.315 235.975 398.645 236.305 ;
        RECT 398.315 233.925 398.645 234.255 ;
        RECT 398.315 231.995 398.645 232.325 ;
        RECT 398.315 230.155 398.645 230.485 ;
        RECT 398.315 228.665 398.645 228.995 ;
        RECT 398.315 226.995 398.645 227.325 ;
        RECT 398.315 225.505 398.645 225.835 ;
        RECT 398.315 223.835 398.645 224.165 ;
        RECT 398.315 222.345 398.645 222.675 ;
        RECT 398.315 220.675 398.645 221.005 ;
        RECT 398.315 219.185 398.645 219.515 ;
        RECT 398.315 217.775 398.645 218.105 ;
        RECT 398.315 215.935 398.645 216.265 ;
        RECT 398.315 214.445 398.645 214.775 ;
        RECT 398.315 212.775 398.645 213.105 ;
        RECT 398.315 211.285 398.645 211.615 ;
        RECT 398.315 209.615 398.645 209.945 ;
        RECT 398.315 208.125 398.645 208.455 ;
        RECT 398.315 206.455 398.645 206.785 ;
        RECT 398.315 204.965 398.645 205.295 ;
        RECT 398.315 203.555 398.645 203.885 ;
        RECT 398.315 201.715 398.645 202.045 ;
        RECT 398.315 200.225 398.645 200.555 ;
        RECT 398.315 198.555 398.645 198.885 ;
        RECT 398.315 197.065 398.645 197.395 ;
        RECT 398.315 195.395 398.645 195.725 ;
        RECT 398.315 193.905 398.645 194.235 ;
        RECT 398.315 192.235 398.645 192.565 ;
        RECT 398.315 190.745 398.645 191.075 ;
        RECT 398.315 189.335 398.645 189.665 ;
        RECT 398.315 187.495 398.645 187.825 ;
        RECT 398.315 186.005 398.645 186.335 ;
        RECT 398.315 184.335 398.645 184.665 ;
        RECT 398.315 182.845 398.645 183.175 ;
        RECT 398.315 181.175 398.645 181.505 ;
        RECT 398.315 179.685 398.645 180.015 ;
        RECT 398.315 178.015 398.645 178.345 ;
        RECT 398.315 176.525 398.645 176.855 ;
        RECT 398.315 175.115 398.645 175.445 ;
        RECT 398.315 173.275 398.645 173.605 ;
        RECT 398.315 171.785 398.645 172.115 ;
        RECT 398.315 170.115 398.645 170.445 ;
        RECT 398.315 168.625 398.645 168.955 ;
        RECT 398.315 166.955 398.645 167.285 ;
        RECT 398.315 165.465 398.645 165.795 ;
        RECT 398.315 163.795 398.645 164.125 ;
        RECT 398.315 162.305 398.645 162.635 ;
        RECT 398.315 160.895 398.645 161.225 ;
        RECT 398.315 159.055 398.645 159.385 ;
        RECT 398.315 157.565 398.645 157.895 ;
        RECT 398.315 155.895 398.645 156.225 ;
        RECT 398.315 154.405 398.645 154.735 ;
        RECT 398.315 152.735 398.645 153.065 ;
        RECT 398.315 151.245 398.645 151.575 ;
        RECT 398.315 149.575 398.645 149.905 ;
        RECT 398.315 148.085 398.645 148.415 ;
        RECT 398.315 146.675 398.645 147.005 ;
        RECT 398.315 144.835 398.645 145.165 ;
        RECT 398.315 143.345 398.645 143.675 ;
        RECT 398.315 141.675 398.645 142.005 ;
        RECT 398.315 140.185 398.645 140.515 ;
        RECT 398.315 138.515 398.645 138.845 ;
        RECT 398.315 137.025 398.645 137.355 ;
        RECT 398.315 135.355 398.645 135.685 ;
        RECT 398.315 133.865 398.645 134.195 ;
        RECT 398.315 132.455 398.645 132.785 ;
        RECT 398.315 130.615 398.645 130.945 ;
        RECT 398.315 129.125 398.645 129.455 ;
        RECT 398.315 127.455 398.645 127.785 ;
        RECT 398.315 125.965 398.645 126.295 ;
        RECT 398.315 124.295 398.645 124.625 ;
        RECT 398.315 122.805 398.645 123.135 ;
        RECT 398.315 121.135 398.645 121.465 ;
        RECT 398.315 119.645 398.645 119.975 ;
        RECT 398.315 118.235 398.645 118.565 ;
        RECT 398.315 116.395 398.645 116.725 ;
        RECT 398.315 114.905 398.645 115.235 ;
        RECT 398.315 113.235 398.645 113.565 ;
        RECT 398.315 111.745 398.645 112.075 ;
        RECT 398.315 110.075 398.645 110.405 ;
        RECT 398.315 108.585 398.645 108.915 ;
        RECT 398.315 106.915 398.645 107.245 ;
        RECT 398.315 105.425 398.645 105.755 ;
        RECT 398.315 104.015 398.645 104.345 ;
        RECT 398.315 102.175 398.645 102.505 ;
        RECT 398.315 100.685 398.645 101.015 ;
        RECT 398.315 99.015 398.645 99.345 ;
        RECT 398.315 97.525 398.645 97.855 ;
        RECT 398.315 95.855 398.645 96.185 ;
        RECT 398.315 94.365 398.645 94.695 ;
        RECT 398.315 92.695 398.645 93.025 ;
        RECT 398.315 91.205 398.645 91.535 ;
        RECT 398.315 89.795 398.645 90.125 ;
        RECT 398.315 87.955 398.645 88.285 ;
        RECT 398.315 86.465 398.645 86.795 ;
        RECT 398.315 84.795 398.645 85.125 ;
        RECT 398.315 83.305 398.645 83.635 ;
        RECT 398.315 81.635 398.645 81.965 ;
        RECT 398.315 80.145 398.645 80.475 ;
        RECT 398.315 78.475 398.645 78.805 ;
        RECT 398.315 76.985 398.645 77.315 ;
        RECT 398.315 75.575 398.645 75.905 ;
        RECT 398.315 73.735 398.645 74.065 ;
        RECT 398.315 72.245 398.645 72.575 ;
        RECT 398.315 70.575 398.645 70.905 ;
        RECT 398.315 69.085 398.645 69.415 ;
        RECT 398.315 67.415 398.645 67.745 ;
        RECT 398.315 65.925 398.645 66.255 ;
        RECT 398.315 64.255 398.645 64.585 ;
        RECT 398.315 62.765 398.645 63.095 ;
        RECT 398.315 61.355 398.645 61.685 ;
        RECT 398.315 59.515 398.645 59.845 ;
        RECT 398.315 58.025 398.645 58.355 ;
        RECT 398.315 56.355 398.645 56.685 ;
        RECT 398.315 54.865 398.645 55.195 ;
        RECT 398.315 53.195 398.645 53.525 ;
        RECT 398.315 51.705 398.645 52.035 ;
        RECT 398.315 50.035 398.645 50.365 ;
        RECT 398.315 48.545 398.645 48.875 ;
        RECT 398.315 47.135 398.645 47.465 ;
        RECT 398.315 45.295 398.645 45.625 ;
        RECT 398.315 43.805 398.645 44.135 ;
        RECT 398.315 42.135 398.645 42.465 ;
        RECT 398.315 40.645 398.645 40.975 ;
        RECT 398.315 38.975 398.645 39.305 ;
        RECT 398.315 37.485 398.645 37.815 ;
        RECT 398.315 35.815 398.645 36.145 ;
        RECT 398.315 34.325 398.645 34.655 ;
        RECT 398.315 32.915 398.645 33.245 ;
        RECT 398.315 31.075 398.645 31.405 ;
        RECT 398.315 29.585 398.645 29.915 ;
        RECT 398.315 27.915 398.645 28.245 ;
        RECT 398.315 26.425 398.645 26.755 ;
        RECT 398.315 24.755 398.645 25.085 ;
        RECT 398.315 23.265 398.645 23.595 ;
        RECT 398.315 21.595 398.645 21.925 ;
        RECT 398.315 20.105 398.645 20.435 ;
        RECT 398.315 18.695 398.645 19.025 ;
        RECT 398.315 16.855 398.645 17.185 ;
        RECT 398.315 15.365 398.645 15.695 ;
        RECT 398.315 13.695 398.645 14.025 ;
        RECT 398.315 12.205 398.645 12.535 ;
        RECT 398.315 10.535 398.645 10.865 ;
        RECT 398.315 9.045 398.645 9.375 ;
        RECT 398.315 7.375 398.645 7.705 ;
        RECT 398.315 5.885 398.645 6.215 ;
        RECT 398.315 4.475 398.645 4.805 ;
        RECT 398.315 2.115 398.645 2.445 ;
        RECT 398.315 0.06 398.645 0.39 ;
        RECT 398.315 -1.525 398.645 -1.195 ;
        RECT 398.315 -2.885 398.645 -2.555 ;
        RECT 398.315 -4.245 398.645 -3.915 ;
        RECT 398.315 -5.605 398.645 -5.275 ;
        RECT 398.315 -6.965 398.645 -6.635 ;
        RECT 398.315 -8.325 398.645 -7.995 ;
        RECT 398.315 -9.685 398.645 -9.355 ;
        RECT 398.315 -11.045 398.645 -10.715 ;
        RECT 398.315 -12.405 398.645 -12.075 ;
        RECT 398.315 -13.765 398.645 -13.435 ;
        RECT 398.315 -15.125 398.645 -14.795 ;
        RECT 398.315 -16.485 398.645 -16.155 ;
        RECT 398.315 -17.845 398.645 -17.515 ;
        RECT 398.315 -19.205 398.645 -18.875 ;
        RECT 398.315 -20.565 398.645 -20.235 ;
        RECT 398.315 -21.925 398.645 -21.595 ;
        RECT 398.315 -23.285 398.645 -22.955 ;
        RECT 398.315 -24.645 398.645 -24.315 ;
        RECT 398.315 -26.005 398.645 -25.675 ;
        RECT 398.315 -27.365 398.645 -27.035 ;
        RECT 398.315 -28.725 398.645 -28.395 ;
        RECT 398.315 -30.085 398.645 -29.755 ;
        RECT 398.315 -31.445 398.645 -31.115 ;
        RECT 398.315 -32.805 398.645 -32.475 ;
        RECT 398.315 -34.165 398.645 -33.835 ;
        RECT 398.315 -35.525 398.645 -35.195 ;
        RECT 398.315 -36.885 398.645 -36.555 ;
        RECT 398.315 -38.245 398.645 -37.915 ;
        RECT 398.315 -39.605 398.645 -39.275 ;
        RECT 398.315 -40.965 398.645 -40.635 ;
        RECT 398.315 -42.325 398.645 -41.995 ;
        RECT 398.315 -43.685 398.645 -43.355 ;
        RECT 398.315 -45.045 398.645 -44.715 ;
        RECT 398.315 -46.405 398.645 -46.075 ;
        RECT 398.315 -47.765 398.645 -47.435 ;
        RECT 398.315 -49.125 398.645 -48.795 ;
        RECT 398.315 -50.485 398.645 -50.155 ;
        RECT 398.315 -51.845 398.645 -51.515 ;
        RECT 398.315 -53.205 398.645 -52.875 ;
        RECT 398.315 -54.565 398.645 -54.235 ;
        RECT 398.315 -55.925 398.645 -55.595 ;
        RECT 398.315 -57.285 398.645 -56.955 ;
        RECT 398.315 -58.645 398.645 -58.315 ;
        RECT 398.315 -60.005 398.645 -59.675 ;
        RECT 398.315 -61.365 398.645 -61.035 ;
        RECT 398.315 -62.725 398.645 -62.395 ;
        RECT 398.315 -64.085 398.645 -63.755 ;
        RECT 398.315 -65.445 398.645 -65.115 ;
        RECT 398.315 -66.805 398.645 -66.475 ;
        RECT 398.315 -68.165 398.645 -67.835 ;
        RECT 398.315 -69.525 398.645 -69.195 ;
        RECT 398.315 -70.885 398.645 -70.555 ;
        RECT 398.315 -72.245 398.645 -71.915 ;
        RECT 398.315 -73.605 398.645 -73.275 ;
        RECT 398.315 -74.965 398.645 -74.635 ;
        RECT 398.315 -76.325 398.645 -75.995 ;
        RECT 398.315 -77.685 398.645 -77.355 ;
        RECT 398.315 -79.045 398.645 -78.715 ;
        RECT 398.315 -80.405 398.645 -80.075 ;
        RECT 398.315 -81.765 398.645 -81.435 ;
        RECT 398.315 -83.125 398.645 -82.795 ;
        RECT 398.315 -84.485 398.645 -84.155 ;
        RECT 398.315 -85.845 398.645 -85.515 ;
        RECT 398.315 -87.205 398.645 -86.875 ;
        RECT 398.315 -88.565 398.645 -88.235 ;
        RECT 398.315 -89.925 398.645 -89.595 ;
        RECT 398.315 -91.285 398.645 -90.955 ;
        RECT 398.315 -92.645 398.645 -92.315 ;
        RECT 398.315 -94.005 398.645 -93.675 ;
        RECT 398.315 -95.365 398.645 -95.035 ;
        RECT 398.315 -96.725 398.645 -96.395 ;
        RECT 398.315 -98.085 398.645 -97.755 ;
        RECT 398.315 -99.445 398.645 -99.115 ;
        RECT 398.315 -100.805 398.645 -100.475 ;
        RECT 398.315 -102.165 398.645 -101.835 ;
        RECT 398.315 -103.525 398.645 -103.195 ;
        RECT 398.315 -104.885 398.645 -104.555 ;
        RECT 398.315 -106.245 398.645 -105.915 ;
        RECT 398.315 -107.605 398.645 -107.275 ;
        RECT 398.315 -108.965 398.645 -108.635 ;
        RECT 398.315 -110.325 398.645 -109.995 ;
        RECT 398.315 -111.685 398.645 -111.355 ;
        RECT 398.315 -113.045 398.645 -112.715 ;
        RECT 398.315 -114.405 398.645 -114.075 ;
        RECT 398.315 -115.765 398.645 -115.435 ;
        RECT 398.315 -117.125 398.645 -116.795 ;
        RECT 398.315 -118.485 398.645 -118.155 ;
        RECT 398.315 -119.845 398.645 -119.515 ;
        RECT 398.315 -121.205 398.645 -120.875 ;
        RECT 398.315 -122.565 398.645 -122.235 ;
        RECT 398.315 -123.925 398.645 -123.595 ;
        RECT 398.315 -125.285 398.645 -124.955 ;
        RECT 398.315 -126.645 398.645 -126.315 ;
        RECT 398.315 -128.005 398.645 -127.675 ;
        RECT 398.315 -129.365 398.645 -129.035 ;
        RECT 398.315 -130.725 398.645 -130.395 ;
        RECT 398.315 -132.085 398.645 -131.755 ;
        RECT 398.315 -133.445 398.645 -133.115 ;
        RECT 398.315 -134.805 398.645 -134.475 ;
        RECT 398.315 -136.165 398.645 -135.835 ;
        RECT 398.315 -137.525 398.645 -137.195 ;
        RECT 398.315 -138.885 398.645 -138.555 ;
        RECT 398.315 -140.245 398.645 -139.915 ;
        RECT 398.315 -141.605 398.645 -141.275 ;
        RECT 398.315 -142.965 398.645 -142.635 ;
        RECT 398.315 -144.325 398.645 -143.995 ;
        RECT 398.315 -145.685 398.645 -145.355 ;
        RECT 398.315 -147.045 398.645 -146.715 ;
        RECT 398.315 -148.405 398.645 -148.075 ;
        RECT 398.315 -149.765 398.645 -149.435 ;
        RECT 398.315 -151.125 398.645 -150.795 ;
        RECT 398.315 -152.485 398.645 -152.155 ;
        RECT 398.315 -153.845 398.645 -153.515 ;
        RECT 398.315 -155.205 398.645 -154.875 ;
        RECT 398.315 -156.565 398.645 -156.235 ;
        RECT 398.315 -157.925 398.645 -157.595 ;
        RECT 398.315 -159.285 398.645 -158.955 ;
        RECT 398.315 -160.645 398.645 -160.315 ;
        RECT 398.315 -162.005 398.645 -161.675 ;
        RECT 398.315 -163.365 398.645 -163.035 ;
        RECT 398.315 -164.725 398.645 -164.395 ;
        RECT 398.315 -166.085 398.645 -165.755 ;
        RECT 398.315 -167.445 398.645 -167.115 ;
        RECT 398.315 -168.805 398.645 -168.475 ;
        RECT 398.315 -170.165 398.645 -169.835 ;
        RECT 398.315 -171.525 398.645 -171.195 ;
        RECT 398.315 -172.885 398.645 -172.555 ;
        RECT 398.315 -174.245 398.645 -173.915 ;
        RECT 398.315 -175.605 398.645 -175.275 ;
        RECT 398.315 -176.965 398.645 -176.635 ;
        RECT 398.315 -178.325 398.645 -177.995 ;
        RECT 398.315 -180.57 398.645 -179.44 ;
        RECT 398.32 -180.685 398.64 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 399.675 241.32 400.005 242.45 ;
        RECT 399.675 239.195 400.005 239.525 ;
        RECT 399.675 237.835 400.005 238.165 ;
        RECT 399.675 235.975 400.005 236.305 ;
        RECT 399.675 233.925 400.005 234.255 ;
        RECT 399.675 231.995 400.005 232.325 ;
        RECT 399.675 230.155 400.005 230.485 ;
        RECT 399.675 228.665 400.005 228.995 ;
        RECT 399.675 226.995 400.005 227.325 ;
        RECT 399.675 225.505 400.005 225.835 ;
        RECT 399.675 223.835 400.005 224.165 ;
        RECT 399.675 222.345 400.005 222.675 ;
        RECT 399.675 220.675 400.005 221.005 ;
        RECT 399.675 219.185 400.005 219.515 ;
        RECT 399.675 217.775 400.005 218.105 ;
        RECT 399.675 215.935 400.005 216.265 ;
        RECT 399.675 214.445 400.005 214.775 ;
        RECT 399.675 212.775 400.005 213.105 ;
        RECT 399.675 211.285 400.005 211.615 ;
        RECT 399.675 209.615 400.005 209.945 ;
        RECT 399.675 208.125 400.005 208.455 ;
        RECT 399.675 206.455 400.005 206.785 ;
        RECT 399.675 204.965 400.005 205.295 ;
        RECT 399.675 203.555 400.005 203.885 ;
        RECT 399.675 201.715 400.005 202.045 ;
        RECT 399.675 200.225 400.005 200.555 ;
        RECT 399.675 198.555 400.005 198.885 ;
        RECT 399.675 197.065 400.005 197.395 ;
        RECT 399.675 195.395 400.005 195.725 ;
        RECT 399.675 193.905 400.005 194.235 ;
        RECT 399.675 192.235 400.005 192.565 ;
        RECT 399.675 190.745 400.005 191.075 ;
        RECT 399.675 189.335 400.005 189.665 ;
        RECT 399.675 187.495 400.005 187.825 ;
        RECT 399.675 186.005 400.005 186.335 ;
        RECT 399.675 184.335 400.005 184.665 ;
        RECT 399.675 182.845 400.005 183.175 ;
        RECT 399.675 181.175 400.005 181.505 ;
        RECT 399.675 179.685 400.005 180.015 ;
        RECT 399.675 178.015 400.005 178.345 ;
        RECT 399.675 176.525 400.005 176.855 ;
        RECT 399.675 175.115 400.005 175.445 ;
        RECT 399.675 173.275 400.005 173.605 ;
        RECT 399.675 171.785 400.005 172.115 ;
        RECT 399.675 170.115 400.005 170.445 ;
        RECT 399.675 168.625 400.005 168.955 ;
        RECT 399.675 166.955 400.005 167.285 ;
        RECT 399.675 165.465 400.005 165.795 ;
        RECT 399.675 163.795 400.005 164.125 ;
        RECT 399.675 162.305 400.005 162.635 ;
        RECT 399.675 160.895 400.005 161.225 ;
        RECT 399.675 159.055 400.005 159.385 ;
        RECT 399.675 157.565 400.005 157.895 ;
        RECT 399.675 155.895 400.005 156.225 ;
        RECT 399.675 154.405 400.005 154.735 ;
        RECT 399.675 152.735 400.005 153.065 ;
        RECT 399.675 151.245 400.005 151.575 ;
        RECT 399.675 149.575 400.005 149.905 ;
        RECT 399.675 148.085 400.005 148.415 ;
        RECT 399.675 146.675 400.005 147.005 ;
        RECT 399.675 144.835 400.005 145.165 ;
        RECT 399.675 143.345 400.005 143.675 ;
        RECT 399.675 141.675 400.005 142.005 ;
        RECT 399.675 140.185 400.005 140.515 ;
        RECT 399.675 138.515 400.005 138.845 ;
        RECT 399.675 137.025 400.005 137.355 ;
        RECT 399.675 135.355 400.005 135.685 ;
        RECT 399.675 133.865 400.005 134.195 ;
        RECT 399.675 132.455 400.005 132.785 ;
        RECT 399.675 130.615 400.005 130.945 ;
        RECT 399.675 129.125 400.005 129.455 ;
        RECT 399.675 127.455 400.005 127.785 ;
        RECT 399.675 125.965 400.005 126.295 ;
        RECT 399.675 124.295 400.005 124.625 ;
        RECT 399.675 122.805 400.005 123.135 ;
        RECT 399.675 121.135 400.005 121.465 ;
        RECT 399.675 119.645 400.005 119.975 ;
        RECT 399.675 118.235 400.005 118.565 ;
        RECT 399.675 116.395 400.005 116.725 ;
        RECT 399.675 114.905 400.005 115.235 ;
        RECT 399.675 113.235 400.005 113.565 ;
        RECT 399.675 111.745 400.005 112.075 ;
        RECT 399.675 110.075 400.005 110.405 ;
        RECT 399.675 108.585 400.005 108.915 ;
        RECT 399.675 106.915 400.005 107.245 ;
        RECT 399.675 105.425 400.005 105.755 ;
        RECT 399.675 104.015 400.005 104.345 ;
        RECT 399.675 102.175 400.005 102.505 ;
        RECT 399.675 100.685 400.005 101.015 ;
        RECT 399.675 99.015 400.005 99.345 ;
        RECT 399.675 97.525 400.005 97.855 ;
        RECT 399.675 95.855 400.005 96.185 ;
        RECT 399.675 94.365 400.005 94.695 ;
        RECT 399.675 92.695 400.005 93.025 ;
        RECT 399.675 91.205 400.005 91.535 ;
        RECT 399.675 89.795 400.005 90.125 ;
        RECT 399.675 87.955 400.005 88.285 ;
        RECT 399.675 86.465 400.005 86.795 ;
        RECT 399.675 84.795 400.005 85.125 ;
        RECT 399.675 83.305 400.005 83.635 ;
        RECT 399.675 81.635 400.005 81.965 ;
        RECT 399.675 80.145 400.005 80.475 ;
        RECT 399.675 78.475 400.005 78.805 ;
        RECT 399.675 76.985 400.005 77.315 ;
        RECT 399.675 75.575 400.005 75.905 ;
        RECT 399.675 73.735 400.005 74.065 ;
        RECT 399.675 72.245 400.005 72.575 ;
        RECT 399.675 70.575 400.005 70.905 ;
        RECT 399.675 69.085 400.005 69.415 ;
        RECT 399.675 67.415 400.005 67.745 ;
        RECT 399.675 65.925 400.005 66.255 ;
        RECT 399.675 64.255 400.005 64.585 ;
        RECT 399.675 62.765 400.005 63.095 ;
        RECT 399.675 61.355 400.005 61.685 ;
        RECT 399.675 59.515 400.005 59.845 ;
        RECT 399.675 58.025 400.005 58.355 ;
        RECT 399.675 56.355 400.005 56.685 ;
        RECT 399.675 54.865 400.005 55.195 ;
        RECT 399.675 53.195 400.005 53.525 ;
        RECT 399.675 51.705 400.005 52.035 ;
        RECT 399.675 50.035 400.005 50.365 ;
        RECT 399.675 48.545 400.005 48.875 ;
        RECT 399.675 47.135 400.005 47.465 ;
        RECT 399.675 45.295 400.005 45.625 ;
        RECT 399.675 43.805 400.005 44.135 ;
        RECT 399.675 42.135 400.005 42.465 ;
        RECT 399.675 40.645 400.005 40.975 ;
        RECT 399.675 38.975 400.005 39.305 ;
        RECT 399.675 37.485 400.005 37.815 ;
        RECT 399.675 35.815 400.005 36.145 ;
        RECT 399.675 34.325 400.005 34.655 ;
        RECT 399.675 32.915 400.005 33.245 ;
        RECT 399.675 31.075 400.005 31.405 ;
        RECT 399.675 29.585 400.005 29.915 ;
        RECT 399.675 27.915 400.005 28.245 ;
        RECT 399.675 26.425 400.005 26.755 ;
        RECT 399.675 24.755 400.005 25.085 ;
        RECT 399.675 23.265 400.005 23.595 ;
        RECT 399.675 21.595 400.005 21.925 ;
        RECT 399.675 20.105 400.005 20.435 ;
        RECT 399.675 18.695 400.005 19.025 ;
        RECT 399.675 16.855 400.005 17.185 ;
        RECT 399.675 15.365 400.005 15.695 ;
        RECT 399.675 13.695 400.005 14.025 ;
        RECT 399.675 12.205 400.005 12.535 ;
        RECT 399.675 10.535 400.005 10.865 ;
        RECT 399.675 9.045 400.005 9.375 ;
        RECT 399.675 7.375 400.005 7.705 ;
        RECT 399.675 5.885 400.005 6.215 ;
        RECT 399.675 4.475 400.005 4.805 ;
        RECT 399.675 2.115 400.005 2.445 ;
        RECT 399.675 0.06 400.005 0.39 ;
        RECT 399.675 -1.525 400.005 -1.195 ;
        RECT 399.675 -2.885 400.005 -2.555 ;
        RECT 399.675 -4.245 400.005 -3.915 ;
        RECT 399.675 -5.605 400.005 -5.275 ;
        RECT 399.675 -6.965 400.005 -6.635 ;
        RECT 399.675 -8.325 400.005 -7.995 ;
        RECT 399.675 -9.685 400.005 -9.355 ;
        RECT 399.675 -11.045 400.005 -10.715 ;
        RECT 399.675 -12.405 400.005 -12.075 ;
        RECT 399.675 -13.765 400.005 -13.435 ;
        RECT 399.675 -15.125 400.005 -14.795 ;
        RECT 399.675 -16.485 400.005 -16.155 ;
        RECT 399.675 -17.845 400.005 -17.515 ;
        RECT 399.675 -19.205 400.005 -18.875 ;
        RECT 399.675 -20.565 400.005 -20.235 ;
        RECT 399.675 -21.925 400.005 -21.595 ;
        RECT 399.675 -23.285 400.005 -22.955 ;
        RECT 399.675 -24.645 400.005 -24.315 ;
        RECT 399.675 -26.005 400.005 -25.675 ;
        RECT 399.675 -27.365 400.005 -27.035 ;
        RECT 399.675 -28.725 400.005 -28.395 ;
        RECT 399.675 -30.085 400.005 -29.755 ;
        RECT 399.675 -31.445 400.005 -31.115 ;
        RECT 399.675 -32.805 400.005 -32.475 ;
        RECT 399.675 -34.165 400.005 -33.835 ;
        RECT 399.675 -35.525 400.005 -35.195 ;
        RECT 399.675 -36.885 400.005 -36.555 ;
        RECT 399.675 -38.245 400.005 -37.915 ;
        RECT 399.675 -39.605 400.005 -39.275 ;
        RECT 399.675 -40.965 400.005 -40.635 ;
        RECT 399.675 -42.325 400.005 -41.995 ;
        RECT 399.675 -43.685 400.005 -43.355 ;
        RECT 399.675 -45.045 400.005 -44.715 ;
        RECT 399.675 -46.405 400.005 -46.075 ;
        RECT 399.675 -47.765 400.005 -47.435 ;
        RECT 399.675 -49.125 400.005 -48.795 ;
        RECT 399.675 -50.485 400.005 -50.155 ;
        RECT 399.675 -51.845 400.005 -51.515 ;
        RECT 399.675 -53.205 400.005 -52.875 ;
        RECT 399.675 -54.565 400.005 -54.235 ;
        RECT 399.675 -55.925 400.005 -55.595 ;
        RECT 399.675 -57.285 400.005 -56.955 ;
        RECT 399.675 -58.645 400.005 -58.315 ;
        RECT 399.675 -60.005 400.005 -59.675 ;
        RECT 399.675 -61.365 400.005 -61.035 ;
        RECT 399.675 -62.725 400.005 -62.395 ;
        RECT 399.675 -64.085 400.005 -63.755 ;
        RECT 399.675 -65.445 400.005 -65.115 ;
        RECT 399.675 -66.805 400.005 -66.475 ;
        RECT 399.675 -68.165 400.005 -67.835 ;
        RECT 399.675 -69.525 400.005 -69.195 ;
        RECT 399.675 -70.885 400.005 -70.555 ;
        RECT 399.675 -72.245 400.005 -71.915 ;
        RECT 399.675 -73.605 400.005 -73.275 ;
        RECT 399.675 -74.965 400.005 -74.635 ;
        RECT 399.675 -76.325 400.005 -75.995 ;
        RECT 399.675 -77.685 400.005 -77.355 ;
        RECT 399.675 -79.045 400.005 -78.715 ;
        RECT 399.675 -80.405 400.005 -80.075 ;
        RECT 399.675 -81.765 400.005 -81.435 ;
        RECT 399.675 -83.125 400.005 -82.795 ;
        RECT 399.675 -84.485 400.005 -84.155 ;
        RECT 399.675 -85.845 400.005 -85.515 ;
        RECT 399.675 -87.205 400.005 -86.875 ;
        RECT 399.675 -88.565 400.005 -88.235 ;
        RECT 399.675 -89.925 400.005 -89.595 ;
        RECT 399.675 -91.285 400.005 -90.955 ;
        RECT 399.675 -92.645 400.005 -92.315 ;
        RECT 399.675 -94.005 400.005 -93.675 ;
        RECT 399.675 -95.365 400.005 -95.035 ;
        RECT 399.675 -96.725 400.005 -96.395 ;
        RECT 399.675 -98.085 400.005 -97.755 ;
        RECT 399.675 -99.445 400.005 -99.115 ;
        RECT 399.675 -100.805 400.005 -100.475 ;
        RECT 399.675 -102.165 400.005 -101.835 ;
        RECT 399.675 -103.525 400.005 -103.195 ;
        RECT 399.675 -104.885 400.005 -104.555 ;
        RECT 399.675 -106.245 400.005 -105.915 ;
        RECT 399.675 -107.605 400.005 -107.275 ;
        RECT 399.675 -108.965 400.005 -108.635 ;
        RECT 399.675 -110.325 400.005 -109.995 ;
        RECT 399.675 -111.685 400.005 -111.355 ;
        RECT 399.675 -113.045 400.005 -112.715 ;
        RECT 399.675 -114.405 400.005 -114.075 ;
        RECT 399.675 -115.765 400.005 -115.435 ;
        RECT 399.675 -117.125 400.005 -116.795 ;
        RECT 399.675 -118.485 400.005 -118.155 ;
        RECT 399.675 -119.845 400.005 -119.515 ;
        RECT 399.675 -121.205 400.005 -120.875 ;
        RECT 399.675 -122.565 400.005 -122.235 ;
        RECT 399.675 -123.925 400.005 -123.595 ;
        RECT 399.675 -125.285 400.005 -124.955 ;
        RECT 399.675 -126.645 400.005 -126.315 ;
        RECT 399.675 -128.005 400.005 -127.675 ;
        RECT 399.675 -129.365 400.005 -129.035 ;
        RECT 399.675 -130.725 400.005 -130.395 ;
        RECT 399.675 -132.085 400.005 -131.755 ;
        RECT 399.675 -133.445 400.005 -133.115 ;
        RECT 399.675 -134.805 400.005 -134.475 ;
        RECT 399.675 -136.165 400.005 -135.835 ;
        RECT 399.675 -137.525 400.005 -137.195 ;
        RECT 399.675 -138.885 400.005 -138.555 ;
        RECT 399.675 -140.245 400.005 -139.915 ;
        RECT 399.675 -141.605 400.005 -141.275 ;
        RECT 399.675 -142.965 400.005 -142.635 ;
        RECT 399.675 -144.325 400.005 -143.995 ;
        RECT 399.675 -145.685 400.005 -145.355 ;
        RECT 399.675 -147.045 400.005 -146.715 ;
        RECT 399.675 -148.405 400.005 -148.075 ;
        RECT 399.675 -149.765 400.005 -149.435 ;
        RECT 399.675 -151.125 400.005 -150.795 ;
        RECT 399.675 -152.485 400.005 -152.155 ;
        RECT 399.675 -153.845 400.005 -153.515 ;
        RECT 399.675 -155.205 400.005 -154.875 ;
        RECT 399.675 -156.565 400.005 -156.235 ;
        RECT 399.675 -157.925 400.005 -157.595 ;
        RECT 399.675 -159.285 400.005 -158.955 ;
        RECT 399.675 -160.645 400.005 -160.315 ;
        RECT 399.675 -162.005 400.005 -161.675 ;
        RECT 399.675 -163.365 400.005 -163.035 ;
        RECT 399.675 -164.725 400.005 -164.395 ;
        RECT 399.675 -166.085 400.005 -165.755 ;
        RECT 399.675 -167.445 400.005 -167.115 ;
        RECT 399.675 -168.805 400.005 -168.475 ;
        RECT 399.675 -170.165 400.005 -169.835 ;
        RECT 399.675 -171.525 400.005 -171.195 ;
        RECT 399.675 -172.885 400.005 -172.555 ;
        RECT 399.675 -174.245 400.005 -173.915 ;
        RECT 399.675 -175.605 400.005 -175.275 ;
        RECT 399.675 -176.965 400.005 -176.635 ;
        RECT 399.675 -178.325 400.005 -177.995 ;
        RECT 399.675 -180.57 400.005 -179.44 ;
        RECT 399.68 -180.685 400 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 401.035 241.32 401.365 242.45 ;
        RECT 401.035 239.195 401.365 239.525 ;
        RECT 401.035 237.835 401.365 238.165 ;
        RECT 401.035 235.975 401.365 236.305 ;
        RECT 401.035 233.925 401.365 234.255 ;
        RECT 401.035 231.995 401.365 232.325 ;
        RECT 401.035 230.155 401.365 230.485 ;
        RECT 401.035 228.665 401.365 228.995 ;
        RECT 401.035 226.995 401.365 227.325 ;
        RECT 401.035 225.505 401.365 225.835 ;
        RECT 401.035 223.835 401.365 224.165 ;
        RECT 401.035 222.345 401.365 222.675 ;
        RECT 401.035 220.675 401.365 221.005 ;
        RECT 401.035 219.185 401.365 219.515 ;
        RECT 401.035 217.775 401.365 218.105 ;
        RECT 401.035 215.935 401.365 216.265 ;
        RECT 401.035 214.445 401.365 214.775 ;
        RECT 401.035 212.775 401.365 213.105 ;
        RECT 401.035 211.285 401.365 211.615 ;
        RECT 401.035 209.615 401.365 209.945 ;
        RECT 401.035 208.125 401.365 208.455 ;
        RECT 401.035 206.455 401.365 206.785 ;
        RECT 401.035 204.965 401.365 205.295 ;
        RECT 401.035 203.555 401.365 203.885 ;
        RECT 401.035 201.715 401.365 202.045 ;
        RECT 401.035 200.225 401.365 200.555 ;
        RECT 401.035 198.555 401.365 198.885 ;
        RECT 401.035 197.065 401.365 197.395 ;
        RECT 401.035 195.395 401.365 195.725 ;
        RECT 401.035 193.905 401.365 194.235 ;
        RECT 401.035 192.235 401.365 192.565 ;
        RECT 401.035 190.745 401.365 191.075 ;
        RECT 401.035 189.335 401.365 189.665 ;
        RECT 401.035 187.495 401.365 187.825 ;
        RECT 401.035 186.005 401.365 186.335 ;
        RECT 401.035 184.335 401.365 184.665 ;
        RECT 401.035 182.845 401.365 183.175 ;
        RECT 401.035 181.175 401.365 181.505 ;
        RECT 401.035 179.685 401.365 180.015 ;
        RECT 401.035 178.015 401.365 178.345 ;
        RECT 401.035 176.525 401.365 176.855 ;
        RECT 401.035 175.115 401.365 175.445 ;
        RECT 401.035 173.275 401.365 173.605 ;
        RECT 401.035 171.785 401.365 172.115 ;
        RECT 401.035 170.115 401.365 170.445 ;
        RECT 401.035 168.625 401.365 168.955 ;
        RECT 401.035 166.955 401.365 167.285 ;
        RECT 401.035 165.465 401.365 165.795 ;
        RECT 401.035 163.795 401.365 164.125 ;
        RECT 401.035 162.305 401.365 162.635 ;
        RECT 401.035 160.895 401.365 161.225 ;
        RECT 401.035 159.055 401.365 159.385 ;
        RECT 401.035 157.565 401.365 157.895 ;
        RECT 401.035 155.895 401.365 156.225 ;
        RECT 401.035 154.405 401.365 154.735 ;
        RECT 401.035 152.735 401.365 153.065 ;
        RECT 401.035 151.245 401.365 151.575 ;
        RECT 401.035 149.575 401.365 149.905 ;
        RECT 401.035 148.085 401.365 148.415 ;
        RECT 401.035 146.675 401.365 147.005 ;
        RECT 401.035 144.835 401.365 145.165 ;
        RECT 401.035 143.345 401.365 143.675 ;
        RECT 401.035 141.675 401.365 142.005 ;
        RECT 401.035 140.185 401.365 140.515 ;
        RECT 401.035 138.515 401.365 138.845 ;
        RECT 401.035 137.025 401.365 137.355 ;
        RECT 401.035 135.355 401.365 135.685 ;
        RECT 401.035 133.865 401.365 134.195 ;
        RECT 401.035 132.455 401.365 132.785 ;
        RECT 401.035 130.615 401.365 130.945 ;
        RECT 401.035 129.125 401.365 129.455 ;
        RECT 401.035 127.455 401.365 127.785 ;
        RECT 401.035 125.965 401.365 126.295 ;
        RECT 401.035 124.295 401.365 124.625 ;
        RECT 401.035 122.805 401.365 123.135 ;
        RECT 401.035 121.135 401.365 121.465 ;
        RECT 401.035 119.645 401.365 119.975 ;
        RECT 401.035 118.235 401.365 118.565 ;
        RECT 401.035 116.395 401.365 116.725 ;
        RECT 401.035 114.905 401.365 115.235 ;
        RECT 401.035 113.235 401.365 113.565 ;
        RECT 401.035 111.745 401.365 112.075 ;
        RECT 401.035 110.075 401.365 110.405 ;
        RECT 401.035 108.585 401.365 108.915 ;
        RECT 401.035 106.915 401.365 107.245 ;
        RECT 401.035 105.425 401.365 105.755 ;
        RECT 401.035 104.015 401.365 104.345 ;
        RECT 401.035 102.175 401.365 102.505 ;
        RECT 401.035 100.685 401.365 101.015 ;
        RECT 401.035 99.015 401.365 99.345 ;
        RECT 401.035 97.525 401.365 97.855 ;
        RECT 401.035 95.855 401.365 96.185 ;
        RECT 401.035 94.365 401.365 94.695 ;
        RECT 401.035 92.695 401.365 93.025 ;
        RECT 401.035 91.205 401.365 91.535 ;
        RECT 401.035 89.795 401.365 90.125 ;
        RECT 401.035 87.955 401.365 88.285 ;
        RECT 401.035 86.465 401.365 86.795 ;
        RECT 401.035 84.795 401.365 85.125 ;
        RECT 401.035 83.305 401.365 83.635 ;
        RECT 401.035 81.635 401.365 81.965 ;
        RECT 401.035 80.145 401.365 80.475 ;
        RECT 401.035 78.475 401.365 78.805 ;
        RECT 401.035 76.985 401.365 77.315 ;
        RECT 401.035 75.575 401.365 75.905 ;
        RECT 401.035 73.735 401.365 74.065 ;
        RECT 401.035 72.245 401.365 72.575 ;
        RECT 401.035 70.575 401.365 70.905 ;
        RECT 401.035 69.085 401.365 69.415 ;
        RECT 401.035 67.415 401.365 67.745 ;
        RECT 401.035 65.925 401.365 66.255 ;
        RECT 401.035 64.255 401.365 64.585 ;
        RECT 401.035 62.765 401.365 63.095 ;
        RECT 401.035 61.355 401.365 61.685 ;
        RECT 401.035 59.515 401.365 59.845 ;
        RECT 401.035 58.025 401.365 58.355 ;
        RECT 401.035 56.355 401.365 56.685 ;
        RECT 401.035 54.865 401.365 55.195 ;
        RECT 401.035 53.195 401.365 53.525 ;
        RECT 401.035 51.705 401.365 52.035 ;
        RECT 401.035 50.035 401.365 50.365 ;
        RECT 401.035 48.545 401.365 48.875 ;
        RECT 401.035 47.135 401.365 47.465 ;
        RECT 401.035 45.295 401.365 45.625 ;
        RECT 401.035 43.805 401.365 44.135 ;
        RECT 401.035 42.135 401.365 42.465 ;
        RECT 401.035 40.645 401.365 40.975 ;
        RECT 401.035 38.975 401.365 39.305 ;
        RECT 401.035 37.485 401.365 37.815 ;
        RECT 401.035 35.815 401.365 36.145 ;
        RECT 401.035 34.325 401.365 34.655 ;
        RECT 401.035 32.915 401.365 33.245 ;
        RECT 401.035 31.075 401.365 31.405 ;
        RECT 401.035 29.585 401.365 29.915 ;
        RECT 401.035 27.915 401.365 28.245 ;
        RECT 401.035 26.425 401.365 26.755 ;
        RECT 401.035 24.755 401.365 25.085 ;
        RECT 401.035 23.265 401.365 23.595 ;
        RECT 401.035 21.595 401.365 21.925 ;
        RECT 401.035 20.105 401.365 20.435 ;
        RECT 401.035 18.695 401.365 19.025 ;
        RECT 401.035 16.855 401.365 17.185 ;
        RECT 401.035 15.365 401.365 15.695 ;
        RECT 401.035 13.695 401.365 14.025 ;
        RECT 401.035 12.205 401.365 12.535 ;
        RECT 401.035 10.535 401.365 10.865 ;
        RECT 401.035 9.045 401.365 9.375 ;
        RECT 401.035 7.375 401.365 7.705 ;
        RECT 401.035 5.885 401.365 6.215 ;
        RECT 401.035 4.475 401.365 4.805 ;
        RECT 401.035 2.115 401.365 2.445 ;
        RECT 401.035 0.06 401.365 0.39 ;
        RECT 401.035 -1.525 401.365 -1.195 ;
        RECT 401.035 -2.885 401.365 -2.555 ;
        RECT 401.035 -4.245 401.365 -3.915 ;
        RECT 401.035 -5.605 401.365 -5.275 ;
        RECT 401.035 -6.965 401.365 -6.635 ;
        RECT 401.035 -8.325 401.365 -7.995 ;
        RECT 401.035 -9.685 401.365 -9.355 ;
        RECT 401.035 -11.045 401.365 -10.715 ;
        RECT 401.035 -12.405 401.365 -12.075 ;
        RECT 401.035 -13.765 401.365 -13.435 ;
        RECT 401.035 -15.125 401.365 -14.795 ;
        RECT 401.035 -16.485 401.365 -16.155 ;
        RECT 401.035 -17.845 401.365 -17.515 ;
        RECT 401.035 -19.205 401.365 -18.875 ;
        RECT 401.035 -20.565 401.365 -20.235 ;
        RECT 401.035 -21.925 401.365 -21.595 ;
        RECT 401.035 -23.285 401.365 -22.955 ;
        RECT 401.035 -24.645 401.365 -24.315 ;
        RECT 401.035 -26.005 401.365 -25.675 ;
        RECT 401.035 -27.365 401.365 -27.035 ;
        RECT 401.035 -28.725 401.365 -28.395 ;
        RECT 401.035 -30.085 401.365 -29.755 ;
        RECT 401.035 -31.445 401.365 -31.115 ;
        RECT 401.035 -32.805 401.365 -32.475 ;
        RECT 401.035 -34.165 401.365 -33.835 ;
        RECT 401.035 -35.525 401.365 -35.195 ;
        RECT 401.035 -36.885 401.365 -36.555 ;
        RECT 401.035 -38.245 401.365 -37.915 ;
        RECT 401.035 -39.605 401.365 -39.275 ;
        RECT 401.035 -40.965 401.365 -40.635 ;
        RECT 401.035 -42.325 401.365 -41.995 ;
        RECT 401.035 -43.685 401.365 -43.355 ;
        RECT 401.035 -45.045 401.365 -44.715 ;
        RECT 401.035 -46.405 401.365 -46.075 ;
        RECT 401.035 -47.765 401.365 -47.435 ;
        RECT 401.035 -49.125 401.365 -48.795 ;
        RECT 401.035 -50.485 401.365 -50.155 ;
        RECT 401.035 -51.845 401.365 -51.515 ;
        RECT 401.035 -53.205 401.365 -52.875 ;
        RECT 401.035 -54.565 401.365 -54.235 ;
        RECT 401.035 -55.925 401.365 -55.595 ;
        RECT 401.035 -57.285 401.365 -56.955 ;
        RECT 401.035 -58.645 401.365 -58.315 ;
        RECT 401.035 -60.005 401.365 -59.675 ;
        RECT 401.035 -61.365 401.365 -61.035 ;
        RECT 401.035 -62.725 401.365 -62.395 ;
        RECT 401.035 -64.085 401.365 -63.755 ;
        RECT 401.035 -65.445 401.365 -65.115 ;
        RECT 401.035 -66.805 401.365 -66.475 ;
        RECT 401.035 -68.165 401.365 -67.835 ;
        RECT 401.035 -69.525 401.365 -69.195 ;
        RECT 401.035 -70.885 401.365 -70.555 ;
        RECT 401.035 -72.245 401.365 -71.915 ;
        RECT 401.035 -73.605 401.365 -73.275 ;
        RECT 401.035 -74.965 401.365 -74.635 ;
        RECT 401.035 -76.325 401.365 -75.995 ;
        RECT 401.035 -77.685 401.365 -77.355 ;
        RECT 401.035 -79.045 401.365 -78.715 ;
        RECT 401.035 -80.405 401.365 -80.075 ;
        RECT 401.035 -81.765 401.365 -81.435 ;
        RECT 401.035 -83.125 401.365 -82.795 ;
        RECT 401.035 -84.485 401.365 -84.155 ;
        RECT 401.035 -85.845 401.365 -85.515 ;
        RECT 401.035 -87.205 401.365 -86.875 ;
        RECT 401.035 -88.565 401.365 -88.235 ;
        RECT 401.035 -89.925 401.365 -89.595 ;
        RECT 401.035 -91.285 401.365 -90.955 ;
        RECT 401.035 -92.645 401.365 -92.315 ;
        RECT 401.035 -94.005 401.365 -93.675 ;
        RECT 401.035 -95.365 401.365 -95.035 ;
        RECT 401.035 -96.725 401.365 -96.395 ;
        RECT 401.035 -98.085 401.365 -97.755 ;
        RECT 401.035 -99.445 401.365 -99.115 ;
        RECT 401.035 -100.805 401.365 -100.475 ;
        RECT 401.035 -102.165 401.365 -101.835 ;
        RECT 401.035 -103.525 401.365 -103.195 ;
        RECT 401.035 -104.885 401.365 -104.555 ;
        RECT 401.035 -106.245 401.365 -105.915 ;
        RECT 401.035 -107.605 401.365 -107.275 ;
        RECT 401.035 -108.965 401.365 -108.635 ;
        RECT 401.035 -110.325 401.365 -109.995 ;
        RECT 401.035 -111.685 401.365 -111.355 ;
        RECT 401.035 -113.045 401.365 -112.715 ;
        RECT 401.035 -114.405 401.365 -114.075 ;
        RECT 401.035 -115.765 401.365 -115.435 ;
        RECT 401.035 -117.125 401.365 -116.795 ;
        RECT 401.035 -118.485 401.365 -118.155 ;
        RECT 401.035 -119.845 401.365 -119.515 ;
        RECT 401.035 -121.205 401.365 -120.875 ;
        RECT 401.035 -122.565 401.365 -122.235 ;
        RECT 401.035 -123.925 401.365 -123.595 ;
        RECT 401.035 -125.285 401.365 -124.955 ;
        RECT 401.035 -126.645 401.365 -126.315 ;
        RECT 401.035 -128.005 401.365 -127.675 ;
        RECT 401.035 -129.365 401.365 -129.035 ;
        RECT 401.035 -130.725 401.365 -130.395 ;
        RECT 401.035 -132.085 401.365 -131.755 ;
        RECT 401.035 -133.445 401.365 -133.115 ;
        RECT 401.035 -134.805 401.365 -134.475 ;
        RECT 401.035 -136.165 401.365 -135.835 ;
        RECT 401.035 -137.525 401.365 -137.195 ;
        RECT 401.035 -138.885 401.365 -138.555 ;
        RECT 401.035 -140.245 401.365 -139.915 ;
        RECT 401.035 -141.605 401.365 -141.275 ;
        RECT 401.035 -142.965 401.365 -142.635 ;
        RECT 401.035 -144.325 401.365 -143.995 ;
        RECT 401.035 -145.685 401.365 -145.355 ;
        RECT 401.035 -147.045 401.365 -146.715 ;
        RECT 401.035 -148.405 401.365 -148.075 ;
        RECT 401.035 -149.765 401.365 -149.435 ;
        RECT 401.035 -151.125 401.365 -150.795 ;
        RECT 401.035 -152.485 401.365 -152.155 ;
        RECT 401.035 -153.845 401.365 -153.515 ;
        RECT 401.035 -155.205 401.365 -154.875 ;
        RECT 401.035 -156.565 401.365 -156.235 ;
        RECT 401.035 -157.925 401.365 -157.595 ;
        RECT 401.035 -159.285 401.365 -158.955 ;
        RECT 401.035 -160.645 401.365 -160.315 ;
        RECT 401.035 -162.005 401.365 -161.675 ;
        RECT 401.035 -163.365 401.365 -163.035 ;
        RECT 401.035 -164.725 401.365 -164.395 ;
        RECT 401.035 -166.085 401.365 -165.755 ;
        RECT 401.035 -167.445 401.365 -167.115 ;
        RECT 401.035 -168.805 401.365 -168.475 ;
        RECT 401.035 -170.165 401.365 -169.835 ;
        RECT 401.035 -171.525 401.365 -171.195 ;
        RECT 401.035 -172.885 401.365 -172.555 ;
        RECT 401.035 -174.245 401.365 -173.915 ;
        RECT 401.035 -175.605 401.365 -175.275 ;
        RECT 401.035 -176.965 401.365 -176.635 ;
        RECT 401.035 -178.325 401.365 -177.995 ;
        RECT 401.035 -180.57 401.365 -179.44 ;
        RECT 401.04 -180.685 401.36 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 402.395 241.32 402.725 242.45 ;
        RECT 402.395 239.195 402.725 239.525 ;
        RECT 402.395 237.835 402.725 238.165 ;
        RECT 402.395 -1.525 402.725 -1.195 ;
        RECT 402.395 -2.885 402.725 -2.555 ;
        RECT 402.395 -4.245 402.725 -3.915 ;
        RECT 402.395 -5.605 402.725 -5.275 ;
        RECT 402.395 -6.965 402.725 -6.635 ;
        RECT 402.395 -8.325 402.725 -7.995 ;
        RECT 402.395 -9.685 402.725 -9.355 ;
        RECT 402.395 -11.045 402.725 -10.715 ;
        RECT 402.395 -12.405 402.725 -12.075 ;
        RECT 402.395 -13.765 402.725 -13.435 ;
        RECT 402.395 -15.125 402.725 -14.795 ;
        RECT 402.395 -16.485 402.725 -16.155 ;
        RECT 402.395 -17.845 402.725 -17.515 ;
        RECT 402.395 -19.205 402.725 -18.875 ;
        RECT 402.395 -20.565 402.725 -20.235 ;
        RECT 402.395 -21.925 402.725 -21.595 ;
        RECT 402.395 -23.285 402.725 -22.955 ;
        RECT 402.395 -24.645 402.725 -24.315 ;
        RECT 402.395 -26.005 402.725 -25.675 ;
        RECT 402.395 -27.365 402.725 -27.035 ;
        RECT 402.395 -28.725 402.725 -28.395 ;
        RECT 402.395 -30.085 402.725 -29.755 ;
        RECT 402.395 -31.445 402.725 -31.115 ;
        RECT 402.395 -32.805 402.725 -32.475 ;
        RECT 402.395 -34.165 402.725 -33.835 ;
        RECT 402.395 -35.525 402.725 -35.195 ;
        RECT 402.395 -36.885 402.725 -36.555 ;
        RECT 402.395 -38.245 402.725 -37.915 ;
        RECT 402.395 -39.605 402.725 -39.275 ;
        RECT 402.395 -40.965 402.725 -40.635 ;
        RECT 402.395 -42.325 402.725 -41.995 ;
        RECT 402.395 -43.685 402.725 -43.355 ;
        RECT 402.395 -45.045 402.725 -44.715 ;
        RECT 402.395 -46.405 402.725 -46.075 ;
        RECT 402.395 -47.765 402.725 -47.435 ;
        RECT 402.395 -49.125 402.725 -48.795 ;
        RECT 402.395 -50.485 402.725 -50.155 ;
        RECT 402.395 -51.845 402.725 -51.515 ;
        RECT 402.395 -53.205 402.725 -52.875 ;
        RECT 402.395 -54.565 402.725 -54.235 ;
        RECT 402.395 -55.925 402.725 -55.595 ;
        RECT 402.395 -57.285 402.725 -56.955 ;
        RECT 402.395 -58.645 402.725 -58.315 ;
        RECT 402.395 -60.005 402.725 -59.675 ;
        RECT 402.395 -61.365 402.725 -61.035 ;
        RECT 402.395 -62.725 402.725 -62.395 ;
        RECT 402.395 -64.085 402.725 -63.755 ;
        RECT 402.395 -65.445 402.725 -65.115 ;
        RECT 402.395 -66.805 402.725 -66.475 ;
        RECT 402.395 -68.165 402.725 -67.835 ;
        RECT 402.395 -69.525 402.725 -69.195 ;
        RECT 402.395 -70.885 402.725 -70.555 ;
        RECT 402.395 -72.245 402.725 -71.915 ;
        RECT 402.395 -73.605 402.725 -73.275 ;
        RECT 402.395 -74.965 402.725 -74.635 ;
        RECT 402.395 -76.325 402.725 -75.995 ;
        RECT 402.395 -77.685 402.725 -77.355 ;
        RECT 402.395 -79.045 402.725 -78.715 ;
        RECT 402.395 -80.405 402.725 -80.075 ;
        RECT 402.395 -81.765 402.725 -81.435 ;
        RECT 402.395 -83.125 402.725 -82.795 ;
        RECT 402.395 -84.485 402.725 -84.155 ;
        RECT 402.395 -85.845 402.725 -85.515 ;
        RECT 402.395 -87.205 402.725 -86.875 ;
        RECT 402.395 -88.565 402.725 -88.235 ;
        RECT 402.395 -89.925 402.725 -89.595 ;
        RECT 402.395 -91.285 402.725 -90.955 ;
        RECT 402.395 -92.645 402.725 -92.315 ;
        RECT 402.395 -94.005 402.725 -93.675 ;
        RECT 402.395 -95.365 402.725 -95.035 ;
        RECT 402.395 -96.725 402.725 -96.395 ;
        RECT 402.395 -98.085 402.725 -97.755 ;
        RECT 402.395 -99.445 402.725 -99.115 ;
        RECT 402.395 -100.805 402.725 -100.475 ;
        RECT 402.395 -102.165 402.725 -101.835 ;
        RECT 402.395 -103.525 402.725 -103.195 ;
        RECT 402.395 -104.885 402.725 -104.555 ;
        RECT 402.395 -106.245 402.725 -105.915 ;
        RECT 402.395 -107.605 402.725 -107.275 ;
        RECT 402.395 -108.965 402.725 -108.635 ;
        RECT 402.395 -110.325 402.725 -109.995 ;
        RECT 402.395 -111.685 402.725 -111.355 ;
        RECT 402.395 -113.045 402.725 -112.715 ;
        RECT 402.395 -114.405 402.725 -114.075 ;
        RECT 402.395 -115.765 402.725 -115.435 ;
        RECT 402.395 -117.125 402.725 -116.795 ;
        RECT 402.395 -118.485 402.725 -118.155 ;
        RECT 402.395 -119.845 402.725 -119.515 ;
        RECT 402.395 -121.205 402.725 -120.875 ;
        RECT 402.395 -122.565 402.725 -122.235 ;
        RECT 402.395 -123.925 402.725 -123.595 ;
        RECT 402.395 -125.285 402.725 -124.955 ;
        RECT 402.395 -126.645 402.725 -126.315 ;
        RECT 402.395 -128.005 402.725 -127.675 ;
        RECT 402.395 -129.365 402.725 -129.035 ;
        RECT 402.395 -130.725 402.725 -130.395 ;
        RECT 402.395 -132.085 402.725 -131.755 ;
        RECT 402.395 -133.445 402.725 -133.115 ;
        RECT 402.395 -134.805 402.725 -134.475 ;
        RECT 402.395 -136.165 402.725 -135.835 ;
        RECT 402.395 -137.525 402.725 -137.195 ;
        RECT 402.395 -138.885 402.725 -138.555 ;
        RECT 402.395 -140.245 402.725 -139.915 ;
        RECT 402.395 -141.605 402.725 -141.275 ;
        RECT 402.395 -142.965 402.725 -142.635 ;
        RECT 402.395 -144.325 402.725 -143.995 ;
        RECT 402.395 -145.685 402.725 -145.355 ;
        RECT 402.395 -147.045 402.725 -146.715 ;
        RECT 402.395 -148.405 402.725 -148.075 ;
        RECT 402.395 -149.765 402.725 -149.435 ;
        RECT 402.395 -151.125 402.725 -150.795 ;
        RECT 402.395 -152.485 402.725 -152.155 ;
        RECT 402.395 -153.845 402.725 -153.515 ;
        RECT 402.395 -155.205 402.725 -154.875 ;
        RECT 402.395 -156.565 402.725 -156.235 ;
        RECT 402.395 -157.925 402.725 -157.595 ;
        RECT 402.395 -159.285 402.725 -158.955 ;
        RECT 402.395 -160.645 402.725 -160.315 ;
        RECT 402.395 -162.005 402.725 -161.675 ;
        RECT 402.395 -163.365 402.725 -163.035 ;
        RECT 402.395 -164.725 402.725 -164.395 ;
        RECT 402.395 -166.085 402.725 -165.755 ;
        RECT 402.395 -167.445 402.725 -167.115 ;
        RECT 402.395 -168.805 402.725 -168.475 ;
        RECT 402.395 -170.165 402.725 -169.835 ;
        RECT 402.395 -171.525 402.725 -171.195 ;
        RECT 402.395 -172.885 402.725 -172.555 ;
        RECT 402.395 -174.245 402.725 -173.915 ;
        RECT 402.395 -175.605 402.725 -175.275 ;
        RECT 402.395 -176.965 402.725 -176.635 ;
        RECT 402.395 -178.325 402.725 -177.995 ;
        RECT 402.395 -180.57 402.725 -179.44 ;
        RECT 402.4 -180.685 402.72 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 369.31 -94.075 369.64 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 369.755 241.32 370.085 242.45 ;
        RECT 369.755 239.195 370.085 239.525 ;
        RECT 369.755 237.835 370.085 238.165 ;
        RECT 369.76 237.16 370.08 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 371.115 241.32 371.445 242.45 ;
        RECT 371.115 239.195 371.445 239.525 ;
        RECT 371.115 237.835 371.445 238.165 ;
        RECT 371.12 237.16 371.44 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 371.115 -1.525 371.445 -1.195 ;
        RECT 371.115 -2.885 371.445 -2.555 ;
        RECT 371.12 -3.56 371.44 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 372.475 241.32 372.805 242.45 ;
        RECT 372.475 239.195 372.805 239.525 ;
        RECT 372.475 237.835 372.805 238.165 ;
        RECT 372.48 237.16 372.8 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 372.475 -1.525 372.805 -1.195 ;
        RECT 372.475 -2.885 372.805 -2.555 ;
        RECT 372.48 -3.56 372.8 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 372.475 -91.285 372.805 -90.955 ;
        RECT 372.475 -92.645 372.805 -92.315 ;
        RECT 372.475 -94.005 372.805 -93.675 ;
        RECT 372.475 -95.365 372.805 -95.035 ;
        RECT 372.475 -96.725 372.805 -96.395 ;
        RECT 372.475 -98.085 372.805 -97.755 ;
        RECT 372.475 -99.445 372.805 -99.115 ;
        RECT 372.475 -100.805 372.805 -100.475 ;
        RECT 372.475 -102.165 372.805 -101.835 ;
        RECT 372.475 -103.525 372.805 -103.195 ;
        RECT 372.475 -104.885 372.805 -104.555 ;
        RECT 372.475 -106.245 372.805 -105.915 ;
        RECT 372.475 -107.605 372.805 -107.275 ;
        RECT 372.475 -108.965 372.805 -108.635 ;
        RECT 372.475 -110.325 372.805 -109.995 ;
        RECT 372.475 -111.685 372.805 -111.355 ;
        RECT 372.475 -113.045 372.805 -112.715 ;
        RECT 372.475 -114.405 372.805 -114.075 ;
        RECT 372.475 -115.765 372.805 -115.435 ;
        RECT 372.475 -117.125 372.805 -116.795 ;
        RECT 372.475 -118.485 372.805 -118.155 ;
        RECT 372.475 -119.845 372.805 -119.515 ;
        RECT 372.475 -121.205 372.805 -120.875 ;
        RECT 372.475 -122.565 372.805 -122.235 ;
        RECT 372.475 -123.925 372.805 -123.595 ;
        RECT 372.475 -125.285 372.805 -124.955 ;
        RECT 372.475 -126.645 372.805 -126.315 ;
        RECT 372.475 -128.005 372.805 -127.675 ;
        RECT 372.475 -129.365 372.805 -129.035 ;
        RECT 372.475 -130.725 372.805 -130.395 ;
        RECT 372.475 -132.085 372.805 -131.755 ;
        RECT 372.475 -133.445 372.805 -133.115 ;
        RECT 372.475 -134.805 372.805 -134.475 ;
        RECT 372.475 -136.165 372.805 -135.835 ;
        RECT 372.475 -137.525 372.805 -137.195 ;
        RECT 372.475 -138.885 372.805 -138.555 ;
        RECT 372.475 -140.245 372.805 -139.915 ;
        RECT 372.475 -141.605 372.805 -141.275 ;
        RECT 372.475 -142.965 372.805 -142.635 ;
        RECT 372.475 -144.325 372.805 -143.995 ;
        RECT 372.475 -145.685 372.805 -145.355 ;
        RECT 372.475 -147.045 372.805 -146.715 ;
        RECT 372.475 -148.405 372.805 -148.075 ;
        RECT 372.475 -149.765 372.805 -149.435 ;
        RECT 372.475 -151.125 372.805 -150.795 ;
        RECT 372.475 -152.485 372.805 -152.155 ;
        RECT 372.475 -153.845 372.805 -153.515 ;
        RECT 372.475 -155.205 372.805 -154.875 ;
        RECT 372.475 -156.565 372.805 -156.235 ;
        RECT 372.475 -157.925 372.805 -157.595 ;
        RECT 372.475 -159.285 372.805 -158.955 ;
        RECT 372.475 -160.645 372.805 -160.315 ;
        RECT 372.475 -162.005 372.805 -161.675 ;
        RECT 372.475 -163.365 372.805 -163.035 ;
        RECT 372.475 -164.725 372.805 -164.395 ;
        RECT 372.475 -166.085 372.805 -165.755 ;
        RECT 372.475 -167.445 372.805 -167.115 ;
        RECT 372.475 -168.805 372.805 -168.475 ;
        RECT 372.475 -170.165 372.805 -169.835 ;
        RECT 372.475 -171.525 372.805 -171.195 ;
        RECT 372.475 -172.885 372.805 -172.555 ;
        RECT 372.475 -174.245 372.805 -173.915 ;
        RECT 372.475 -175.605 372.805 -175.275 ;
        RECT 372.475 -176.965 372.805 -176.635 ;
        RECT 372.475 -178.325 372.805 -177.995 ;
        RECT 372.475 -180.57 372.805 -179.44 ;
        RECT 372.48 -180.685 372.8 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 373.835 241.32 374.165 242.45 ;
        RECT 373.835 239.195 374.165 239.525 ;
        RECT 373.835 237.835 374.165 238.165 ;
        RECT 373.84 237.16 374.16 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 373.835 -1.525 374.165 -1.195 ;
        RECT 373.835 -2.885 374.165 -2.555 ;
        RECT 373.84 -3.56 374.16 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 373.835 -91.285 374.165 -90.955 ;
        RECT 373.835 -92.645 374.165 -92.315 ;
        RECT 373.835 -94.005 374.165 -93.675 ;
        RECT 373.835 -95.365 374.165 -95.035 ;
        RECT 373.835 -96.725 374.165 -96.395 ;
        RECT 373.835 -98.085 374.165 -97.755 ;
        RECT 373.835 -99.445 374.165 -99.115 ;
        RECT 373.835 -100.805 374.165 -100.475 ;
        RECT 373.835 -102.165 374.165 -101.835 ;
        RECT 373.835 -103.525 374.165 -103.195 ;
        RECT 373.835 -104.885 374.165 -104.555 ;
        RECT 373.835 -106.245 374.165 -105.915 ;
        RECT 373.835 -107.605 374.165 -107.275 ;
        RECT 373.835 -108.965 374.165 -108.635 ;
        RECT 373.835 -110.325 374.165 -109.995 ;
        RECT 373.835 -111.685 374.165 -111.355 ;
        RECT 373.835 -113.045 374.165 -112.715 ;
        RECT 373.835 -114.405 374.165 -114.075 ;
        RECT 373.835 -115.765 374.165 -115.435 ;
        RECT 373.835 -117.125 374.165 -116.795 ;
        RECT 373.835 -118.485 374.165 -118.155 ;
        RECT 373.835 -119.845 374.165 -119.515 ;
        RECT 373.835 -121.205 374.165 -120.875 ;
        RECT 373.835 -122.565 374.165 -122.235 ;
        RECT 373.835 -123.925 374.165 -123.595 ;
        RECT 373.835 -125.285 374.165 -124.955 ;
        RECT 373.835 -126.645 374.165 -126.315 ;
        RECT 373.835 -128.005 374.165 -127.675 ;
        RECT 373.835 -129.365 374.165 -129.035 ;
        RECT 373.835 -130.725 374.165 -130.395 ;
        RECT 373.835 -132.085 374.165 -131.755 ;
        RECT 373.835 -133.445 374.165 -133.115 ;
        RECT 373.835 -134.805 374.165 -134.475 ;
        RECT 373.835 -136.165 374.165 -135.835 ;
        RECT 373.835 -137.525 374.165 -137.195 ;
        RECT 373.835 -138.885 374.165 -138.555 ;
        RECT 373.835 -140.245 374.165 -139.915 ;
        RECT 373.835 -141.605 374.165 -141.275 ;
        RECT 373.835 -142.965 374.165 -142.635 ;
        RECT 373.835 -144.325 374.165 -143.995 ;
        RECT 373.835 -145.685 374.165 -145.355 ;
        RECT 373.835 -147.045 374.165 -146.715 ;
        RECT 373.835 -148.405 374.165 -148.075 ;
        RECT 373.835 -149.765 374.165 -149.435 ;
        RECT 373.835 -151.125 374.165 -150.795 ;
        RECT 373.835 -152.485 374.165 -152.155 ;
        RECT 373.835 -153.845 374.165 -153.515 ;
        RECT 373.835 -155.205 374.165 -154.875 ;
        RECT 373.835 -156.565 374.165 -156.235 ;
        RECT 373.835 -157.925 374.165 -157.595 ;
        RECT 373.835 -159.285 374.165 -158.955 ;
        RECT 373.835 -160.645 374.165 -160.315 ;
        RECT 373.835 -162.005 374.165 -161.675 ;
        RECT 373.835 -163.365 374.165 -163.035 ;
        RECT 373.835 -164.725 374.165 -164.395 ;
        RECT 373.835 -166.085 374.165 -165.755 ;
        RECT 373.835 -167.445 374.165 -167.115 ;
        RECT 373.835 -168.805 374.165 -168.475 ;
        RECT 373.835 -170.165 374.165 -169.835 ;
        RECT 373.835 -171.525 374.165 -171.195 ;
        RECT 373.835 -172.885 374.165 -172.555 ;
        RECT 373.835 -174.245 374.165 -173.915 ;
        RECT 373.835 -175.605 374.165 -175.275 ;
        RECT 373.835 -176.965 374.165 -176.635 ;
        RECT 373.835 -178.325 374.165 -177.995 ;
        RECT 373.835 -180.57 374.165 -179.44 ;
        RECT 373.84 -180.685 374.16 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 375.195 241.32 375.525 242.45 ;
        RECT 375.195 239.195 375.525 239.525 ;
        RECT 375.195 237.835 375.525 238.165 ;
        RECT 375.2 237.16 375.52 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 375.195 -95.365 375.525 -95.035 ;
        RECT 375.195 -96.725 375.525 -96.395 ;
        RECT 375.195 -98.085 375.525 -97.755 ;
        RECT 375.195 -99.445 375.525 -99.115 ;
        RECT 375.195 -100.805 375.525 -100.475 ;
        RECT 375.195 -102.165 375.525 -101.835 ;
        RECT 375.195 -103.525 375.525 -103.195 ;
        RECT 375.195 -104.885 375.525 -104.555 ;
        RECT 375.195 -106.245 375.525 -105.915 ;
        RECT 375.195 -107.605 375.525 -107.275 ;
        RECT 375.195 -108.965 375.525 -108.635 ;
        RECT 375.195 -110.325 375.525 -109.995 ;
        RECT 375.195 -111.685 375.525 -111.355 ;
        RECT 375.195 -113.045 375.525 -112.715 ;
        RECT 375.195 -114.405 375.525 -114.075 ;
        RECT 375.195 -115.765 375.525 -115.435 ;
        RECT 375.195 -117.125 375.525 -116.795 ;
        RECT 375.195 -118.485 375.525 -118.155 ;
        RECT 375.195 -119.845 375.525 -119.515 ;
        RECT 375.195 -121.205 375.525 -120.875 ;
        RECT 375.195 -122.565 375.525 -122.235 ;
        RECT 375.195 -123.925 375.525 -123.595 ;
        RECT 375.195 -125.285 375.525 -124.955 ;
        RECT 375.195 -126.645 375.525 -126.315 ;
        RECT 375.195 -128.005 375.525 -127.675 ;
        RECT 375.195 -129.365 375.525 -129.035 ;
        RECT 375.195 -130.725 375.525 -130.395 ;
        RECT 375.195 -132.085 375.525 -131.755 ;
        RECT 375.195 -133.445 375.525 -133.115 ;
        RECT 375.195 -134.805 375.525 -134.475 ;
        RECT 375.195 -136.165 375.525 -135.835 ;
        RECT 375.195 -137.525 375.525 -137.195 ;
        RECT 375.195 -138.885 375.525 -138.555 ;
        RECT 375.195 -140.245 375.525 -139.915 ;
        RECT 375.195 -141.605 375.525 -141.275 ;
        RECT 375.195 -142.965 375.525 -142.635 ;
        RECT 375.195 -144.325 375.525 -143.995 ;
        RECT 375.195 -145.685 375.525 -145.355 ;
        RECT 375.195 -147.045 375.525 -146.715 ;
        RECT 375.195 -148.405 375.525 -148.075 ;
        RECT 375.195 -149.765 375.525 -149.435 ;
        RECT 375.195 -151.125 375.525 -150.795 ;
        RECT 375.195 -152.485 375.525 -152.155 ;
        RECT 375.195 -153.845 375.525 -153.515 ;
        RECT 375.195 -155.205 375.525 -154.875 ;
        RECT 375.195 -156.565 375.525 -156.235 ;
        RECT 375.195 -157.925 375.525 -157.595 ;
        RECT 375.195 -159.285 375.525 -158.955 ;
        RECT 375.195 -160.645 375.525 -160.315 ;
        RECT 375.195 -162.005 375.525 -161.675 ;
        RECT 375.195 -163.365 375.525 -163.035 ;
        RECT 375.195 -164.725 375.525 -164.395 ;
        RECT 375.195 -166.085 375.525 -165.755 ;
        RECT 375.195 -167.445 375.525 -167.115 ;
        RECT 375.195 -168.805 375.525 -168.475 ;
        RECT 375.195 -170.165 375.525 -169.835 ;
        RECT 375.195 -171.525 375.525 -171.195 ;
        RECT 375.195 -172.885 375.525 -172.555 ;
        RECT 375.195 -174.245 375.525 -173.915 ;
        RECT 375.195 -175.605 375.525 -175.275 ;
        RECT 375.195 -176.965 375.525 -176.635 ;
        RECT 375.195 -178.325 375.525 -177.995 ;
        RECT 375.195 -180.57 375.525 -179.44 ;
        RECT 375.2 -180.685 375.52 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 375.41 -94.075 375.74 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 376.555 241.32 376.885 242.45 ;
        RECT 376.555 239.195 376.885 239.525 ;
        RECT 376.555 237.835 376.885 238.165 ;
        RECT 376.56 237.16 376.88 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 376.555 -1.525 376.885 -1.195 ;
        RECT 376.555 -2.885 376.885 -2.555 ;
        RECT 376.56 -3.56 376.88 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 377.915 241.32 378.245 242.45 ;
        RECT 377.915 239.195 378.245 239.525 ;
        RECT 377.915 237.835 378.245 238.165 ;
        RECT 377.92 237.16 378.24 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 377.915 -1.525 378.245 -1.195 ;
        RECT 377.915 -2.885 378.245 -2.555 ;
        RECT 377.92 -3.56 378.24 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 379.275 241.32 379.605 242.45 ;
        RECT 379.275 239.195 379.605 239.525 ;
        RECT 379.275 237.835 379.605 238.165 ;
        RECT 379.28 237.16 379.6 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 379.275 -1.525 379.605 -1.195 ;
        RECT 379.275 -2.885 379.605 -2.555 ;
        RECT 379.28 -3.56 379.6 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 379.275 -91.285 379.605 -90.955 ;
        RECT 379.275 -92.645 379.605 -92.315 ;
        RECT 379.275 -94.005 379.605 -93.675 ;
        RECT 379.275 -95.365 379.605 -95.035 ;
        RECT 379.275 -96.725 379.605 -96.395 ;
        RECT 379.275 -98.085 379.605 -97.755 ;
        RECT 379.275 -99.445 379.605 -99.115 ;
        RECT 379.275 -100.805 379.605 -100.475 ;
        RECT 379.275 -102.165 379.605 -101.835 ;
        RECT 379.275 -103.525 379.605 -103.195 ;
        RECT 379.275 -104.885 379.605 -104.555 ;
        RECT 379.275 -106.245 379.605 -105.915 ;
        RECT 379.275 -107.605 379.605 -107.275 ;
        RECT 379.275 -108.965 379.605 -108.635 ;
        RECT 379.275 -110.325 379.605 -109.995 ;
        RECT 379.275 -111.685 379.605 -111.355 ;
        RECT 379.275 -113.045 379.605 -112.715 ;
        RECT 379.275 -114.405 379.605 -114.075 ;
        RECT 379.275 -115.765 379.605 -115.435 ;
        RECT 379.275 -117.125 379.605 -116.795 ;
        RECT 379.275 -118.485 379.605 -118.155 ;
        RECT 379.275 -119.845 379.605 -119.515 ;
        RECT 379.275 -121.205 379.605 -120.875 ;
        RECT 379.275 -122.565 379.605 -122.235 ;
        RECT 379.275 -123.925 379.605 -123.595 ;
        RECT 379.275 -125.285 379.605 -124.955 ;
        RECT 379.275 -126.645 379.605 -126.315 ;
        RECT 379.275 -128.005 379.605 -127.675 ;
        RECT 379.275 -129.365 379.605 -129.035 ;
        RECT 379.275 -130.725 379.605 -130.395 ;
        RECT 379.275 -132.085 379.605 -131.755 ;
        RECT 379.275 -133.445 379.605 -133.115 ;
        RECT 379.275 -134.805 379.605 -134.475 ;
        RECT 379.275 -136.165 379.605 -135.835 ;
        RECT 379.275 -137.525 379.605 -137.195 ;
        RECT 379.275 -138.885 379.605 -138.555 ;
        RECT 379.275 -140.245 379.605 -139.915 ;
        RECT 379.275 -141.605 379.605 -141.275 ;
        RECT 379.275 -142.965 379.605 -142.635 ;
        RECT 379.275 -144.325 379.605 -143.995 ;
        RECT 379.275 -145.685 379.605 -145.355 ;
        RECT 379.275 -147.045 379.605 -146.715 ;
        RECT 379.275 -148.405 379.605 -148.075 ;
        RECT 379.275 -149.765 379.605 -149.435 ;
        RECT 379.275 -151.125 379.605 -150.795 ;
        RECT 379.275 -152.485 379.605 -152.155 ;
        RECT 379.275 -153.845 379.605 -153.515 ;
        RECT 379.275 -155.205 379.605 -154.875 ;
        RECT 379.275 -156.565 379.605 -156.235 ;
        RECT 379.275 -157.925 379.605 -157.595 ;
        RECT 379.275 -159.285 379.605 -158.955 ;
        RECT 379.275 -160.645 379.605 -160.315 ;
        RECT 379.275 -162.005 379.605 -161.675 ;
        RECT 379.275 -163.365 379.605 -163.035 ;
        RECT 379.275 -164.725 379.605 -164.395 ;
        RECT 379.275 -166.085 379.605 -165.755 ;
        RECT 379.275 -167.445 379.605 -167.115 ;
        RECT 379.275 -168.805 379.605 -168.475 ;
        RECT 379.275 -170.165 379.605 -169.835 ;
        RECT 379.275 -171.525 379.605 -171.195 ;
        RECT 379.275 -172.885 379.605 -172.555 ;
        RECT 379.275 -174.245 379.605 -173.915 ;
        RECT 379.275 -175.605 379.605 -175.275 ;
        RECT 379.275 -176.965 379.605 -176.635 ;
        RECT 379.275 -178.325 379.605 -177.995 ;
        RECT 379.275 -180.57 379.605 -179.44 ;
        RECT 379.28 -180.685 379.6 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 380.635 241.32 380.965 242.45 ;
        RECT 380.635 239.195 380.965 239.525 ;
        RECT 380.635 237.835 380.965 238.165 ;
        RECT 380.64 237.16 380.96 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 380.635 -95.365 380.965 -95.035 ;
        RECT 380.635 -96.725 380.965 -96.395 ;
        RECT 380.635 -98.085 380.965 -97.755 ;
        RECT 380.635 -99.445 380.965 -99.115 ;
        RECT 380.635 -100.805 380.965 -100.475 ;
        RECT 380.635 -102.165 380.965 -101.835 ;
        RECT 380.635 -103.525 380.965 -103.195 ;
        RECT 380.635 -104.885 380.965 -104.555 ;
        RECT 380.635 -106.245 380.965 -105.915 ;
        RECT 380.635 -107.605 380.965 -107.275 ;
        RECT 380.635 -108.965 380.965 -108.635 ;
        RECT 380.635 -110.325 380.965 -109.995 ;
        RECT 380.635 -111.685 380.965 -111.355 ;
        RECT 380.635 -113.045 380.965 -112.715 ;
        RECT 380.635 -114.405 380.965 -114.075 ;
        RECT 380.635 -115.765 380.965 -115.435 ;
        RECT 380.635 -117.125 380.965 -116.795 ;
        RECT 380.635 -118.485 380.965 -118.155 ;
        RECT 380.635 -119.845 380.965 -119.515 ;
        RECT 380.635 -121.205 380.965 -120.875 ;
        RECT 380.635 -122.565 380.965 -122.235 ;
        RECT 380.635 -123.925 380.965 -123.595 ;
        RECT 380.635 -125.285 380.965 -124.955 ;
        RECT 380.635 -126.645 380.965 -126.315 ;
        RECT 380.635 -128.005 380.965 -127.675 ;
        RECT 380.635 -129.365 380.965 -129.035 ;
        RECT 380.635 -130.725 380.965 -130.395 ;
        RECT 380.635 -132.085 380.965 -131.755 ;
        RECT 380.635 -133.445 380.965 -133.115 ;
        RECT 380.635 -134.805 380.965 -134.475 ;
        RECT 380.635 -136.165 380.965 -135.835 ;
        RECT 380.635 -137.525 380.965 -137.195 ;
        RECT 380.635 -138.885 380.965 -138.555 ;
        RECT 380.635 -140.245 380.965 -139.915 ;
        RECT 380.635 -141.605 380.965 -141.275 ;
        RECT 380.635 -142.965 380.965 -142.635 ;
        RECT 380.635 -144.325 380.965 -143.995 ;
        RECT 380.635 -145.685 380.965 -145.355 ;
        RECT 380.635 -147.045 380.965 -146.715 ;
        RECT 380.635 -148.405 380.965 -148.075 ;
        RECT 380.635 -149.765 380.965 -149.435 ;
        RECT 380.635 -151.125 380.965 -150.795 ;
        RECT 380.635 -152.485 380.965 -152.155 ;
        RECT 380.635 -153.845 380.965 -153.515 ;
        RECT 380.635 -155.205 380.965 -154.875 ;
        RECT 380.635 -156.565 380.965 -156.235 ;
        RECT 380.635 -157.925 380.965 -157.595 ;
        RECT 380.635 -159.285 380.965 -158.955 ;
        RECT 380.635 -160.645 380.965 -160.315 ;
        RECT 380.635 -162.005 380.965 -161.675 ;
        RECT 380.635 -163.365 380.965 -163.035 ;
        RECT 380.635 -164.725 380.965 -164.395 ;
        RECT 380.635 -166.085 380.965 -165.755 ;
        RECT 380.635 -167.445 380.965 -167.115 ;
        RECT 380.635 -168.805 380.965 -168.475 ;
        RECT 380.635 -170.165 380.965 -169.835 ;
        RECT 380.635 -171.525 380.965 -171.195 ;
        RECT 380.635 -172.885 380.965 -172.555 ;
        RECT 380.635 -174.245 380.965 -173.915 ;
        RECT 380.635 -175.605 380.965 -175.275 ;
        RECT 380.635 -176.965 380.965 -176.635 ;
        RECT 380.635 -178.325 380.965 -177.995 ;
        RECT 380.635 -180.57 380.965 -179.44 ;
        RECT 380.64 -180.685 380.96 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 381.51 -94.075 381.84 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 381.995 241.32 382.325 242.45 ;
        RECT 381.995 239.195 382.325 239.525 ;
        RECT 381.995 237.835 382.325 238.165 ;
        RECT 382 237.16 382.32 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 383.355 241.32 383.685 242.45 ;
        RECT 383.355 239.195 383.685 239.525 ;
        RECT 383.355 237.835 383.685 238.165 ;
        RECT 383.36 237.16 383.68 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 383.355 -1.525 383.685 -1.195 ;
        RECT 383.355 -2.885 383.685 -2.555 ;
        RECT 383.36 -3.56 383.68 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 384.715 241.32 385.045 242.45 ;
        RECT 384.715 239.195 385.045 239.525 ;
        RECT 384.715 237.835 385.045 238.165 ;
        RECT 384.72 237.16 385.04 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 384.715 -1.525 385.045 -1.195 ;
        RECT 384.715 -2.885 385.045 -2.555 ;
        RECT 384.72 -3.56 385.04 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 384.715 -91.285 385.045 -90.955 ;
        RECT 384.715 -92.645 385.045 -92.315 ;
        RECT 384.715 -94.005 385.045 -93.675 ;
        RECT 384.715 -95.365 385.045 -95.035 ;
        RECT 384.715 -96.725 385.045 -96.395 ;
        RECT 384.715 -98.085 385.045 -97.755 ;
        RECT 384.715 -99.445 385.045 -99.115 ;
        RECT 384.715 -100.805 385.045 -100.475 ;
        RECT 384.715 -102.165 385.045 -101.835 ;
        RECT 384.715 -103.525 385.045 -103.195 ;
        RECT 384.715 -104.885 385.045 -104.555 ;
        RECT 384.715 -106.245 385.045 -105.915 ;
        RECT 384.715 -107.605 385.045 -107.275 ;
        RECT 384.715 -108.965 385.045 -108.635 ;
        RECT 384.715 -110.325 385.045 -109.995 ;
        RECT 384.715 -111.685 385.045 -111.355 ;
        RECT 384.715 -113.045 385.045 -112.715 ;
        RECT 384.715 -114.405 385.045 -114.075 ;
        RECT 384.715 -115.765 385.045 -115.435 ;
        RECT 384.715 -117.125 385.045 -116.795 ;
        RECT 384.715 -118.485 385.045 -118.155 ;
        RECT 384.715 -119.845 385.045 -119.515 ;
        RECT 384.715 -121.205 385.045 -120.875 ;
        RECT 384.715 -122.565 385.045 -122.235 ;
        RECT 384.715 -123.925 385.045 -123.595 ;
        RECT 384.715 -125.285 385.045 -124.955 ;
        RECT 384.715 -126.645 385.045 -126.315 ;
        RECT 384.715 -128.005 385.045 -127.675 ;
        RECT 384.715 -129.365 385.045 -129.035 ;
        RECT 384.715 -130.725 385.045 -130.395 ;
        RECT 384.715 -132.085 385.045 -131.755 ;
        RECT 384.715 -133.445 385.045 -133.115 ;
        RECT 384.715 -134.805 385.045 -134.475 ;
        RECT 384.715 -136.165 385.045 -135.835 ;
        RECT 384.715 -137.525 385.045 -137.195 ;
        RECT 384.715 -138.885 385.045 -138.555 ;
        RECT 384.715 -140.245 385.045 -139.915 ;
        RECT 384.715 -141.605 385.045 -141.275 ;
        RECT 384.715 -142.965 385.045 -142.635 ;
        RECT 384.715 -144.325 385.045 -143.995 ;
        RECT 384.715 -145.685 385.045 -145.355 ;
        RECT 384.715 -147.045 385.045 -146.715 ;
        RECT 384.715 -148.405 385.045 -148.075 ;
        RECT 384.715 -149.765 385.045 -149.435 ;
        RECT 384.715 -151.125 385.045 -150.795 ;
        RECT 384.715 -152.485 385.045 -152.155 ;
        RECT 384.715 -153.845 385.045 -153.515 ;
        RECT 384.715 -155.205 385.045 -154.875 ;
        RECT 384.715 -156.565 385.045 -156.235 ;
        RECT 384.715 -157.925 385.045 -157.595 ;
        RECT 384.715 -159.285 385.045 -158.955 ;
        RECT 384.715 -160.645 385.045 -160.315 ;
        RECT 384.715 -162.005 385.045 -161.675 ;
        RECT 384.715 -163.365 385.045 -163.035 ;
        RECT 384.715 -164.725 385.045 -164.395 ;
        RECT 384.715 -166.085 385.045 -165.755 ;
        RECT 384.715 -167.445 385.045 -167.115 ;
        RECT 384.715 -168.805 385.045 -168.475 ;
        RECT 384.715 -170.165 385.045 -169.835 ;
        RECT 384.715 -171.525 385.045 -171.195 ;
        RECT 384.715 -172.885 385.045 -172.555 ;
        RECT 384.715 -174.245 385.045 -173.915 ;
        RECT 384.715 -175.605 385.045 -175.275 ;
        RECT 384.715 -176.965 385.045 -176.635 ;
        RECT 384.715 -178.325 385.045 -177.995 ;
        RECT 384.715 -180.57 385.045 -179.44 ;
        RECT 384.72 -180.685 385.04 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 386.075 241.32 386.405 242.45 ;
        RECT 386.075 239.195 386.405 239.525 ;
        RECT 386.075 237.835 386.405 238.165 ;
        RECT 386.08 237.16 386.4 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 386.075 -1.525 386.405 -1.195 ;
        RECT 386.075 -2.885 386.405 -2.555 ;
        RECT 386.08 -3.56 386.4 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 386.075 -91.285 386.405 -90.955 ;
        RECT 386.075 -92.645 386.405 -92.315 ;
        RECT 386.075 -94.005 386.405 -93.675 ;
        RECT 386.075 -95.365 386.405 -95.035 ;
        RECT 386.075 -96.725 386.405 -96.395 ;
        RECT 386.075 -98.085 386.405 -97.755 ;
        RECT 386.075 -99.445 386.405 -99.115 ;
        RECT 386.075 -100.805 386.405 -100.475 ;
        RECT 386.075 -102.165 386.405 -101.835 ;
        RECT 386.075 -103.525 386.405 -103.195 ;
        RECT 386.075 -104.885 386.405 -104.555 ;
        RECT 386.075 -106.245 386.405 -105.915 ;
        RECT 386.075 -107.605 386.405 -107.275 ;
        RECT 386.075 -108.965 386.405 -108.635 ;
        RECT 386.075 -110.325 386.405 -109.995 ;
        RECT 386.075 -111.685 386.405 -111.355 ;
        RECT 386.075 -113.045 386.405 -112.715 ;
        RECT 386.075 -114.405 386.405 -114.075 ;
        RECT 386.075 -115.765 386.405 -115.435 ;
        RECT 386.075 -117.125 386.405 -116.795 ;
        RECT 386.075 -118.485 386.405 -118.155 ;
        RECT 386.075 -119.845 386.405 -119.515 ;
        RECT 386.075 -121.205 386.405 -120.875 ;
        RECT 386.075 -122.565 386.405 -122.235 ;
        RECT 386.075 -123.925 386.405 -123.595 ;
        RECT 386.075 -125.285 386.405 -124.955 ;
        RECT 386.075 -126.645 386.405 -126.315 ;
        RECT 386.075 -128.005 386.405 -127.675 ;
        RECT 386.075 -129.365 386.405 -129.035 ;
        RECT 386.075 -130.725 386.405 -130.395 ;
        RECT 386.075 -132.085 386.405 -131.755 ;
        RECT 386.075 -133.445 386.405 -133.115 ;
        RECT 386.075 -134.805 386.405 -134.475 ;
        RECT 386.075 -136.165 386.405 -135.835 ;
        RECT 386.075 -137.525 386.405 -137.195 ;
        RECT 386.075 -138.885 386.405 -138.555 ;
        RECT 386.075 -140.245 386.405 -139.915 ;
        RECT 386.075 -141.605 386.405 -141.275 ;
        RECT 386.075 -142.965 386.405 -142.635 ;
        RECT 386.075 -144.325 386.405 -143.995 ;
        RECT 386.075 -145.685 386.405 -145.355 ;
        RECT 386.075 -147.045 386.405 -146.715 ;
        RECT 386.075 -148.405 386.405 -148.075 ;
        RECT 386.075 -149.765 386.405 -149.435 ;
        RECT 386.075 -151.125 386.405 -150.795 ;
        RECT 386.075 -152.485 386.405 -152.155 ;
        RECT 386.075 -153.845 386.405 -153.515 ;
        RECT 386.075 -155.205 386.405 -154.875 ;
        RECT 386.075 -156.565 386.405 -156.235 ;
        RECT 386.075 -157.925 386.405 -157.595 ;
        RECT 386.075 -159.285 386.405 -158.955 ;
        RECT 386.075 -160.645 386.405 -160.315 ;
        RECT 386.075 -162.005 386.405 -161.675 ;
        RECT 386.075 -163.365 386.405 -163.035 ;
        RECT 386.075 -164.725 386.405 -164.395 ;
        RECT 386.075 -166.085 386.405 -165.755 ;
        RECT 386.075 -167.445 386.405 -167.115 ;
        RECT 386.075 -168.805 386.405 -168.475 ;
        RECT 386.075 -170.165 386.405 -169.835 ;
        RECT 386.075 -171.525 386.405 -171.195 ;
        RECT 386.075 -172.885 386.405 -172.555 ;
        RECT 386.075 -174.245 386.405 -173.915 ;
        RECT 386.075 -175.605 386.405 -175.275 ;
        RECT 386.075 -176.965 386.405 -176.635 ;
        RECT 386.075 -178.325 386.405 -177.995 ;
        RECT 386.075 -180.57 386.405 -179.44 ;
        RECT 386.08 -180.685 386.4 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 387.435 241.32 387.765 242.45 ;
        RECT 387.435 239.195 387.765 239.525 ;
        RECT 387.435 237.835 387.765 238.165 ;
        RECT 387.44 237.16 387.76 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 387.435 -95.365 387.765 -95.035 ;
        RECT 387.435 -96.725 387.765 -96.395 ;
        RECT 387.435 -98.085 387.765 -97.755 ;
        RECT 387.435 -99.445 387.765 -99.115 ;
        RECT 387.435 -100.805 387.765 -100.475 ;
        RECT 387.435 -102.165 387.765 -101.835 ;
        RECT 387.435 -103.525 387.765 -103.195 ;
        RECT 387.435 -104.885 387.765 -104.555 ;
        RECT 387.435 -106.245 387.765 -105.915 ;
        RECT 387.435 -107.605 387.765 -107.275 ;
        RECT 387.435 -108.965 387.765 -108.635 ;
        RECT 387.435 -110.325 387.765 -109.995 ;
        RECT 387.435 -111.685 387.765 -111.355 ;
        RECT 387.435 -113.045 387.765 -112.715 ;
        RECT 387.435 -114.405 387.765 -114.075 ;
        RECT 387.435 -115.765 387.765 -115.435 ;
        RECT 387.435 -117.125 387.765 -116.795 ;
        RECT 387.435 -118.485 387.765 -118.155 ;
        RECT 387.435 -119.845 387.765 -119.515 ;
        RECT 387.435 -121.205 387.765 -120.875 ;
        RECT 387.435 -122.565 387.765 -122.235 ;
        RECT 387.435 -123.925 387.765 -123.595 ;
        RECT 387.435 -125.285 387.765 -124.955 ;
        RECT 387.435 -126.645 387.765 -126.315 ;
        RECT 387.435 -128.005 387.765 -127.675 ;
        RECT 387.435 -129.365 387.765 -129.035 ;
        RECT 387.435 -130.725 387.765 -130.395 ;
        RECT 387.435 -132.085 387.765 -131.755 ;
        RECT 387.435 -133.445 387.765 -133.115 ;
        RECT 387.435 -134.805 387.765 -134.475 ;
        RECT 387.435 -136.165 387.765 -135.835 ;
        RECT 387.435 -137.525 387.765 -137.195 ;
        RECT 387.435 -138.885 387.765 -138.555 ;
        RECT 387.435 -140.245 387.765 -139.915 ;
        RECT 387.435 -141.605 387.765 -141.275 ;
        RECT 387.435 -142.965 387.765 -142.635 ;
        RECT 387.435 -144.325 387.765 -143.995 ;
        RECT 387.435 -145.685 387.765 -145.355 ;
        RECT 387.435 -147.045 387.765 -146.715 ;
        RECT 387.435 -148.405 387.765 -148.075 ;
        RECT 387.435 -149.765 387.765 -149.435 ;
        RECT 387.435 -151.125 387.765 -150.795 ;
        RECT 387.435 -152.485 387.765 -152.155 ;
        RECT 387.435 -153.845 387.765 -153.515 ;
        RECT 387.435 -155.205 387.765 -154.875 ;
        RECT 387.435 -156.565 387.765 -156.235 ;
        RECT 387.435 -157.925 387.765 -157.595 ;
        RECT 387.435 -159.285 387.765 -158.955 ;
        RECT 387.435 -160.645 387.765 -160.315 ;
        RECT 387.435 -162.005 387.765 -161.675 ;
        RECT 387.435 -163.365 387.765 -163.035 ;
        RECT 387.435 -164.725 387.765 -164.395 ;
        RECT 387.435 -166.085 387.765 -165.755 ;
        RECT 387.435 -167.445 387.765 -167.115 ;
        RECT 387.435 -168.805 387.765 -168.475 ;
        RECT 387.435 -170.165 387.765 -169.835 ;
        RECT 387.435 -171.525 387.765 -171.195 ;
        RECT 387.435 -172.885 387.765 -172.555 ;
        RECT 387.435 -174.245 387.765 -173.915 ;
        RECT 387.435 -175.605 387.765 -175.275 ;
        RECT 387.435 -176.965 387.765 -176.635 ;
        RECT 387.435 -178.325 387.765 -177.995 ;
        RECT 387.435 -180.57 387.765 -179.44 ;
        RECT 387.44 -180.685 387.76 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 387.61 -94.075 387.94 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 388.795 241.32 389.125 242.45 ;
        RECT 388.795 239.195 389.125 239.525 ;
        RECT 388.795 237.835 389.125 238.165 ;
        RECT 388.8 237.16 389.12 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 388.795 -1.525 389.125 -1.195 ;
        RECT 388.795 -2.885 389.125 -2.555 ;
        RECT 388.8 -3.56 389.12 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 390.155 241.32 390.485 242.45 ;
        RECT 390.155 239.195 390.485 239.525 ;
        RECT 390.155 237.835 390.485 238.165 ;
        RECT 390.16 237.16 390.48 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 390.155 -1.525 390.485 -1.195 ;
        RECT 390.155 -2.885 390.485 -2.555 ;
        RECT 390.16 -3.56 390.48 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 391.515 241.32 391.845 242.45 ;
        RECT 391.515 239.195 391.845 239.525 ;
        RECT 391.515 237.835 391.845 238.165 ;
        RECT 391.52 237.16 391.84 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 391.515 -1.525 391.845 -1.195 ;
        RECT 391.515 -2.885 391.845 -2.555 ;
        RECT 391.52 -3.56 391.84 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 391.515 -91.285 391.845 -90.955 ;
        RECT 391.515 -92.645 391.845 -92.315 ;
        RECT 391.515 -94.005 391.845 -93.675 ;
        RECT 391.515 -95.365 391.845 -95.035 ;
        RECT 391.515 -96.725 391.845 -96.395 ;
        RECT 391.515 -98.085 391.845 -97.755 ;
        RECT 391.515 -99.445 391.845 -99.115 ;
        RECT 391.515 -100.805 391.845 -100.475 ;
        RECT 391.515 -102.165 391.845 -101.835 ;
        RECT 391.515 -103.525 391.845 -103.195 ;
        RECT 391.515 -104.885 391.845 -104.555 ;
        RECT 391.515 -106.245 391.845 -105.915 ;
        RECT 391.515 -107.605 391.845 -107.275 ;
        RECT 391.515 -108.965 391.845 -108.635 ;
        RECT 391.515 -110.325 391.845 -109.995 ;
        RECT 391.515 -111.685 391.845 -111.355 ;
        RECT 391.515 -113.045 391.845 -112.715 ;
        RECT 391.515 -114.405 391.845 -114.075 ;
        RECT 391.515 -115.765 391.845 -115.435 ;
        RECT 391.515 -117.125 391.845 -116.795 ;
        RECT 391.515 -118.485 391.845 -118.155 ;
        RECT 391.515 -119.845 391.845 -119.515 ;
        RECT 391.515 -121.205 391.845 -120.875 ;
        RECT 391.515 -122.565 391.845 -122.235 ;
        RECT 391.515 -123.925 391.845 -123.595 ;
        RECT 391.515 -125.285 391.845 -124.955 ;
        RECT 391.515 -126.645 391.845 -126.315 ;
        RECT 391.515 -128.005 391.845 -127.675 ;
        RECT 391.515 -129.365 391.845 -129.035 ;
        RECT 391.515 -130.725 391.845 -130.395 ;
        RECT 391.515 -132.085 391.845 -131.755 ;
        RECT 391.515 -133.445 391.845 -133.115 ;
        RECT 391.515 -134.805 391.845 -134.475 ;
        RECT 391.515 -136.165 391.845 -135.835 ;
        RECT 391.515 -137.525 391.845 -137.195 ;
        RECT 391.515 -138.885 391.845 -138.555 ;
        RECT 391.515 -140.245 391.845 -139.915 ;
        RECT 391.515 -141.605 391.845 -141.275 ;
        RECT 391.515 -142.965 391.845 -142.635 ;
        RECT 391.515 -144.325 391.845 -143.995 ;
        RECT 391.515 -145.685 391.845 -145.355 ;
        RECT 391.515 -147.045 391.845 -146.715 ;
        RECT 391.515 -148.405 391.845 -148.075 ;
        RECT 391.515 -149.765 391.845 -149.435 ;
        RECT 391.515 -151.125 391.845 -150.795 ;
        RECT 391.515 -152.485 391.845 -152.155 ;
        RECT 391.515 -153.845 391.845 -153.515 ;
        RECT 391.515 -155.205 391.845 -154.875 ;
        RECT 391.515 -156.565 391.845 -156.235 ;
        RECT 391.515 -157.925 391.845 -157.595 ;
        RECT 391.515 -159.285 391.845 -158.955 ;
        RECT 391.515 -160.645 391.845 -160.315 ;
        RECT 391.515 -162.005 391.845 -161.675 ;
        RECT 391.515 -163.365 391.845 -163.035 ;
        RECT 391.515 -164.725 391.845 -164.395 ;
        RECT 391.515 -166.085 391.845 -165.755 ;
        RECT 391.515 -167.445 391.845 -167.115 ;
        RECT 391.515 -168.805 391.845 -168.475 ;
        RECT 391.515 -170.165 391.845 -169.835 ;
        RECT 391.515 -171.525 391.845 -171.195 ;
        RECT 391.515 -172.885 391.845 -172.555 ;
        RECT 391.515 -174.245 391.845 -173.915 ;
        RECT 391.515 -175.605 391.845 -175.275 ;
        RECT 391.515 -176.965 391.845 -176.635 ;
        RECT 391.515 -178.325 391.845 -177.995 ;
        RECT 391.515 -180.57 391.845 -179.44 ;
        RECT 391.52 -180.685 391.84 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 392.875 241.32 393.205 242.45 ;
        RECT 392.875 239.195 393.205 239.525 ;
        RECT 392.875 237.835 393.205 238.165 ;
        RECT 392.88 237.16 393.2 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 392.875 -95.365 393.205 -95.035 ;
        RECT 392.875 -96.725 393.205 -96.395 ;
        RECT 392.875 -98.085 393.205 -97.755 ;
        RECT 392.875 -99.445 393.205 -99.115 ;
        RECT 392.875 -100.805 393.205 -100.475 ;
        RECT 392.875 -102.165 393.205 -101.835 ;
        RECT 392.875 -103.525 393.205 -103.195 ;
        RECT 392.875 -104.885 393.205 -104.555 ;
        RECT 392.875 -106.245 393.205 -105.915 ;
        RECT 392.875 -107.605 393.205 -107.275 ;
        RECT 392.875 -108.965 393.205 -108.635 ;
        RECT 392.875 -110.325 393.205 -109.995 ;
        RECT 392.875 -111.685 393.205 -111.355 ;
        RECT 392.875 -113.045 393.205 -112.715 ;
        RECT 392.875 -114.405 393.205 -114.075 ;
        RECT 392.875 -115.765 393.205 -115.435 ;
        RECT 392.875 -117.125 393.205 -116.795 ;
        RECT 392.875 -118.485 393.205 -118.155 ;
        RECT 392.875 -119.845 393.205 -119.515 ;
        RECT 392.875 -121.205 393.205 -120.875 ;
        RECT 392.875 -122.565 393.205 -122.235 ;
        RECT 392.875 -123.925 393.205 -123.595 ;
        RECT 392.875 -125.285 393.205 -124.955 ;
        RECT 392.875 -126.645 393.205 -126.315 ;
        RECT 392.875 -128.005 393.205 -127.675 ;
        RECT 392.875 -129.365 393.205 -129.035 ;
        RECT 392.875 -130.725 393.205 -130.395 ;
        RECT 392.875 -132.085 393.205 -131.755 ;
        RECT 392.875 -133.445 393.205 -133.115 ;
        RECT 392.875 -134.805 393.205 -134.475 ;
        RECT 392.875 -136.165 393.205 -135.835 ;
        RECT 392.875 -137.525 393.205 -137.195 ;
        RECT 392.875 -138.885 393.205 -138.555 ;
        RECT 392.875 -140.245 393.205 -139.915 ;
        RECT 392.875 -141.605 393.205 -141.275 ;
        RECT 392.875 -142.965 393.205 -142.635 ;
        RECT 392.875 -144.325 393.205 -143.995 ;
        RECT 392.875 -145.685 393.205 -145.355 ;
        RECT 392.875 -147.045 393.205 -146.715 ;
        RECT 392.875 -148.405 393.205 -148.075 ;
        RECT 392.875 -149.765 393.205 -149.435 ;
        RECT 392.875 -151.125 393.205 -150.795 ;
        RECT 392.875 -152.485 393.205 -152.155 ;
        RECT 392.875 -153.845 393.205 -153.515 ;
        RECT 392.875 -155.205 393.205 -154.875 ;
        RECT 392.875 -156.565 393.205 -156.235 ;
        RECT 392.875 -157.925 393.205 -157.595 ;
        RECT 392.875 -159.285 393.205 -158.955 ;
        RECT 392.875 -160.645 393.205 -160.315 ;
        RECT 392.875 -162.005 393.205 -161.675 ;
        RECT 392.875 -163.365 393.205 -163.035 ;
        RECT 392.875 -164.725 393.205 -164.395 ;
        RECT 392.875 -166.085 393.205 -165.755 ;
        RECT 392.875 -167.445 393.205 -167.115 ;
        RECT 392.875 -168.805 393.205 -168.475 ;
        RECT 392.875 -170.165 393.205 -169.835 ;
        RECT 392.875 -171.525 393.205 -171.195 ;
        RECT 392.875 -172.885 393.205 -172.555 ;
        RECT 392.875 -174.245 393.205 -173.915 ;
        RECT 392.875 -175.605 393.205 -175.275 ;
        RECT 392.875 -176.965 393.205 -176.635 ;
        RECT 392.875 -178.325 393.205 -177.995 ;
        RECT 392.875 -180.57 393.205 -179.44 ;
        RECT 392.88 -180.685 393.2 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 393.06 -94.075 393.39 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 394.235 241.32 394.565 242.45 ;
        RECT 394.235 239.195 394.565 239.525 ;
        RECT 394.235 237.835 394.565 238.165 ;
        RECT 394.24 237.16 394.56 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 394.235 -95.365 394.565 -95.035 ;
        RECT 394.235 -96.725 394.565 -96.395 ;
        RECT 394.235 -98.085 394.565 -97.755 ;
        RECT 394.235 -99.445 394.565 -99.115 ;
        RECT 394.235 -100.805 394.565 -100.475 ;
        RECT 394.235 -102.165 394.565 -101.835 ;
        RECT 394.235 -103.525 394.565 -103.195 ;
        RECT 394.235 -104.885 394.565 -104.555 ;
        RECT 394.235 -106.245 394.565 -105.915 ;
        RECT 394.235 -107.605 394.565 -107.275 ;
        RECT 394.235 -108.965 394.565 -108.635 ;
        RECT 394.235 -110.325 394.565 -109.995 ;
        RECT 394.235 -111.685 394.565 -111.355 ;
        RECT 394.235 -113.045 394.565 -112.715 ;
        RECT 394.235 -114.405 394.565 -114.075 ;
        RECT 394.235 -115.765 394.565 -115.435 ;
        RECT 394.235 -117.125 394.565 -116.795 ;
        RECT 394.235 -118.485 394.565 -118.155 ;
        RECT 394.235 -119.845 394.565 -119.515 ;
        RECT 394.235 -121.205 394.565 -120.875 ;
        RECT 394.235 -122.565 394.565 -122.235 ;
        RECT 394.235 -123.925 394.565 -123.595 ;
        RECT 394.235 -125.285 394.565 -124.955 ;
        RECT 394.235 -126.645 394.565 -126.315 ;
        RECT 394.235 -128.005 394.565 -127.675 ;
        RECT 394.235 -129.365 394.565 -129.035 ;
        RECT 394.235 -130.725 394.565 -130.395 ;
        RECT 394.235 -132.085 394.565 -131.755 ;
        RECT 394.235 -133.445 394.565 -133.115 ;
        RECT 394.235 -134.805 394.565 -134.475 ;
        RECT 394.235 -136.165 394.565 -135.835 ;
        RECT 394.235 -137.525 394.565 -137.195 ;
        RECT 394.235 -138.885 394.565 -138.555 ;
        RECT 394.235 -140.245 394.565 -139.915 ;
        RECT 394.235 -141.605 394.565 -141.275 ;
        RECT 394.235 -142.965 394.565 -142.635 ;
        RECT 394.235 -144.325 394.565 -143.995 ;
        RECT 394.235 -145.685 394.565 -145.355 ;
        RECT 394.235 -147.045 394.565 -146.715 ;
        RECT 394.235 -148.405 394.565 -148.075 ;
        RECT 394.235 -149.765 394.565 -149.435 ;
        RECT 394.235 -151.125 394.565 -150.795 ;
        RECT 394.235 -152.485 394.565 -152.155 ;
        RECT 394.235 -153.845 394.565 -153.515 ;
        RECT 394.235 -155.205 394.565 -154.875 ;
        RECT 394.235 -156.565 394.565 -156.235 ;
        RECT 394.235 -157.925 394.565 -157.595 ;
        RECT 394.235 -159.285 394.565 -158.955 ;
        RECT 394.235 -160.645 394.565 -160.315 ;
        RECT 394.235 -162.005 394.565 -161.675 ;
        RECT 394.235 -163.365 394.565 -163.035 ;
        RECT 394.235 -164.725 394.565 -164.395 ;
        RECT 394.235 -166.085 394.565 -165.755 ;
        RECT 394.235 -167.445 394.565 -167.115 ;
        RECT 394.235 -168.805 394.565 -168.475 ;
        RECT 394.235 -170.165 394.565 -169.835 ;
        RECT 394.235 -171.525 394.565 -171.195 ;
        RECT 394.235 -172.885 394.565 -172.555 ;
        RECT 394.235 -174.245 394.565 -173.915 ;
        RECT 394.235 -175.605 394.565 -175.275 ;
        RECT 394.235 -176.965 394.565 -176.635 ;
        RECT 394.235 -178.325 394.565 -177.995 ;
        RECT 394.235 -180.57 394.565 -179.44 ;
        RECT 394.24 -180.685 394.56 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 395.595 241.32 395.925 242.45 ;
        RECT 395.595 239.195 395.925 239.525 ;
        RECT 395.595 237.835 395.925 238.165 ;
        RECT 395.6 237.16 395.92 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 395.595 -1.525 395.925 -1.195 ;
        RECT 395.595 -2.885 395.925 -2.555 ;
        RECT 395.6 -3.56 395.92 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 395.595 -91.285 395.925 -90.955 ;
        RECT 395.595 -92.645 395.925 -92.315 ;
        RECT 395.595 -94.005 395.925 -93.675 ;
        RECT 395.595 -95.365 395.925 -95.035 ;
        RECT 395.595 -96.725 395.925 -96.395 ;
        RECT 395.595 -98.085 395.925 -97.755 ;
        RECT 395.595 -99.445 395.925 -99.115 ;
        RECT 395.595 -100.805 395.925 -100.475 ;
        RECT 395.595 -102.165 395.925 -101.835 ;
        RECT 395.595 -103.525 395.925 -103.195 ;
        RECT 395.595 -104.885 395.925 -104.555 ;
        RECT 395.595 -106.245 395.925 -105.915 ;
        RECT 395.595 -107.605 395.925 -107.275 ;
        RECT 395.595 -108.965 395.925 -108.635 ;
        RECT 395.595 -110.325 395.925 -109.995 ;
        RECT 395.595 -111.685 395.925 -111.355 ;
        RECT 395.595 -113.045 395.925 -112.715 ;
        RECT 395.595 -114.405 395.925 -114.075 ;
        RECT 395.595 -115.765 395.925 -115.435 ;
        RECT 395.595 -117.125 395.925 -116.795 ;
        RECT 395.595 -118.485 395.925 -118.155 ;
        RECT 395.595 -119.845 395.925 -119.515 ;
        RECT 395.595 -121.205 395.925 -120.875 ;
        RECT 395.595 -122.565 395.925 -122.235 ;
        RECT 395.595 -123.925 395.925 -123.595 ;
        RECT 395.595 -125.285 395.925 -124.955 ;
        RECT 395.595 -126.645 395.925 -126.315 ;
        RECT 395.595 -128.005 395.925 -127.675 ;
        RECT 395.595 -129.365 395.925 -129.035 ;
        RECT 395.595 -130.725 395.925 -130.395 ;
        RECT 395.595 -132.085 395.925 -131.755 ;
        RECT 395.595 -133.445 395.925 -133.115 ;
        RECT 395.595 -134.805 395.925 -134.475 ;
        RECT 395.595 -136.165 395.925 -135.835 ;
        RECT 395.595 -137.525 395.925 -137.195 ;
        RECT 395.595 -138.885 395.925 -138.555 ;
        RECT 395.595 -140.245 395.925 -139.915 ;
        RECT 395.595 -141.605 395.925 -141.275 ;
        RECT 395.595 -142.965 395.925 -142.635 ;
        RECT 395.595 -144.325 395.925 -143.995 ;
        RECT 395.595 -145.685 395.925 -145.355 ;
        RECT 395.595 -147.045 395.925 -146.715 ;
        RECT 395.595 -148.405 395.925 -148.075 ;
        RECT 395.595 -149.765 395.925 -149.435 ;
        RECT 395.595 -151.125 395.925 -150.795 ;
        RECT 395.595 -152.485 395.925 -152.155 ;
        RECT 395.595 -153.845 395.925 -153.515 ;
        RECT 395.595 -155.205 395.925 -154.875 ;
        RECT 395.595 -156.565 395.925 -156.235 ;
        RECT 395.595 -157.925 395.925 -157.595 ;
        RECT 395.595 -159.285 395.925 -158.955 ;
        RECT 395.595 -160.645 395.925 -160.315 ;
        RECT 395.595 -162.005 395.925 -161.675 ;
        RECT 395.595 -163.365 395.925 -163.035 ;
        RECT 395.595 -164.725 395.925 -164.395 ;
        RECT 395.595 -166.085 395.925 -165.755 ;
        RECT 395.595 -167.445 395.925 -167.115 ;
        RECT 395.595 -168.805 395.925 -168.475 ;
        RECT 395.595 -170.165 395.925 -169.835 ;
        RECT 395.595 -171.525 395.925 -171.195 ;
        RECT 395.595 -172.885 395.925 -172.555 ;
        RECT 395.595 -174.245 395.925 -173.915 ;
        RECT 395.595 -175.605 395.925 -175.275 ;
        RECT 395.595 -176.965 395.925 -176.635 ;
        RECT 395.595 -178.325 395.925 -177.995 ;
        RECT 395.595 -180.57 395.925 -179.44 ;
        RECT 395.6 -180.685 395.92 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 396.955 241.32 397.285 242.45 ;
        RECT 396.955 239.195 397.285 239.525 ;
        RECT 396.955 237.835 397.285 238.165 ;
        RECT 396.96 237.16 397.28 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 396.955 -1.525 397.285 -1.195 ;
        RECT 396.955 -2.885 397.285 -2.555 ;
        RECT 396.96 -3.56 397.28 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 396.955 -103.525 397.285 -103.195 ;
        RECT 396.955 -104.885 397.285 -104.555 ;
        RECT 396.955 -106.245 397.285 -105.915 ;
        RECT 396.955 -107.605 397.285 -107.275 ;
        RECT 396.955 -108.965 397.285 -108.635 ;
        RECT 396.955 -110.325 397.285 -109.995 ;
        RECT 396.955 -111.685 397.285 -111.355 ;
        RECT 396.955 -113.045 397.285 -112.715 ;
        RECT 396.955 -114.405 397.285 -114.075 ;
        RECT 396.955 -115.765 397.285 -115.435 ;
        RECT 396.955 -117.125 397.285 -116.795 ;
        RECT 396.955 -118.485 397.285 -118.155 ;
        RECT 396.955 -119.845 397.285 -119.515 ;
        RECT 396.955 -121.205 397.285 -120.875 ;
        RECT 396.955 -122.565 397.285 -122.235 ;
        RECT 396.955 -123.925 397.285 -123.595 ;
        RECT 396.955 -125.285 397.285 -124.955 ;
        RECT 396.955 -126.645 397.285 -126.315 ;
        RECT 396.955 -128.005 397.285 -127.675 ;
        RECT 396.955 -129.365 397.285 -129.035 ;
        RECT 396.955 -130.725 397.285 -130.395 ;
        RECT 396.955 -132.085 397.285 -131.755 ;
        RECT 396.955 -133.445 397.285 -133.115 ;
        RECT 396.955 -134.805 397.285 -134.475 ;
        RECT 396.955 -136.165 397.285 -135.835 ;
        RECT 396.955 -137.525 397.285 -137.195 ;
        RECT 396.955 -138.885 397.285 -138.555 ;
        RECT 396.955 -140.245 397.285 -139.915 ;
        RECT 396.955 -141.605 397.285 -141.275 ;
        RECT 396.955 -142.965 397.285 -142.635 ;
        RECT 396.955 -144.325 397.285 -143.995 ;
        RECT 396.955 -145.685 397.285 -145.355 ;
        RECT 396.955 -147.045 397.285 -146.715 ;
        RECT 396.955 -148.405 397.285 -148.075 ;
        RECT 396.955 -149.765 397.285 -149.435 ;
        RECT 396.955 -151.125 397.285 -150.795 ;
        RECT 396.955 -152.485 397.285 -152.155 ;
        RECT 396.955 -153.845 397.285 -153.515 ;
        RECT 396.955 -155.205 397.285 -154.875 ;
        RECT 396.955 -156.565 397.285 -156.235 ;
        RECT 396.955 -157.925 397.285 -157.595 ;
        RECT 396.955 -159.285 397.285 -158.955 ;
        RECT 396.955 -160.645 397.285 -160.315 ;
        RECT 396.955 -162.005 397.285 -161.675 ;
        RECT 396.955 -163.365 397.285 -163.035 ;
        RECT 396.955 -164.725 397.285 -164.395 ;
        RECT 396.955 -166.085 397.285 -165.755 ;
        RECT 396.955 -167.445 397.285 -167.115 ;
        RECT 396.955 -168.805 397.285 -168.475 ;
        RECT 396.955 -170.165 397.285 -169.835 ;
        RECT 396.955 -171.525 397.285 -171.195 ;
        RECT 396.955 -172.885 397.285 -172.555 ;
        RECT 396.955 -174.245 397.285 -173.915 ;
        RECT 396.955 -175.605 397.285 -175.275 ;
        RECT 396.955 -176.965 397.285 -176.635 ;
        RECT 396.955 -178.325 397.285 -177.995 ;
        RECT 396.955 -180.57 397.285 -179.44 ;
        RECT 396.96 -180.685 397.28 -90.955 ;
        RECT 396.955 -91.285 397.285 -90.955 ;
        RECT 396.955 -92.645 397.285 -92.315 ;
        RECT 396.955 -94.005 397.285 -93.675 ;
        RECT 396.955 -95.365 397.285 -95.035 ;
        RECT 396.955 -96.725 397.285 -96.395 ;
        RECT 396.955 -98.085 397.285 -97.755 ;
        RECT 396.955 -99.445 397.285 -99.115 ;
        RECT 396.955 -100.805 397.285 -100.475 ;
        RECT 396.955 -102.165 397.285 -101.835 ;
    END
    PORT
      LAYER met3 ;
        RECT 337.115 241.32 337.445 242.45 ;
        RECT 337.115 239.195 337.445 239.525 ;
        RECT 337.115 237.835 337.445 238.165 ;
        RECT 337.12 237.16 337.44 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 337.115 -1.525 337.445 -1.195 ;
        RECT 337.115 -2.885 337.445 -2.555 ;
        RECT 337.12 -3.56 337.44 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 337.115 -91.285 337.445 -90.955 ;
        RECT 337.115 -92.645 337.445 -92.315 ;
        RECT 337.115 -94.005 337.445 -93.675 ;
        RECT 337.115 -95.365 337.445 -95.035 ;
        RECT 337.115 -96.725 337.445 -96.395 ;
        RECT 337.115 -98.085 337.445 -97.755 ;
        RECT 337.115 -99.445 337.445 -99.115 ;
        RECT 337.115 -100.805 337.445 -100.475 ;
        RECT 337.115 -102.165 337.445 -101.835 ;
        RECT 337.115 -103.525 337.445 -103.195 ;
        RECT 337.115 -104.885 337.445 -104.555 ;
        RECT 337.115 -106.245 337.445 -105.915 ;
        RECT 337.115 -107.605 337.445 -107.275 ;
        RECT 337.115 -108.965 337.445 -108.635 ;
        RECT 337.115 -110.325 337.445 -109.995 ;
        RECT 337.115 -111.685 337.445 -111.355 ;
        RECT 337.115 -113.045 337.445 -112.715 ;
        RECT 337.115 -114.405 337.445 -114.075 ;
        RECT 337.115 -115.765 337.445 -115.435 ;
        RECT 337.115 -117.125 337.445 -116.795 ;
        RECT 337.115 -118.485 337.445 -118.155 ;
        RECT 337.115 -119.845 337.445 -119.515 ;
        RECT 337.115 -121.205 337.445 -120.875 ;
        RECT 337.115 -122.565 337.445 -122.235 ;
        RECT 337.115 -123.925 337.445 -123.595 ;
        RECT 337.115 -125.285 337.445 -124.955 ;
        RECT 337.115 -126.645 337.445 -126.315 ;
        RECT 337.115 -128.005 337.445 -127.675 ;
        RECT 337.115 -129.365 337.445 -129.035 ;
        RECT 337.115 -130.725 337.445 -130.395 ;
        RECT 337.115 -132.085 337.445 -131.755 ;
        RECT 337.115 -133.445 337.445 -133.115 ;
        RECT 337.115 -134.805 337.445 -134.475 ;
        RECT 337.115 -136.165 337.445 -135.835 ;
        RECT 337.115 -137.525 337.445 -137.195 ;
        RECT 337.115 -138.885 337.445 -138.555 ;
        RECT 337.115 -140.245 337.445 -139.915 ;
        RECT 337.115 -141.605 337.445 -141.275 ;
        RECT 337.115 -142.965 337.445 -142.635 ;
        RECT 337.115 -144.325 337.445 -143.995 ;
        RECT 337.115 -145.685 337.445 -145.355 ;
        RECT 337.115 -147.045 337.445 -146.715 ;
        RECT 337.115 -148.405 337.445 -148.075 ;
        RECT 337.115 -149.765 337.445 -149.435 ;
        RECT 337.115 -151.125 337.445 -150.795 ;
        RECT 337.115 -152.485 337.445 -152.155 ;
        RECT 337.115 -153.845 337.445 -153.515 ;
        RECT 337.115 -155.205 337.445 -154.875 ;
        RECT 337.115 -156.565 337.445 -156.235 ;
        RECT 337.115 -157.925 337.445 -157.595 ;
        RECT 337.115 -159.285 337.445 -158.955 ;
        RECT 337.115 -160.645 337.445 -160.315 ;
        RECT 337.115 -162.005 337.445 -161.675 ;
        RECT 337.115 -163.365 337.445 -163.035 ;
        RECT 337.115 -164.725 337.445 -164.395 ;
        RECT 337.115 -166.085 337.445 -165.755 ;
        RECT 337.115 -167.445 337.445 -167.115 ;
        RECT 337.115 -168.805 337.445 -168.475 ;
        RECT 337.115 -170.165 337.445 -169.835 ;
        RECT 337.115 -171.525 337.445 -171.195 ;
        RECT 337.115 -172.885 337.445 -172.555 ;
        RECT 337.115 -174.245 337.445 -173.915 ;
        RECT 337.115 -175.605 337.445 -175.275 ;
        RECT 337.115 -176.965 337.445 -176.635 ;
        RECT 337.115 -178.325 337.445 -177.995 ;
        RECT 337.115 -180.57 337.445 -179.44 ;
        RECT 337.12 -180.685 337.44 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 338.475 241.32 338.805 242.45 ;
        RECT 338.475 239.195 338.805 239.525 ;
        RECT 338.475 237.835 338.805 238.165 ;
        RECT 338.48 237.16 338.8 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 338.475 -95.365 338.805 -95.035 ;
        RECT 338.475 -96.725 338.805 -96.395 ;
        RECT 338.475 -98.085 338.805 -97.755 ;
        RECT 338.475 -99.445 338.805 -99.115 ;
        RECT 338.475 -100.805 338.805 -100.475 ;
        RECT 338.475 -102.165 338.805 -101.835 ;
        RECT 338.475 -103.525 338.805 -103.195 ;
        RECT 338.475 -104.885 338.805 -104.555 ;
        RECT 338.475 -106.245 338.805 -105.915 ;
        RECT 338.475 -107.605 338.805 -107.275 ;
        RECT 338.475 -108.965 338.805 -108.635 ;
        RECT 338.475 -110.325 338.805 -109.995 ;
        RECT 338.475 -111.685 338.805 -111.355 ;
        RECT 338.475 -113.045 338.805 -112.715 ;
        RECT 338.475 -114.405 338.805 -114.075 ;
        RECT 338.475 -115.765 338.805 -115.435 ;
        RECT 338.475 -117.125 338.805 -116.795 ;
        RECT 338.475 -118.485 338.805 -118.155 ;
        RECT 338.475 -119.845 338.805 -119.515 ;
        RECT 338.475 -121.205 338.805 -120.875 ;
        RECT 338.475 -122.565 338.805 -122.235 ;
        RECT 338.475 -123.925 338.805 -123.595 ;
        RECT 338.475 -125.285 338.805 -124.955 ;
        RECT 338.475 -126.645 338.805 -126.315 ;
        RECT 338.475 -128.005 338.805 -127.675 ;
        RECT 338.475 -129.365 338.805 -129.035 ;
        RECT 338.475 -130.725 338.805 -130.395 ;
        RECT 338.475 -132.085 338.805 -131.755 ;
        RECT 338.475 -133.445 338.805 -133.115 ;
        RECT 338.475 -134.805 338.805 -134.475 ;
        RECT 338.475 -136.165 338.805 -135.835 ;
        RECT 338.475 -137.525 338.805 -137.195 ;
        RECT 338.475 -138.885 338.805 -138.555 ;
        RECT 338.475 -140.245 338.805 -139.915 ;
        RECT 338.475 -141.605 338.805 -141.275 ;
        RECT 338.475 -142.965 338.805 -142.635 ;
        RECT 338.475 -144.325 338.805 -143.995 ;
        RECT 338.475 -145.685 338.805 -145.355 ;
        RECT 338.475 -147.045 338.805 -146.715 ;
        RECT 338.475 -148.405 338.805 -148.075 ;
        RECT 338.475 -149.765 338.805 -149.435 ;
        RECT 338.475 -151.125 338.805 -150.795 ;
        RECT 338.475 -152.485 338.805 -152.155 ;
        RECT 338.475 -153.845 338.805 -153.515 ;
        RECT 338.475 -155.205 338.805 -154.875 ;
        RECT 338.475 -156.565 338.805 -156.235 ;
        RECT 338.475 -157.925 338.805 -157.595 ;
        RECT 338.475 -159.285 338.805 -158.955 ;
        RECT 338.475 -160.645 338.805 -160.315 ;
        RECT 338.475 -162.005 338.805 -161.675 ;
        RECT 338.475 -163.365 338.805 -163.035 ;
        RECT 338.475 -164.725 338.805 -164.395 ;
        RECT 338.475 -166.085 338.805 -165.755 ;
        RECT 338.475 -167.445 338.805 -167.115 ;
        RECT 338.475 -168.805 338.805 -168.475 ;
        RECT 338.475 -170.165 338.805 -169.835 ;
        RECT 338.475 -171.525 338.805 -171.195 ;
        RECT 338.475 -172.885 338.805 -172.555 ;
        RECT 338.475 -174.245 338.805 -173.915 ;
        RECT 338.475 -175.605 338.805 -175.275 ;
        RECT 338.475 -176.965 338.805 -176.635 ;
        RECT 338.475 -178.325 338.805 -177.995 ;
        RECT 338.475 -180.57 338.805 -179.44 ;
        RECT 338.48 -180.685 338.8 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 338.81 -94.075 339.14 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 339.835 241.32 340.165 242.45 ;
        RECT 339.835 239.195 340.165 239.525 ;
        RECT 339.835 237.835 340.165 238.165 ;
        RECT 339.84 237.16 340.16 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 339.835 -1.525 340.165 -1.195 ;
        RECT 339.835 -2.885 340.165 -2.555 ;
        RECT 339.84 -3.56 340.16 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 341.195 241.32 341.525 242.45 ;
        RECT 341.195 239.195 341.525 239.525 ;
        RECT 341.195 237.835 341.525 238.165 ;
        RECT 341.2 237.16 341.52 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 341.195 -1.525 341.525 -1.195 ;
        RECT 341.195 -2.885 341.525 -2.555 ;
        RECT 341.2 -3.56 341.52 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 342.555 241.32 342.885 242.45 ;
        RECT 342.555 239.195 342.885 239.525 ;
        RECT 342.555 237.835 342.885 238.165 ;
        RECT 342.56 237.16 342.88 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 342.555 -1.525 342.885 -1.195 ;
        RECT 342.555 -2.885 342.885 -2.555 ;
        RECT 342.56 -3.56 342.88 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 342.555 -91.285 342.885 -90.955 ;
        RECT 342.555 -92.645 342.885 -92.315 ;
        RECT 342.555 -94.005 342.885 -93.675 ;
        RECT 342.555 -95.365 342.885 -95.035 ;
        RECT 342.555 -96.725 342.885 -96.395 ;
        RECT 342.555 -98.085 342.885 -97.755 ;
        RECT 342.555 -99.445 342.885 -99.115 ;
        RECT 342.555 -100.805 342.885 -100.475 ;
        RECT 342.555 -102.165 342.885 -101.835 ;
        RECT 342.555 -103.525 342.885 -103.195 ;
        RECT 342.555 -104.885 342.885 -104.555 ;
        RECT 342.555 -106.245 342.885 -105.915 ;
        RECT 342.555 -107.605 342.885 -107.275 ;
        RECT 342.555 -108.965 342.885 -108.635 ;
        RECT 342.555 -110.325 342.885 -109.995 ;
        RECT 342.555 -111.685 342.885 -111.355 ;
        RECT 342.555 -113.045 342.885 -112.715 ;
        RECT 342.555 -114.405 342.885 -114.075 ;
        RECT 342.555 -115.765 342.885 -115.435 ;
        RECT 342.555 -117.125 342.885 -116.795 ;
        RECT 342.555 -118.485 342.885 -118.155 ;
        RECT 342.555 -119.845 342.885 -119.515 ;
        RECT 342.555 -121.205 342.885 -120.875 ;
        RECT 342.555 -122.565 342.885 -122.235 ;
        RECT 342.555 -123.925 342.885 -123.595 ;
        RECT 342.555 -125.285 342.885 -124.955 ;
        RECT 342.555 -126.645 342.885 -126.315 ;
        RECT 342.555 -128.005 342.885 -127.675 ;
        RECT 342.555 -129.365 342.885 -129.035 ;
        RECT 342.555 -130.725 342.885 -130.395 ;
        RECT 342.555 -132.085 342.885 -131.755 ;
        RECT 342.555 -133.445 342.885 -133.115 ;
        RECT 342.555 -134.805 342.885 -134.475 ;
        RECT 342.555 -136.165 342.885 -135.835 ;
        RECT 342.555 -137.525 342.885 -137.195 ;
        RECT 342.555 -138.885 342.885 -138.555 ;
        RECT 342.555 -140.245 342.885 -139.915 ;
        RECT 342.555 -141.605 342.885 -141.275 ;
        RECT 342.555 -142.965 342.885 -142.635 ;
        RECT 342.555 -144.325 342.885 -143.995 ;
        RECT 342.555 -145.685 342.885 -145.355 ;
        RECT 342.555 -147.045 342.885 -146.715 ;
        RECT 342.555 -148.405 342.885 -148.075 ;
        RECT 342.555 -149.765 342.885 -149.435 ;
        RECT 342.555 -151.125 342.885 -150.795 ;
        RECT 342.555 -152.485 342.885 -152.155 ;
        RECT 342.555 -153.845 342.885 -153.515 ;
        RECT 342.555 -155.205 342.885 -154.875 ;
        RECT 342.555 -156.565 342.885 -156.235 ;
        RECT 342.555 -157.925 342.885 -157.595 ;
        RECT 342.555 -159.285 342.885 -158.955 ;
        RECT 342.555 -160.645 342.885 -160.315 ;
        RECT 342.555 -162.005 342.885 -161.675 ;
        RECT 342.555 -163.365 342.885 -163.035 ;
        RECT 342.555 -164.725 342.885 -164.395 ;
        RECT 342.555 -166.085 342.885 -165.755 ;
        RECT 342.555 -167.445 342.885 -167.115 ;
        RECT 342.555 -168.805 342.885 -168.475 ;
        RECT 342.555 -170.165 342.885 -169.835 ;
        RECT 342.555 -171.525 342.885 -171.195 ;
        RECT 342.555 -172.885 342.885 -172.555 ;
        RECT 342.555 -174.245 342.885 -173.915 ;
        RECT 342.555 -175.605 342.885 -175.275 ;
        RECT 342.555 -176.965 342.885 -176.635 ;
        RECT 342.555 -178.325 342.885 -177.995 ;
        RECT 342.555 -180.57 342.885 -179.44 ;
        RECT 342.56 -180.685 342.88 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 343.915 241.32 344.245 242.45 ;
        RECT 343.915 239.195 344.245 239.525 ;
        RECT 343.915 237.835 344.245 238.165 ;
        RECT 343.92 237.16 344.24 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 343.915 -95.365 344.245 -95.035 ;
        RECT 343.915 -96.725 344.245 -96.395 ;
        RECT 343.915 -98.085 344.245 -97.755 ;
        RECT 343.915 -99.445 344.245 -99.115 ;
        RECT 343.915 -100.805 344.245 -100.475 ;
        RECT 343.915 -102.165 344.245 -101.835 ;
        RECT 343.915 -103.525 344.245 -103.195 ;
        RECT 343.915 -104.885 344.245 -104.555 ;
        RECT 343.915 -106.245 344.245 -105.915 ;
        RECT 343.915 -107.605 344.245 -107.275 ;
        RECT 343.915 -108.965 344.245 -108.635 ;
        RECT 343.915 -110.325 344.245 -109.995 ;
        RECT 343.915 -111.685 344.245 -111.355 ;
        RECT 343.915 -113.045 344.245 -112.715 ;
        RECT 343.915 -114.405 344.245 -114.075 ;
        RECT 343.915 -115.765 344.245 -115.435 ;
        RECT 343.915 -117.125 344.245 -116.795 ;
        RECT 343.915 -118.485 344.245 -118.155 ;
        RECT 343.915 -119.845 344.245 -119.515 ;
        RECT 343.915 -121.205 344.245 -120.875 ;
        RECT 343.915 -122.565 344.245 -122.235 ;
        RECT 343.915 -123.925 344.245 -123.595 ;
        RECT 343.915 -125.285 344.245 -124.955 ;
        RECT 343.915 -126.645 344.245 -126.315 ;
        RECT 343.915 -128.005 344.245 -127.675 ;
        RECT 343.915 -129.365 344.245 -129.035 ;
        RECT 343.915 -130.725 344.245 -130.395 ;
        RECT 343.915 -132.085 344.245 -131.755 ;
        RECT 343.915 -133.445 344.245 -133.115 ;
        RECT 343.915 -134.805 344.245 -134.475 ;
        RECT 343.915 -136.165 344.245 -135.835 ;
        RECT 343.915 -137.525 344.245 -137.195 ;
        RECT 343.915 -138.885 344.245 -138.555 ;
        RECT 343.915 -140.245 344.245 -139.915 ;
        RECT 343.915 -141.605 344.245 -141.275 ;
        RECT 343.915 -142.965 344.245 -142.635 ;
        RECT 343.915 -144.325 344.245 -143.995 ;
        RECT 343.915 -145.685 344.245 -145.355 ;
        RECT 343.915 -147.045 344.245 -146.715 ;
        RECT 343.915 -148.405 344.245 -148.075 ;
        RECT 343.915 -149.765 344.245 -149.435 ;
        RECT 343.915 -151.125 344.245 -150.795 ;
        RECT 343.915 -152.485 344.245 -152.155 ;
        RECT 343.915 -153.845 344.245 -153.515 ;
        RECT 343.915 -155.205 344.245 -154.875 ;
        RECT 343.915 -156.565 344.245 -156.235 ;
        RECT 343.915 -157.925 344.245 -157.595 ;
        RECT 343.915 -159.285 344.245 -158.955 ;
        RECT 343.915 -160.645 344.245 -160.315 ;
        RECT 343.915 -162.005 344.245 -161.675 ;
        RECT 343.915 -163.365 344.245 -163.035 ;
        RECT 343.915 -164.725 344.245 -164.395 ;
        RECT 343.915 -166.085 344.245 -165.755 ;
        RECT 343.915 -167.445 344.245 -167.115 ;
        RECT 343.915 -168.805 344.245 -168.475 ;
        RECT 343.915 -170.165 344.245 -169.835 ;
        RECT 343.915 -171.525 344.245 -171.195 ;
        RECT 343.915 -172.885 344.245 -172.555 ;
        RECT 343.915 -174.245 344.245 -173.915 ;
        RECT 343.915 -175.605 344.245 -175.275 ;
        RECT 343.915 -176.965 344.245 -176.635 ;
        RECT 343.915 -178.325 344.245 -177.995 ;
        RECT 343.915 -180.57 344.245 -179.44 ;
        RECT 343.92 -180.685 344.24 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 344.91 -94.075 345.24 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 345.275 241.32 345.605 242.45 ;
        RECT 345.275 239.195 345.605 239.525 ;
        RECT 345.275 237.835 345.605 238.165 ;
        RECT 345.28 237.16 345.6 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 346.635 241.32 346.965 242.45 ;
        RECT 346.635 239.195 346.965 239.525 ;
        RECT 346.635 237.835 346.965 238.165 ;
        RECT 346.64 237.16 346.96 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 346.635 -1.525 346.965 -1.195 ;
        RECT 346.635 -2.885 346.965 -2.555 ;
        RECT 346.64 -3.56 346.96 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 347.995 241.32 348.325 242.45 ;
        RECT 347.995 239.195 348.325 239.525 ;
        RECT 347.995 237.835 348.325 238.165 ;
        RECT 348 237.16 348.32 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 347.995 -1.525 348.325 -1.195 ;
        RECT 347.995 -2.885 348.325 -2.555 ;
        RECT 348 -3.56 348.32 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 349.355 241.32 349.685 242.45 ;
        RECT 349.355 239.195 349.685 239.525 ;
        RECT 349.355 237.835 349.685 238.165 ;
        RECT 349.36 237.16 349.68 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 349.355 -1.525 349.685 -1.195 ;
        RECT 349.355 -2.885 349.685 -2.555 ;
        RECT 349.36 -3.56 349.68 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 349.355 -91.285 349.685 -90.955 ;
        RECT 349.355 -92.645 349.685 -92.315 ;
        RECT 349.355 -94.005 349.685 -93.675 ;
        RECT 349.355 -95.365 349.685 -95.035 ;
        RECT 349.355 -96.725 349.685 -96.395 ;
        RECT 349.355 -98.085 349.685 -97.755 ;
        RECT 349.355 -99.445 349.685 -99.115 ;
        RECT 349.355 -100.805 349.685 -100.475 ;
        RECT 349.355 -102.165 349.685 -101.835 ;
        RECT 349.355 -103.525 349.685 -103.195 ;
        RECT 349.355 -104.885 349.685 -104.555 ;
        RECT 349.355 -106.245 349.685 -105.915 ;
        RECT 349.355 -107.605 349.685 -107.275 ;
        RECT 349.355 -108.965 349.685 -108.635 ;
        RECT 349.355 -110.325 349.685 -109.995 ;
        RECT 349.355 -111.685 349.685 -111.355 ;
        RECT 349.355 -113.045 349.685 -112.715 ;
        RECT 349.355 -114.405 349.685 -114.075 ;
        RECT 349.355 -115.765 349.685 -115.435 ;
        RECT 349.355 -117.125 349.685 -116.795 ;
        RECT 349.355 -118.485 349.685 -118.155 ;
        RECT 349.355 -119.845 349.685 -119.515 ;
        RECT 349.355 -121.205 349.685 -120.875 ;
        RECT 349.355 -122.565 349.685 -122.235 ;
        RECT 349.355 -123.925 349.685 -123.595 ;
        RECT 349.355 -125.285 349.685 -124.955 ;
        RECT 349.355 -126.645 349.685 -126.315 ;
        RECT 349.355 -128.005 349.685 -127.675 ;
        RECT 349.355 -129.365 349.685 -129.035 ;
        RECT 349.355 -130.725 349.685 -130.395 ;
        RECT 349.355 -132.085 349.685 -131.755 ;
        RECT 349.355 -133.445 349.685 -133.115 ;
        RECT 349.355 -134.805 349.685 -134.475 ;
        RECT 349.355 -136.165 349.685 -135.835 ;
        RECT 349.355 -137.525 349.685 -137.195 ;
        RECT 349.355 -138.885 349.685 -138.555 ;
        RECT 349.355 -140.245 349.685 -139.915 ;
        RECT 349.355 -141.605 349.685 -141.275 ;
        RECT 349.355 -142.965 349.685 -142.635 ;
        RECT 349.355 -144.325 349.685 -143.995 ;
        RECT 349.355 -145.685 349.685 -145.355 ;
        RECT 349.355 -147.045 349.685 -146.715 ;
        RECT 349.355 -148.405 349.685 -148.075 ;
        RECT 349.355 -149.765 349.685 -149.435 ;
        RECT 349.355 -151.125 349.685 -150.795 ;
        RECT 349.355 -152.485 349.685 -152.155 ;
        RECT 349.355 -153.845 349.685 -153.515 ;
        RECT 349.355 -155.205 349.685 -154.875 ;
        RECT 349.355 -156.565 349.685 -156.235 ;
        RECT 349.355 -157.925 349.685 -157.595 ;
        RECT 349.355 -159.285 349.685 -158.955 ;
        RECT 349.355 -160.645 349.685 -160.315 ;
        RECT 349.355 -162.005 349.685 -161.675 ;
        RECT 349.355 -163.365 349.685 -163.035 ;
        RECT 349.355 -164.725 349.685 -164.395 ;
        RECT 349.355 -166.085 349.685 -165.755 ;
        RECT 349.355 -167.445 349.685 -167.115 ;
        RECT 349.355 -168.805 349.685 -168.475 ;
        RECT 349.355 -170.165 349.685 -169.835 ;
        RECT 349.355 -171.525 349.685 -171.195 ;
        RECT 349.355 -172.885 349.685 -172.555 ;
        RECT 349.355 -174.245 349.685 -173.915 ;
        RECT 349.355 -175.605 349.685 -175.275 ;
        RECT 349.355 -176.965 349.685 -176.635 ;
        RECT 349.355 -178.325 349.685 -177.995 ;
        RECT 349.355 -180.57 349.685 -179.44 ;
        RECT 349.36 -180.685 349.68 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 350.715 241.32 351.045 242.45 ;
        RECT 350.715 239.195 351.045 239.525 ;
        RECT 350.715 237.835 351.045 238.165 ;
        RECT 350.72 237.16 351.04 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 350.715 -95.365 351.045 -95.035 ;
        RECT 350.715 -96.725 351.045 -96.395 ;
        RECT 350.715 -98.085 351.045 -97.755 ;
        RECT 350.715 -99.445 351.045 -99.115 ;
        RECT 350.715 -100.805 351.045 -100.475 ;
        RECT 350.715 -102.165 351.045 -101.835 ;
        RECT 350.715 -103.525 351.045 -103.195 ;
        RECT 350.715 -104.885 351.045 -104.555 ;
        RECT 350.715 -106.245 351.045 -105.915 ;
        RECT 350.715 -107.605 351.045 -107.275 ;
        RECT 350.715 -108.965 351.045 -108.635 ;
        RECT 350.715 -110.325 351.045 -109.995 ;
        RECT 350.715 -111.685 351.045 -111.355 ;
        RECT 350.715 -113.045 351.045 -112.715 ;
        RECT 350.715 -114.405 351.045 -114.075 ;
        RECT 350.715 -115.765 351.045 -115.435 ;
        RECT 350.715 -117.125 351.045 -116.795 ;
        RECT 350.715 -118.485 351.045 -118.155 ;
        RECT 350.715 -119.845 351.045 -119.515 ;
        RECT 350.715 -121.205 351.045 -120.875 ;
        RECT 350.715 -122.565 351.045 -122.235 ;
        RECT 350.715 -123.925 351.045 -123.595 ;
        RECT 350.715 -125.285 351.045 -124.955 ;
        RECT 350.715 -126.645 351.045 -126.315 ;
        RECT 350.715 -128.005 351.045 -127.675 ;
        RECT 350.715 -129.365 351.045 -129.035 ;
        RECT 350.715 -130.725 351.045 -130.395 ;
        RECT 350.715 -132.085 351.045 -131.755 ;
        RECT 350.715 -133.445 351.045 -133.115 ;
        RECT 350.715 -134.805 351.045 -134.475 ;
        RECT 350.715 -136.165 351.045 -135.835 ;
        RECT 350.715 -137.525 351.045 -137.195 ;
        RECT 350.715 -138.885 351.045 -138.555 ;
        RECT 350.715 -140.245 351.045 -139.915 ;
        RECT 350.715 -141.605 351.045 -141.275 ;
        RECT 350.715 -142.965 351.045 -142.635 ;
        RECT 350.715 -144.325 351.045 -143.995 ;
        RECT 350.715 -145.685 351.045 -145.355 ;
        RECT 350.715 -147.045 351.045 -146.715 ;
        RECT 350.715 -148.405 351.045 -148.075 ;
        RECT 350.715 -149.765 351.045 -149.435 ;
        RECT 350.715 -151.125 351.045 -150.795 ;
        RECT 350.715 -152.485 351.045 -152.155 ;
        RECT 350.715 -153.845 351.045 -153.515 ;
        RECT 350.715 -155.205 351.045 -154.875 ;
        RECT 350.715 -156.565 351.045 -156.235 ;
        RECT 350.715 -157.925 351.045 -157.595 ;
        RECT 350.715 -159.285 351.045 -158.955 ;
        RECT 350.715 -160.645 351.045 -160.315 ;
        RECT 350.715 -162.005 351.045 -161.675 ;
        RECT 350.715 -163.365 351.045 -163.035 ;
        RECT 350.715 -164.725 351.045 -164.395 ;
        RECT 350.715 -166.085 351.045 -165.755 ;
        RECT 350.715 -167.445 351.045 -167.115 ;
        RECT 350.715 -168.805 351.045 -168.475 ;
        RECT 350.715 -170.165 351.045 -169.835 ;
        RECT 350.715 -171.525 351.045 -171.195 ;
        RECT 350.715 -172.885 351.045 -172.555 ;
        RECT 350.715 -174.245 351.045 -173.915 ;
        RECT 350.715 -175.605 351.045 -175.275 ;
        RECT 350.715 -176.965 351.045 -176.635 ;
        RECT 350.715 -178.325 351.045 -177.995 ;
        RECT 350.715 -180.57 351.045 -179.44 ;
        RECT 350.72 -180.685 351.04 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 351.01 -94.075 351.34 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 352.075 241.32 352.405 242.45 ;
        RECT 352.075 239.195 352.405 239.525 ;
        RECT 352.075 237.835 352.405 238.165 ;
        RECT 352.08 237.16 352.4 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 352.075 -1.525 352.405 -1.195 ;
        RECT 352.075 -2.885 352.405 -2.555 ;
        RECT 352.08 -3.56 352.4 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 353.435 241.32 353.765 242.45 ;
        RECT 353.435 239.195 353.765 239.525 ;
        RECT 353.435 237.835 353.765 238.165 ;
        RECT 353.44 237.16 353.76 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 353.435 -1.525 353.765 -1.195 ;
        RECT 353.435 -2.885 353.765 -2.555 ;
        RECT 353.44 -3.56 353.76 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 354.795 241.32 355.125 242.45 ;
        RECT 354.795 239.195 355.125 239.525 ;
        RECT 354.795 237.835 355.125 238.165 ;
        RECT 354.8 237.16 355.12 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 354.795 -1.525 355.125 -1.195 ;
        RECT 354.795 -2.885 355.125 -2.555 ;
        RECT 354.8 -3.56 355.12 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 354.795 -91.285 355.125 -90.955 ;
        RECT 354.795 -92.645 355.125 -92.315 ;
        RECT 354.795 -94.005 355.125 -93.675 ;
        RECT 354.795 -95.365 355.125 -95.035 ;
        RECT 354.795 -96.725 355.125 -96.395 ;
        RECT 354.795 -98.085 355.125 -97.755 ;
        RECT 354.795 -99.445 355.125 -99.115 ;
        RECT 354.795 -100.805 355.125 -100.475 ;
        RECT 354.795 -102.165 355.125 -101.835 ;
        RECT 354.795 -103.525 355.125 -103.195 ;
        RECT 354.795 -104.885 355.125 -104.555 ;
        RECT 354.795 -106.245 355.125 -105.915 ;
        RECT 354.795 -107.605 355.125 -107.275 ;
        RECT 354.795 -108.965 355.125 -108.635 ;
        RECT 354.795 -110.325 355.125 -109.995 ;
        RECT 354.795 -111.685 355.125 -111.355 ;
        RECT 354.795 -113.045 355.125 -112.715 ;
        RECT 354.795 -114.405 355.125 -114.075 ;
        RECT 354.795 -115.765 355.125 -115.435 ;
        RECT 354.795 -117.125 355.125 -116.795 ;
        RECT 354.795 -118.485 355.125 -118.155 ;
        RECT 354.795 -119.845 355.125 -119.515 ;
        RECT 354.795 -121.205 355.125 -120.875 ;
        RECT 354.795 -122.565 355.125 -122.235 ;
        RECT 354.795 -123.925 355.125 -123.595 ;
        RECT 354.795 -125.285 355.125 -124.955 ;
        RECT 354.795 -126.645 355.125 -126.315 ;
        RECT 354.795 -128.005 355.125 -127.675 ;
        RECT 354.795 -129.365 355.125 -129.035 ;
        RECT 354.795 -130.725 355.125 -130.395 ;
        RECT 354.795 -132.085 355.125 -131.755 ;
        RECT 354.795 -133.445 355.125 -133.115 ;
        RECT 354.795 -134.805 355.125 -134.475 ;
        RECT 354.795 -136.165 355.125 -135.835 ;
        RECT 354.795 -137.525 355.125 -137.195 ;
        RECT 354.795 -138.885 355.125 -138.555 ;
        RECT 354.795 -140.245 355.125 -139.915 ;
        RECT 354.795 -141.605 355.125 -141.275 ;
        RECT 354.795 -142.965 355.125 -142.635 ;
        RECT 354.795 -144.325 355.125 -143.995 ;
        RECT 354.795 -145.685 355.125 -145.355 ;
        RECT 354.795 -147.045 355.125 -146.715 ;
        RECT 354.795 -148.405 355.125 -148.075 ;
        RECT 354.795 -149.765 355.125 -149.435 ;
        RECT 354.795 -151.125 355.125 -150.795 ;
        RECT 354.795 -152.485 355.125 -152.155 ;
        RECT 354.795 -153.845 355.125 -153.515 ;
        RECT 354.795 -155.205 355.125 -154.875 ;
        RECT 354.795 -156.565 355.125 -156.235 ;
        RECT 354.795 -157.925 355.125 -157.595 ;
        RECT 354.795 -159.285 355.125 -158.955 ;
        RECT 354.795 -160.645 355.125 -160.315 ;
        RECT 354.795 -162.005 355.125 -161.675 ;
        RECT 354.795 -163.365 355.125 -163.035 ;
        RECT 354.795 -164.725 355.125 -164.395 ;
        RECT 354.795 -166.085 355.125 -165.755 ;
        RECT 354.795 -167.445 355.125 -167.115 ;
        RECT 354.795 -168.805 355.125 -168.475 ;
        RECT 354.795 -170.165 355.125 -169.835 ;
        RECT 354.795 -171.525 355.125 -171.195 ;
        RECT 354.795 -172.885 355.125 -172.555 ;
        RECT 354.795 -174.245 355.125 -173.915 ;
        RECT 354.795 -175.605 355.125 -175.275 ;
        RECT 354.795 -176.965 355.125 -176.635 ;
        RECT 354.795 -178.325 355.125 -177.995 ;
        RECT 354.795 -180.57 355.125 -179.44 ;
        RECT 354.8 -180.685 355.12 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 356.155 241.32 356.485 242.45 ;
        RECT 356.155 239.195 356.485 239.525 ;
        RECT 356.155 237.835 356.485 238.165 ;
        RECT 356.16 237.16 356.48 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 356.155 -95.365 356.485 -95.035 ;
        RECT 356.155 -96.725 356.485 -96.395 ;
        RECT 356.155 -98.085 356.485 -97.755 ;
        RECT 356.155 -99.445 356.485 -99.115 ;
        RECT 356.155 -100.805 356.485 -100.475 ;
        RECT 356.155 -102.165 356.485 -101.835 ;
        RECT 356.155 -103.525 356.485 -103.195 ;
        RECT 356.155 -104.885 356.485 -104.555 ;
        RECT 356.155 -106.245 356.485 -105.915 ;
        RECT 356.155 -107.605 356.485 -107.275 ;
        RECT 356.155 -108.965 356.485 -108.635 ;
        RECT 356.155 -110.325 356.485 -109.995 ;
        RECT 356.155 -111.685 356.485 -111.355 ;
        RECT 356.155 -113.045 356.485 -112.715 ;
        RECT 356.155 -114.405 356.485 -114.075 ;
        RECT 356.155 -115.765 356.485 -115.435 ;
        RECT 356.155 -117.125 356.485 -116.795 ;
        RECT 356.155 -118.485 356.485 -118.155 ;
        RECT 356.155 -119.845 356.485 -119.515 ;
        RECT 356.155 -121.205 356.485 -120.875 ;
        RECT 356.155 -122.565 356.485 -122.235 ;
        RECT 356.155 -123.925 356.485 -123.595 ;
        RECT 356.155 -125.285 356.485 -124.955 ;
        RECT 356.155 -126.645 356.485 -126.315 ;
        RECT 356.155 -128.005 356.485 -127.675 ;
        RECT 356.155 -129.365 356.485 -129.035 ;
        RECT 356.155 -130.725 356.485 -130.395 ;
        RECT 356.155 -132.085 356.485 -131.755 ;
        RECT 356.155 -133.445 356.485 -133.115 ;
        RECT 356.155 -134.805 356.485 -134.475 ;
        RECT 356.155 -136.165 356.485 -135.835 ;
        RECT 356.155 -137.525 356.485 -137.195 ;
        RECT 356.155 -138.885 356.485 -138.555 ;
        RECT 356.155 -140.245 356.485 -139.915 ;
        RECT 356.155 -141.605 356.485 -141.275 ;
        RECT 356.155 -142.965 356.485 -142.635 ;
        RECT 356.155 -144.325 356.485 -143.995 ;
        RECT 356.155 -145.685 356.485 -145.355 ;
        RECT 356.155 -147.045 356.485 -146.715 ;
        RECT 356.155 -148.405 356.485 -148.075 ;
        RECT 356.155 -149.765 356.485 -149.435 ;
        RECT 356.155 -151.125 356.485 -150.795 ;
        RECT 356.155 -152.485 356.485 -152.155 ;
        RECT 356.155 -153.845 356.485 -153.515 ;
        RECT 356.155 -155.205 356.485 -154.875 ;
        RECT 356.155 -156.565 356.485 -156.235 ;
        RECT 356.155 -157.925 356.485 -157.595 ;
        RECT 356.155 -159.285 356.485 -158.955 ;
        RECT 356.155 -160.645 356.485 -160.315 ;
        RECT 356.155 -162.005 356.485 -161.675 ;
        RECT 356.155 -163.365 356.485 -163.035 ;
        RECT 356.155 -164.725 356.485 -164.395 ;
        RECT 356.155 -166.085 356.485 -165.755 ;
        RECT 356.155 -167.445 356.485 -167.115 ;
        RECT 356.155 -168.805 356.485 -168.475 ;
        RECT 356.155 -170.165 356.485 -169.835 ;
        RECT 356.155 -171.525 356.485 -171.195 ;
        RECT 356.155 -172.885 356.485 -172.555 ;
        RECT 356.155 -174.245 356.485 -173.915 ;
        RECT 356.155 -175.605 356.485 -175.275 ;
        RECT 356.155 -176.965 356.485 -176.635 ;
        RECT 356.155 -178.325 356.485 -177.995 ;
        RECT 356.155 -180.57 356.485 -179.44 ;
        RECT 356.16 -180.685 356.48 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 357.11 -94.075 357.44 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 357.515 241.32 357.845 242.45 ;
        RECT 357.515 239.195 357.845 239.525 ;
        RECT 357.515 237.835 357.845 238.165 ;
        RECT 357.52 237.16 357.84 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 358.875 241.32 359.205 242.45 ;
        RECT 358.875 239.195 359.205 239.525 ;
        RECT 358.875 237.835 359.205 238.165 ;
        RECT 358.88 237.16 359.2 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 358.875 -1.525 359.205 -1.195 ;
        RECT 358.875 -2.885 359.205 -2.555 ;
        RECT 358.88 -3.56 359.2 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 360.235 241.32 360.565 242.45 ;
        RECT 360.235 239.195 360.565 239.525 ;
        RECT 360.235 237.835 360.565 238.165 ;
        RECT 360.24 237.16 360.56 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 360.235 -1.525 360.565 -1.195 ;
        RECT 360.235 -2.885 360.565 -2.555 ;
        RECT 360.24 -3.56 360.56 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 360.235 -91.285 360.565 -90.955 ;
        RECT 360.235 -92.645 360.565 -92.315 ;
        RECT 360.235 -94.005 360.565 -93.675 ;
        RECT 360.235 -95.365 360.565 -95.035 ;
        RECT 360.235 -96.725 360.565 -96.395 ;
        RECT 360.235 -98.085 360.565 -97.755 ;
        RECT 360.235 -99.445 360.565 -99.115 ;
        RECT 360.235 -100.805 360.565 -100.475 ;
        RECT 360.235 -102.165 360.565 -101.835 ;
        RECT 360.235 -103.525 360.565 -103.195 ;
        RECT 360.235 -104.885 360.565 -104.555 ;
        RECT 360.235 -106.245 360.565 -105.915 ;
        RECT 360.235 -107.605 360.565 -107.275 ;
        RECT 360.235 -108.965 360.565 -108.635 ;
        RECT 360.235 -110.325 360.565 -109.995 ;
        RECT 360.235 -111.685 360.565 -111.355 ;
        RECT 360.235 -113.045 360.565 -112.715 ;
        RECT 360.235 -114.405 360.565 -114.075 ;
        RECT 360.235 -115.765 360.565 -115.435 ;
        RECT 360.235 -117.125 360.565 -116.795 ;
        RECT 360.235 -118.485 360.565 -118.155 ;
        RECT 360.235 -119.845 360.565 -119.515 ;
        RECT 360.235 -121.205 360.565 -120.875 ;
        RECT 360.235 -122.565 360.565 -122.235 ;
        RECT 360.235 -123.925 360.565 -123.595 ;
        RECT 360.235 -125.285 360.565 -124.955 ;
        RECT 360.235 -126.645 360.565 -126.315 ;
        RECT 360.235 -128.005 360.565 -127.675 ;
        RECT 360.235 -129.365 360.565 -129.035 ;
        RECT 360.235 -130.725 360.565 -130.395 ;
        RECT 360.235 -132.085 360.565 -131.755 ;
        RECT 360.235 -133.445 360.565 -133.115 ;
        RECT 360.235 -134.805 360.565 -134.475 ;
        RECT 360.235 -136.165 360.565 -135.835 ;
        RECT 360.235 -137.525 360.565 -137.195 ;
        RECT 360.235 -138.885 360.565 -138.555 ;
        RECT 360.235 -140.245 360.565 -139.915 ;
        RECT 360.235 -141.605 360.565 -141.275 ;
        RECT 360.235 -142.965 360.565 -142.635 ;
        RECT 360.235 -144.325 360.565 -143.995 ;
        RECT 360.235 -145.685 360.565 -145.355 ;
        RECT 360.235 -147.045 360.565 -146.715 ;
        RECT 360.235 -148.405 360.565 -148.075 ;
        RECT 360.235 -149.765 360.565 -149.435 ;
        RECT 360.235 -151.125 360.565 -150.795 ;
        RECT 360.235 -152.485 360.565 -152.155 ;
        RECT 360.235 -153.845 360.565 -153.515 ;
        RECT 360.235 -155.205 360.565 -154.875 ;
        RECT 360.235 -156.565 360.565 -156.235 ;
        RECT 360.235 -157.925 360.565 -157.595 ;
        RECT 360.235 -159.285 360.565 -158.955 ;
        RECT 360.235 -160.645 360.565 -160.315 ;
        RECT 360.235 -162.005 360.565 -161.675 ;
        RECT 360.235 -163.365 360.565 -163.035 ;
        RECT 360.235 -164.725 360.565 -164.395 ;
        RECT 360.235 -166.085 360.565 -165.755 ;
        RECT 360.235 -167.445 360.565 -167.115 ;
        RECT 360.235 -168.805 360.565 -168.475 ;
        RECT 360.235 -170.165 360.565 -169.835 ;
        RECT 360.235 -171.525 360.565 -171.195 ;
        RECT 360.235 -172.885 360.565 -172.555 ;
        RECT 360.235 -174.245 360.565 -173.915 ;
        RECT 360.235 -175.605 360.565 -175.275 ;
        RECT 360.235 -176.965 360.565 -176.635 ;
        RECT 360.235 -178.325 360.565 -177.995 ;
        RECT 360.235 -180.57 360.565 -179.44 ;
        RECT 360.24 -180.685 360.56 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 361.595 241.32 361.925 242.45 ;
        RECT 361.595 239.195 361.925 239.525 ;
        RECT 361.595 237.835 361.925 238.165 ;
        RECT 361.6 237.16 361.92 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 361.595 -1.525 361.925 -1.195 ;
        RECT 361.595 -2.885 361.925 -2.555 ;
        RECT 361.6 -3.56 361.92 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 361.595 -91.285 361.925 -90.955 ;
        RECT 361.595 -92.645 361.925 -92.315 ;
        RECT 361.595 -94.005 361.925 -93.675 ;
        RECT 361.595 -95.365 361.925 -95.035 ;
        RECT 361.595 -96.725 361.925 -96.395 ;
        RECT 361.595 -98.085 361.925 -97.755 ;
        RECT 361.595 -99.445 361.925 -99.115 ;
        RECT 361.595 -100.805 361.925 -100.475 ;
        RECT 361.595 -102.165 361.925 -101.835 ;
        RECT 361.595 -103.525 361.925 -103.195 ;
        RECT 361.595 -104.885 361.925 -104.555 ;
        RECT 361.595 -106.245 361.925 -105.915 ;
        RECT 361.595 -107.605 361.925 -107.275 ;
        RECT 361.595 -108.965 361.925 -108.635 ;
        RECT 361.595 -110.325 361.925 -109.995 ;
        RECT 361.595 -111.685 361.925 -111.355 ;
        RECT 361.595 -113.045 361.925 -112.715 ;
        RECT 361.595 -114.405 361.925 -114.075 ;
        RECT 361.595 -115.765 361.925 -115.435 ;
        RECT 361.595 -117.125 361.925 -116.795 ;
        RECT 361.595 -118.485 361.925 -118.155 ;
        RECT 361.595 -119.845 361.925 -119.515 ;
        RECT 361.595 -121.205 361.925 -120.875 ;
        RECT 361.595 -122.565 361.925 -122.235 ;
        RECT 361.595 -123.925 361.925 -123.595 ;
        RECT 361.595 -125.285 361.925 -124.955 ;
        RECT 361.595 -126.645 361.925 -126.315 ;
        RECT 361.595 -128.005 361.925 -127.675 ;
        RECT 361.595 -129.365 361.925 -129.035 ;
        RECT 361.595 -130.725 361.925 -130.395 ;
        RECT 361.595 -132.085 361.925 -131.755 ;
        RECT 361.595 -133.445 361.925 -133.115 ;
        RECT 361.595 -134.805 361.925 -134.475 ;
        RECT 361.595 -136.165 361.925 -135.835 ;
        RECT 361.595 -137.525 361.925 -137.195 ;
        RECT 361.595 -138.885 361.925 -138.555 ;
        RECT 361.595 -140.245 361.925 -139.915 ;
        RECT 361.595 -141.605 361.925 -141.275 ;
        RECT 361.595 -142.965 361.925 -142.635 ;
        RECT 361.595 -144.325 361.925 -143.995 ;
        RECT 361.595 -145.685 361.925 -145.355 ;
        RECT 361.595 -147.045 361.925 -146.715 ;
        RECT 361.595 -148.405 361.925 -148.075 ;
        RECT 361.595 -149.765 361.925 -149.435 ;
        RECT 361.595 -151.125 361.925 -150.795 ;
        RECT 361.595 -152.485 361.925 -152.155 ;
        RECT 361.595 -153.845 361.925 -153.515 ;
        RECT 361.595 -155.205 361.925 -154.875 ;
        RECT 361.595 -156.565 361.925 -156.235 ;
        RECT 361.595 -157.925 361.925 -157.595 ;
        RECT 361.595 -159.285 361.925 -158.955 ;
        RECT 361.595 -160.645 361.925 -160.315 ;
        RECT 361.595 -162.005 361.925 -161.675 ;
        RECT 361.595 -163.365 361.925 -163.035 ;
        RECT 361.595 -164.725 361.925 -164.395 ;
        RECT 361.595 -166.085 361.925 -165.755 ;
        RECT 361.595 -167.445 361.925 -167.115 ;
        RECT 361.595 -168.805 361.925 -168.475 ;
        RECT 361.595 -170.165 361.925 -169.835 ;
        RECT 361.595 -171.525 361.925 -171.195 ;
        RECT 361.595 -172.885 361.925 -172.555 ;
        RECT 361.595 -174.245 361.925 -173.915 ;
        RECT 361.595 -175.605 361.925 -175.275 ;
        RECT 361.595 -176.965 361.925 -176.635 ;
        RECT 361.595 -178.325 361.925 -177.995 ;
        RECT 361.595 -180.57 361.925 -179.44 ;
        RECT 361.6 -180.685 361.92 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 362.955 241.32 363.285 242.45 ;
        RECT 362.955 239.195 363.285 239.525 ;
        RECT 362.955 237.835 363.285 238.165 ;
        RECT 362.96 237.16 363.28 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 362.955 -95.365 363.285 -95.035 ;
        RECT 362.955 -96.725 363.285 -96.395 ;
        RECT 362.955 -98.085 363.285 -97.755 ;
        RECT 362.955 -99.445 363.285 -99.115 ;
        RECT 362.955 -100.805 363.285 -100.475 ;
        RECT 362.955 -102.165 363.285 -101.835 ;
        RECT 362.955 -103.525 363.285 -103.195 ;
        RECT 362.955 -104.885 363.285 -104.555 ;
        RECT 362.955 -106.245 363.285 -105.915 ;
        RECT 362.955 -107.605 363.285 -107.275 ;
        RECT 362.955 -108.965 363.285 -108.635 ;
        RECT 362.955 -110.325 363.285 -109.995 ;
        RECT 362.955 -111.685 363.285 -111.355 ;
        RECT 362.955 -113.045 363.285 -112.715 ;
        RECT 362.955 -114.405 363.285 -114.075 ;
        RECT 362.955 -115.765 363.285 -115.435 ;
        RECT 362.955 -117.125 363.285 -116.795 ;
        RECT 362.955 -118.485 363.285 -118.155 ;
        RECT 362.955 -119.845 363.285 -119.515 ;
        RECT 362.955 -121.205 363.285 -120.875 ;
        RECT 362.955 -122.565 363.285 -122.235 ;
        RECT 362.955 -123.925 363.285 -123.595 ;
        RECT 362.955 -125.285 363.285 -124.955 ;
        RECT 362.955 -126.645 363.285 -126.315 ;
        RECT 362.955 -128.005 363.285 -127.675 ;
        RECT 362.955 -129.365 363.285 -129.035 ;
        RECT 362.955 -130.725 363.285 -130.395 ;
        RECT 362.955 -132.085 363.285 -131.755 ;
        RECT 362.955 -133.445 363.285 -133.115 ;
        RECT 362.955 -134.805 363.285 -134.475 ;
        RECT 362.955 -136.165 363.285 -135.835 ;
        RECT 362.955 -137.525 363.285 -137.195 ;
        RECT 362.955 -138.885 363.285 -138.555 ;
        RECT 362.955 -140.245 363.285 -139.915 ;
        RECT 362.955 -141.605 363.285 -141.275 ;
        RECT 362.955 -142.965 363.285 -142.635 ;
        RECT 362.955 -144.325 363.285 -143.995 ;
        RECT 362.955 -145.685 363.285 -145.355 ;
        RECT 362.955 -147.045 363.285 -146.715 ;
        RECT 362.955 -148.405 363.285 -148.075 ;
        RECT 362.955 -149.765 363.285 -149.435 ;
        RECT 362.955 -151.125 363.285 -150.795 ;
        RECT 362.955 -152.485 363.285 -152.155 ;
        RECT 362.955 -153.845 363.285 -153.515 ;
        RECT 362.955 -155.205 363.285 -154.875 ;
        RECT 362.955 -156.565 363.285 -156.235 ;
        RECT 362.955 -157.925 363.285 -157.595 ;
        RECT 362.955 -159.285 363.285 -158.955 ;
        RECT 362.955 -160.645 363.285 -160.315 ;
        RECT 362.955 -162.005 363.285 -161.675 ;
        RECT 362.955 -163.365 363.285 -163.035 ;
        RECT 362.955 -164.725 363.285 -164.395 ;
        RECT 362.955 -166.085 363.285 -165.755 ;
        RECT 362.955 -167.445 363.285 -167.115 ;
        RECT 362.955 -168.805 363.285 -168.475 ;
        RECT 362.955 -170.165 363.285 -169.835 ;
        RECT 362.955 -171.525 363.285 -171.195 ;
        RECT 362.955 -172.885 363.285 -172.555 ;
        RECT 362.955 -174.245 363.285 -173.915 ;
        RECT 362.955 -175.605 363.285 -175.275 ;
        RECT 362.955 -176.965 363.285 -176.635 ;
        RECT 362.955 -178.325 363.285 -177.995 ;
        RECT 362.955 -180.57 363.285 -179.44 ;
        RECT 362.96 -180.685 363.28 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 363.21 -94.075 363.54 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 364.315 241.32 364.645 242.45 ;
        RECT 364.315 239.195 364.645 239.525 ;
        RECT 364.315 237.835 364.645 238.165 ;
        RECT 364.32 237.16 364.64 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 364.315 -1.525 364.645 -1.195 ;
        RECT 364.315 -2.885 364.645 -2.555 ;
        RECT 364.32 -3.56 364.64 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 365.675 241.32 366.005 242.45 ;
        RECT 365.675 239.195 366.005 239.525 ;
        RECT 365.675 237.835 366.005 238.165 ;
        RECT 365.68 237.16 366 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 365.675 -1.525 366.005 -1.195 ;
        RECT 365.675 -2.885 366.005 -2.555 ;
        RECT 365.68 -3.56 366 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 367.035 241.32 367.365 242.45 ;
        RECT 367.035 239.195 367.365 239.525 ;
        RECT 367.035 237.835 367.365 238.165 ;
        RECT 367.04 237.16 367.36 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 367.035 -1.525 367.365 -1.195 ;
        RECT 367.035 -2.885 367.365 -2.555 ;
        RECT 367.04 -3.56 367.36 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 367.035 -91.285 367.365 -90.955 ;
        RECT 367.035 -92.645 367.365 -92.315 ;
        RECT 367.035 -94.005 367.365 -93.675 ;
        RECT 367.035 -95.365 367.365 -95.035 ;
        RECT 367.035 -96.725 367.365 -96.395 ;
        RECT 367.035 -98.085 367.365 -97.755 ;
        RECT 367.035 -99.445 367.365 -99.115 ;
        RECT 367.035 -100.805 367.365 -100.475 ;
        RECT 367.035 -102.165 367.365 -101.835 ;
        RECT 367.035 -103.525 367.365 -103.195 ;
        RECT 367.035 -104.885 367.365 -104.555 ;
        RECT 367.035 -106.245 367.365 -105.915 ;
        RECT 367.035 -107.605 367.365 -107.275 ;
        RECT 367.035 -108.965 367.365 -108.635 ;
        RECT 367.035 -110.325 367.365 -109.995 ;
        RECT 367.035 -111.685 367.365 -111.355 ;
        RECT 367.035 -113.045 367.365 -112.715 ;
        RECT 367.035 -114.405 367.365 -114.075 ;
        RECT 367.035 -115.765 367.365 -115.435 ;
        RECT 367.035 -117.125 367.365 -116.795 ;
        RECT 367.035 -118.485 367.365 -118.155 ;
        RECT 367.035 -119.845 367.365 -119.515 ;
        RECT 367.035 -121.205 367.365 -120.875 ;
        RECT 367.035 -122.565 367.365 -122.235 ;
        RECT 367.035 -123.925 367.365 -123.595 ;
        RECT 367.035 -125.285 367.365 -124.955 ;
        RECT 367.035 -126.645 367.365 -126.315 ;
        RECT 367.035 -128.005 367.365 -127.675 ;
        RECT 367.035 -129.365 367.365 -129.035 ;
        RECT 367.035 -130.725 367.365 -130.395 ;
        RECT 367.035 -132.085 367.365 -131.755 ;
        RECT 367.035 -133.445 367.365 -133.115 ;
        RECT 367.035 -134.805 367.365 -134.475 ;
        RECT 367.035 -136.165 367.365 -135.835 ;
        RECT 367.035 -137.525 367.365 -137.195 ;
        RECT 367.035 -138.885 367.365 -138.555 ;
        RECT 367.035 -140.245 367.365 -139.915 ;
        RECT 367.035 -141.605 367.365 -141.275 ;
        RECT 367.035 -142.965 367.365 -142.635 ;
        RECT 367.035 -144.325 367.365 -143.995 ;
        RECT 367.035 -145.685 367.365 -145.355 ;
        RECT 367.035 -147.045 367.365 -146.715 ;
        RECT 367.035 -148.405 367.365 -148.075 ;
        RECT 367.035 -149.765 367.365 -149.435 ;
        RECT 367.035 -151.125 367.365 -150.795 ;
        RECT 367.035 -152.485 367.365 -152.155 ;
        RECT 367.035 -153.845 367.365 -153.515 ;
        RECT 367.035 -155.205 367.365 -154.875 ;
        RECT 367.035 -156.565 367.365 -156.235 ;
        RECT 367.035 -157.925 367.365 -157.595 ;
        RECT 367.035 -159.285 367.365 -158.955 ;
        RECT 367.035 -160.645 367.365 -160.315 ;
        RECT 367.035 -162.005 367.365 -161.675 ;
        RECT 367.035 -163.365 367.365 -163.035 ;
        RECT 367.035 -164.725 367.365 -164.395 ;
        RECT 367.035 -166.085 367.365 -165.755 ;
        RECT 367.035 -167.445 367.365 -167.115 ;
        RECT 367.035 -168.805 367.365 -168.475 ;
        RECT 367.035 -170.165 367.365 -169.835 ;
        RECT 367.035 -171.525 367.365 -171.195 ;
        RECT 367.035 -172.885 367.365 -172.555 ;
        RECT 367.035 -174.245 367.365 -173.915 ;
        RECT 367.035 -175.605 367.365 -175.275 ;
        RECT 367.035 -176.965 367.365 -176.635 ;
        RECT 367.035 -178.325 367.365 -177.995 ;
        RECT 367.035 -180.57 367.365 -179.44 ;
        RECT 367.04 -180.685 367.36 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 368.395 241.32 368.725 242.45 ;
        RECT 368.395 239.195 368.725 239.525 ;
        RECT 368.395 237.835 368.725 238.165 ;
        RECT 368.4 237.16 368.72 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 368.395 -125.285 368.725 -124.955 ;
        RECT 368.395 -126.645 368.725 -126.315 ;
        RECT 368.395 -128.005 368.725 -127.675 ;
        RECT 368.395 -129.365 368.725 -129.035 ;
        RECT 368.395 -130.725 368.725 -130.395 ;
        RECT 368.395 -132.085 368.725 -131.755 ;
        RECT 368.395 -133.445 368.725 -133.115 ;
        RECT 368.395 -134.805 368.725 -134.475 ;
        RECT 368.395 -136.165 368.725 -135.835 ;
        RECT 368.395 -137.525 368.725 -137.195 ;
        RECT 368.395 -138.885 368.725 -138.555 ;
        RECT 368.395 -140.245 368.725 -139.915 ;
        RECT 368.395 -141.605 368.725 -141.275 ;
        RECT 368.395 -142.965 368.725 -142.635 ;
        RECT 368.395 -144.325 368.725 -143.995 ;
        RECT 368.395 -145.685 368.725 -145.355 ;
        RECT 368.395 -147.045 368.725 -146.715 ;
        RECT 368.395 -148.405 368.725 -148.075 ;
        RECT 368.395 -149.765 368.725 -149.435 ;
        RECT 368.395 -151.125 368.725 -150.795 ;
        RECT 368.395 -152.485 368.725 -152.155 ;
        RECT 368.395 -153.845 368.725 -153.515 ;
        RECT 368.395 -155.205 368.725 -154.875 ;
        RECT 368.395 -156.565 368.725 -156.235 ;
        RECT 368.395 -157.925 368.725 -157.595 ;
        RECT 368.395 -159.285 368.725 -158.955 ;
        RECT 368.395 -160.645 368.725 -160.315 ;
        RECT 368.395 -162.005 368.725 -161.675 ;
        RECT 368.395 -163.365 368.725 -163.035 ;
        RECT 368.395 -164.725 368.725 -164.395 ;
        RECT 368.395 -166.085 368.725 -165.755 ;
        RECT 368.395 -167.445 368.725 -167.115 ;
        RECT 368.395 -168.805 368.725 -168.475 ;
        RECT 368.395 -170.165 368.725 -169.835 ;
        RECT 368.395 -171.525 368.725 -171.195 ;
        RECT 368.395 -172.885 368.725 -172.555 ;
        RECT 368.395 -174.245 368.725 -173.915 ;
        RECT 368.395 -175.605 368.725 -175.275 ;
        RECT 368.395 -176.965 368.725 -176.635 ;
        RECT 368.395 -178.325 368.725 -177.995 ;
        RECT 368.395 -180.57 368.725 -179.44 ;
        RECT 368.4 -180.685 368.72 -95.035 ;
        RECT 368.395 -95.365 368.725 -95.035 ;
        RECT 368.395 -96.725 368.725 -96.395 ;
        RECT 368.395 -98.085 368.725 -97.755 ;
        RECT 368.395 -99.445 368.725 -99.115 ;
        RECT 368.395 -100.805 368.725 -100.475 ;
        RECT 368.395 -102.165 368.725 -101.835 ;
        RECT 368.395 -103.525 368.725 -103.195 ;
        RECT 368.395 -104.885 368.725 -104.555 ;
        RECT 368.395 -106.245 368.725 -105.915 ;
        RECT 368.395 -107.605 368.725 -107.275 ;
        RECT 368.395 -108.965 368.725 -108.635 ;
        RECT 368.395 -110.325 368.725 -109.995 ;
        RECT 368.395 -111.685 368.725 -111.355 ;
        RECT 368.395 -113.045 368.725 -112.715 ;
        RECT 368.395 -114.405 368.725 -114.075 ;
        RECT 368.395 -115.765 368.725 -115.435 ;
        RECT 368.395 -117.125 368.725 -116.795 ;
        RECT 368.395 -118.485 368.725 -118.155 ;
        RECT 368.395 -119.845 368.725 -119.515 ;
        RECT 368.395 -121.205 368.725 -120.875 ;
        RECT 368.395 -122.565 368.725 -122.235 ;
        RECT 368.395 -123.925 368.725 -123.595 ;
    END
    PORT
      LAYER met3 ;
        RECT 301.755 241.32 302.085 242.45 ;
        RECT 301.755 239.195 302.085 239.525 ;
        RECT 301.755 237.835 302.085 238.165 ;
        RECT 301.76 237.16 302.08 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 301.755 -95.365 302.085 -95.035 ;
        RECT 301.755 -96.725 302.085 -96.395 ;
        RECT 301.755 -98.085 302.085 -97.755 ;
        RECT 301.755 -99.445 302.085 -99.115 ;
        RECT 301.755 -100.805 302.085 -100.475 ;
        RECT 301.755 -102.165 302.085 -101.835 ;
        RECT 301.755 -103.525 302.085 -103.195 ;
        RECT 301.755 -104.885 302.085 -104.555 ;
        RECT 301.755 -106.245 302.085 -105.915 ;
        RECT 301.755 -107.605 302.085 -107.275 ;
        RECT 301.755 -108.965 302.085 -108.635 ;
        RECT 301.755 -110.325 302.085 -109.995 ;
        RECT 301.755 -111.685 302.085 -111.355 ;
        RECT 301.755 -113.045 302.085 -112.715 ;
        RECT 301.755 -114.405 302.085 -114.075 ;
        RECT 301.755 -115.765 302.085 -115.435 ;
        RECT 301.755 -117.125 302.085 -116.795 ;
        RECT 301.755 -118.485 302.085 -118.155 ;
        RECT 301.755 -119.845 302.085 -119.515 ;
        RECT 301.755 -121.205 302.085 -120.875 ;
        RECT 301.755 -122.565 302.085 -122.235 ;
        RECT 301.755 -123.925 302.085 -123.595 ;
        RECT 301.755 -125.285 302.085 -124.955 ;
        RECT 301.755 -126.645 302.085 -126.315 ;
        RECT 301.755 -128.005 302.085 -127.675 ;
        RECT 301.755 -129.365 302.085 -129.035 ;
        RECT 301.755 -130.725 302.085 -130.395 ;
        RECT 301.755 -132.085 302.085 -131.755 ;
        RECT 301.755 -133.445 302.085 -133.115 ;
        RECT 301.755 -134.805 302.085 -134.475 ;
        RECT 301.755 -136.165 302.085 -135.835 ;
        RECT 301.755 -137.525 302.085 -137.195 ;
        RECT 301.755 -138.885 302.085 -138.555 ;
        RECT 301.755 -140.245 302.085 -139.915 ;
        RECT 301.755 -141.605 302.085 -141.275 ;
        RECT 301.755 -142.965 302.085 -142.635 ;
        RECT 301.755 -144.325 302.085 -143.995 ;
        RECT 301.755 -145.685 302.085 -145.355 ;
        RECT 301.755 -147.045 302.085 -146.715 ;
        RECT 301.755 -148.405 302.085 -148.075 ;
        RECT 301.755 -149.765 302.085 -149.435 ;
        RECT 301.755 -151.125 302.085 -150.795 ;
        RECT 301.755 -152.485 302.085 -152.155 ;
        RECT 301.755 -153.845 302.085 -153.515 ;
        RECT 301.755 -155.205 302.085 -154.875 ;
        RECT 301.755 -156.565 302.085 -156.235 ;
        RECT 301.755 -157.925 302.085 -157.595 ;
        RECT 301.755 -159.285 302.085 -158.955 ;
        RECT 301.755 -160.645 302.085 -160.315 ;
        RECT 301.755 -162.005 302.085 -161.675 ;
        RECT 301.755 -163.365 302.085 -163.035 ;
        RECT 301.755 -164.725 302.085 -164.395 ;
        RECT 301.755 -166.085 302.085 -165.755 ;
        RECT 301.755 -167.445 302.085 -167.115 ;
        RECT 301.755 -168.805 302.085 -168.475 ;
        RECT 301.755 -170.165 302.085 -169.835 ;
        RECT 301.755 -171.525 302.085 -171.195 ;
        RECT 301.755 -172.885 302.085 -172.555 ;
        RECT 301.755 -174.245 302.085 -173.915 ;
        RECT 301.755 -175.605 302.085 -175.275 ;
        RECT 301.755 -176.965 302.085 -176.635 ;
        RECT 301.755 -178.325 302.085 -177.995 ;
        RECT 301.755 -180.57 302.085 -179.44 ;
        RECT 301.76 -180.685 302.08 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 302.21 -94.075 302.54 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 303.115 241.32 303.445 242.45 ;
        RECT 303.115 239.195 303.445 239.525 ;
        RECT 303.115 237.835 303.445 238.165 ;
        RECT 303.12 237.16 303.44 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 303.115 -1.525 303.445 -1.195 ;
        RECT 303.115 -2.885 303.445 -2.555 ;
        RECT 303.12 -3.56 303.44 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 304.475 241.32 304.805 242.45 ;
        RECT 304.475 239.195 304.805 239.525 ;
        RECT 304.475 237.835 304.805 238.165 ;
        RECT 304.48 237.16 304.8 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 304.475 -1.525 304.805 -1.195 ;
        RECT 304.475 -2.885 304.805 -2.555 ;
        RECT 304.48 -3.56 304.8 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 305.835 241.32 306.165 242.45 ;
        RECT 305.835 239.195 306.165 239.525 ;
        RECT 305.835 237.835 306.165 238.165 ;
        RECT 305.84 237.16 306.16 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 305.835 -1.525 306.165 -1.195 ;
        RECT 305.835 -2.885 306.165 -2.555 ;
        RECT 305.84 -3.56 306.16 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 305.835 -91.285 306.165 -90.955 ;
        RECT 305.835 -92.645 306.165 -92.315 ;
        RECT 305.835 -94.005 306.165 -93.675 ;
        RECT 305.835 -95.365 306.165 -95.035 ;
        RECT 305.835 -96.725 306.165 -96.395 ;
        RECT 305.835 -98.085 306.165 -97.755 ;
        RECT 305.835 -99.445 306.165 -99.115 ;
        RECT 305.835 -100.805 306.165 -100.475 ;
        RECT 305.835 -102.165 306.165 -101.835 ;
        RECT 305.835 -103.525 306.165 -103.195 ;
        RECT 305.835 -104.885 306.165 -104.555 ;
        RECT 305.835 -106.245 306.165 -105.915 ;
        RECT 305.835 -107.605 306.165 -107.275 ;
        RECT 305.835 -108.965 306.165 -108.635 ;
        RECT 305.835 -110.325 306.165 -109.995 ;
        RECT 305.835 -111.685 306.165 -111.355 ;
        RECT 305.835 -113.045 306.165 -112.715 ;
        RECT 305.835 -114.405 306.165 -114.075 ;
        RECT 305.835 -115.765 306.165 -115.435 ;
        RECT 305.835 -117.125 306.165 -116.795 ;
        RECT 305.835 -118.485 306.165 -118.155 ;
        RECT 305.835 -119.845 306.165 -119.515 ;
        RECT 305.835 -121.205 306.165 -120.875 ;
        RECT 305.835 -122.565 306.165 -122.235 ;
        RECT 305.835 -123.925 306.165 -123.595 ;
        RECT 305.835 -125.285 306.165 -124.955 ;
        RECT 305.835 -126.645 306.165 -126.315 ;
        RECT 305.835 -128.005 306.165 -127.675 ;
        RECT 305.835 -129.365 306.165 -129.035 ;
        RECT 305.835 -130.725 306.165 -130.395 ;
        RECT 305.835 -132.085 306.165 -131.755 ;
        RECT 305.835 -133.445 306.165 -133.115 ;
        RECT 305.835 -134.805 306.165 -134.475 ;
        RECT 305.835 -136.165 306.165 -135.835 ;
        RECT 305.835 -137.525 306.165 -137.195 ;
        RECT 305.835 -138.885 306.165 -138.555 ;
        RECT 305.835 -140.245 306.165 -139.915 ;
        RECT 305.835 -141.605 306.165 -141.275 ;
        RECT 305.835 -142.965 306.165 -142.635 ;
        RECT 305.835 -144.325 306.165 -143.995 ;
        RECT 305.835 -145.685 306.165 -145.355 ;
        RECT 305.835 -147.045 306.165 -146.715 ;
        RECT 305.835 -148.405 306.165 -148.075 ;
        RECT 305.835 -149.765 306.165 -149.435 ;
        RECT 305.835 -151.125 306.165 -150.795 ;
        RECT 305.835 -152.485 306.165 -152.155 ;
        RECT 305.835 -153.845 306.165 -153.515 ;
        RECT 305.835 -155.205 306.165 -154.875 ;
        RECT 305.835 -156.565 306.165 -156.235 ;
        RECT 305.835 -157.925 306.165 -157.595 ;
        RECT 305.835 -159.285 306.165 -158.955 ;
        RECT 305.835 -160.645 306.165 -160.315 ;
        RECT 305.835 -162.005 306.165 -161.675 ;
        RECT 305.835 -163.365 306.165 -163.035 ;
        RECT 305.835 -164.725 306.165 -164.395 ;
        RECT 305.835 -166.085 306.165 -165.755 ;
        RECT 305.835 -167.445 306.165 -167.115 ;
        RECT 305.835 -168.805 306.165 -168.475 ;
        RECT 305.835 -170.165 306.165 -169.835 ;
        RECT 305.835 -171.525 306.165 -171.195 ;
        RECT 305.835 -172.885 306.165 -172.555 ;
        RECT 305.835 -174.245 306.165 -173.915 ;
        RECT 305.835 -175.605 306.165 -175.275 ;
        RECT 305.835 -176.965 306.165 -176.635 ;
        RECT 305.835 -178.325 306.165 -177.995 ;
        RECT 305.835 -180.57 306.165 -179.44 ;
        RECT 305.84 -180.685 306.16 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 307.195 241.32 307.525 242.45 ;
        RECT 307.195 239.195 307.525 239.525 ;
        RECT 307.195 237.835 307.525 238.165 ;
        RECT 307.2 237.16 307.52 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 307.195 -95.365 307.525 -95.035 ;
        RECT 307.195 -96.725 307.525 -96.395 ;
        RECT 307.195 -98.085 307.525 -97.755 ;
        RECT 307.195 -99.445 307.525 -99.115 ;
        RECT 307.195 -100.805 307.525 -100.475 ;
        RECT 307.195 -102.165 307.525 -101.835 ;
        RECT 307.195 -103.525 307.525 -103.195 ;
        RECT 307.195 -104.885 307.525 -104.555 ;
        RECT 307.195 -106.245 307.525 -105.915 ;
        RECT 307.195 -107.605 307.525 -107.275 ;
        RECT 307.195 -108.965 307.525 -108.635 ;
        RECT 307.195 -110.325 307.525 -109.995 ;
        RECT 307.195 -111.685 307.525 -111.355 ;
        RECT 307.195 -113.045 307.525 -112.715 ;
        RECT 307.195 -114.405 307.525 -114.075 ;
        RECT 307.195 -115.765 307.525 -115.435 ;
        RECT 307.195 -117.125 307.525 -116.795 ;
        RECT 307.195 -118.485 307.525 -118.155 ;
        RECT 307.195 -119.845 307.525 -119.515 ;
        RECT 307.195 -121.205 307.525 -120.875 ;
        RECT 307.195 -122.565 307.525 -122.235 ;
        RECT 307.195 -123.925 307.525 -123.595 ;
        RECT 307.195 -125.285 307.525 -124.955 ;
        RECT 307.195 -126.645 307.525 -126.315 ;
        RECT 307.195 -128.005 307.525 -127.675 ;
        RECT 307.195 -129.365 307.525 -129.035 ;
        RECT 307.195 -130.725 307.525 -130.395 ;
        RECT 307.195 -132.085 307.525 -131.755 ;
        RECT 307.195 -133.445 307.525 -133.115 ;
        RECT 307.195 -134.805 307.525 -134.475 ;
        RECT 307.195 -136.165 307.525 -135.835 ;
        RECT 307.195 -137.525 307.525 -137.195 ;
        RECT 307.195 -138.885 307.525 -138.555 ;
        RECT 307.195 -140.245 307.525 -139.915 ;
        RECT 307.195 -141.605 307.525 -141.275 ;
        RECT 307.195 -142.965 307.525 -142.635 ;
        RECT 307.195 -144.325 307.525 -143.995 ;
        RECT 307.195 -145.685 307.525 -145.355 ;
        RECT 307.195 -147.045 307.525 -146.715 ;
        RECT 307.195 -148.405 307.525 -148.075 ;
        RECT 307.195 -149.765 307.525 -149.435 ;
        RECT 307.195 -151.125 307.525 -150.795 ;
        RECT 307.195 -152.485 307.525 -152.155 ;
        RECT 307.195 -153.845 307.525 -153.515 ;
        RECT 307.195 -155.205 307.525 -154.875 ;
        RECT 307.195 -156.565 307.525 -156.235 ;
        RECT 307.195 -157.925 307.525 -157.595 ;
        RECT 307.195 -159.285 307.525 -158.955 ;
        RECT 307.195 -160.645 307.525 -160.315 ;
        RECT 307.195 -162.005 307.525 -161.675 ;
        RECT 307.195 -163.365 307.525 -163.035 ;
        RECT 307.195 -164.725 307.525 -164.395 ;
        RECT 307.195 -166.085 307.525 -165.755 ;
        RECT 307.195 -167.445 307.525 -167.115 ;
        RECT 307.195 -168.805 307.525 -168.475 ;
        RECT 307.195 -170.165 307.525 -169.835 ;
        RECT 307.195 -171.525 307.525 -171.195 ;
        RECT 307.195 -172.885 307.525 -172.555 ;
        RECT 307.195 -174.245 307.525 -173.915 ;
        RECT 307.195 -175.605 307.525 -175.275 ;
        RECT 307.195 -176.965 307.525 -176.635 ;
        RECT 307.195 -178.325 307.525 -177.995 ;
        RECT 307.195 -180.57 307.525 -179.44 ;
        RECT 307.2 -180.685 307.52 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 308.31 -94.075 308.64 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 308.555 241.32 308.885 242.45 ;
        RECT 308.555 239.195 308.885 239.525 ;
        RECT 308.555 237.835 308.885 238.165 ;
        RECT 308.56 237.16 308.88 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 309.915 241.32 310.245 242.45 ;
        RECT 309.915 239.195 310.245 239.525 ;
        RECT 309.915 237.835 310.245 238.165 ;
        RECT 309.92 237.16 310.24 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 309.915 -1.525 310.245 -1.195 ;
        RECT 309.915 -2.885 310.245 -2.555 ;
        RECT 309.92 -3.56 310.24 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 309.915 -91.285 310.245 -90.955 ;
        RECT 309.915 -92.645 310.245 -92.315 ;
        RECT 309.915 -94.005 310.245 -93.675 ;
        RECT 309.915 -95.365 310.245 -95.035 ;
        RECT 309.915 -96.725 310.245 -96.395 ;
        RECT 309.915 -98.085 310.245 -97.755 ;
        RECT 309.915 -99.445 310.245 -99.115 ;
        RECT 309.915 -100.805 310.245 -100.475 ;
        RECT 309.915 -102.165 310.245 -101.835 ;
        RECT 309.915 -103.525 310.245 -103.195 ;
        RECT 309.915 -104.885 310.245 -104.555 ;
        RECT 309.915 -106.245 310.245 -105.915 ;
        RECT 309.915 -107.605 310.245 -107.275 ;
        RECT 309.915 -108.965 310.245 -108.635 ;
        RECT 309.915 -110.325 310.245 -109.995 ;
        RECT 309.915 -111.685 310.245 -111.355 ;
        RECT 309.915 -113.045 310.245 -112.715 ;
        RECT 309.915 -114.405 310.245 -114.075 ;
        RECT 309.915 -115.765 310.245 -115.435 ;
        RECT 309.915 -117.125 310.245 -116.795 ;
        RECT 309.915 -118.485 310.245 -118.155 ;
        RECT 309.915 -119.845 310.245 -119.515 ;
        RECT 309.915 -121.205 310.245 -120.875 ;
        RECT 309.915 -122.565 310.245 -122.235 ;
        RECT 309.915 -123.925 310.245 -123.595 ;
        RECT 309.915 -125.285 310.245 -124.955 ;
        RECT 309.915 -126.645 310.245 -126.315 ;
        RECT 309.915 -128.005 310.245 -127.675 ;
        RECT 309.915 -129.365 310.245 -129.035 ;
        RECT 309.915 -130.725 310.245 -130.395 ;
        RECT 309.915 -132.085 310.245 -131.755 ;
        RECT 309.915 -133.445 310.245 -133.115 ;
        RECT 309.915 -134.805 310.245 -134.475 ;
        RECT 309.915 -136.165 310.245 -135.835 ;
        RECT 309.915 -137.525 310.245 -137.195 ;
        RECT 309.915 -138.885 310.245 -138.555 ;
        RECT 309.915 -140.245 310.245 -139.915 ;
        RECT 309.915 -141.605 310.245 -141.275 ;
        RECT 309.915 -142.965 310.245 -142.635 ;
        RECT 309.915 -144.325 310.245 -143.995 ;
        RECT 309.915 -145.685 310.245 -145.355 ;
        RECT 309.915 -147.045 310.245 -146.715 ;
        RECT 309.915 -148.405 310.245 -148.075 ;
        RECT 309.915 -149.765 310.245 -149.435 ;
        RECT 309.915 -151.125 310.245 -150.795 ;
        RECT 309.915 -152.485 310.245 -152.155 ;
        RECT 309.915 -153.845 310.245 -153.515 ;
        RECT 309.915 -155.205 310.245 -154.875 ;
        RECT 309.915 -156.565 310.245 -156.235 ;
        RECT 309.915 -157.925 310.245 -157.595 ;
        RECT 309.915 -159.285 310.245 -158.955 ;
        RECT 309.915 -160.645 310.245 -160.315 ;
        RECT 309.915 -162.005 310.245 -161.675 ;
        RECT 309.915 -163.365 310.245 -163.035 ;
        RECT 309.915 -164.725 310.245 -164.395 ;
        RECT 309.915 -166.085 310.245 -165.755 ;
        RECT 309.915 -167.445 310.245 -167.115 ;
        RECT 309.915 -168.805 310.245 -168.475 ;
        RECT 309.915 -170.165 310.245 -169.835 ;
        RECT 309.915 -171.525 310.245 -171.195 ;
        RECT 309.915 -172.885 310.245 -172.555 ;
        RECT 309.915 -174.245 310.245 -173.915 ;
        RECT 309.915 -175.605 310.245 -175.275 ;
        RECT 309.915 -176.965 310.245 -176.635 ;
        RECT 309.915 -178.325 310.245 -177.995 ;
        RECT 309.915 -180.57 310.245 -179.44 ;
        RECT 309.92 -180.685 310.24 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 311.275 241.32 311.605 242.45 ;
        RECT 311.275 239.195 311.605 239.525 ;
        RECT 311.275 237.835 311.605 238.165 ;
        RECT 311.28 237.16 311.6 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 311.275 -1.525 311.605 -1.195 ;
        RECT 311.275 -2.885 311.605 -2.555 ;
        RECT 311.28 -3.56 311.6 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 312.635 241.32 312.965 242.45 ;
        RECT 312.635 239.195 312.965 239.525 ;
        RECT 312.635 237.835 312.965 238.165 ;
        RECT 312.64 237.16 312.96 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 312.635 -1.525 312.965 -1.195 ;
        RECT 312.635 -2.885 312.965 -2.555 ;
        RECT 312.64 -3.56 312.96 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 312.635 -91.285 312.965 -90.955 ;
        RECT 312.635 -92.645 312.965 -92.315 ;
        RECT 312.635 -94.005 312.965 -93.675 ;
        RECT 312.635 -95.365 312.965 -95.035 ;
        RECT 312.635 -96.725 312.965 -96.395 ;
        RECT 312.635 -98.085 312.965 -97.755 ;
        RECT 312.635 -99.445 312.965 -99.115 ;
        RECT 312.635 -100.805 312.965 -100.475 ;
        RECT 312.635 -102.165 312.965 -101.835 ;
        RECT 312.635 -103.525 312.965 -103.195 ;
        RECT 312.635 -104.885 312.965 -104.555 ;
        RECT 312.635 -106.245 312.965 -105.915 ;
        RECT 312.635 -107.605 312.965 -107.275 ;
        RECT 312.635 -108.965 312.965 -108.635 ;
        RECT 312.635 -110.325 312.965 -109.995 ;
        RECT 312.635 -111.685 312.965 -111.355 ;
        RECT 312.635 -113.045 312.965 -112.715 ;
        RECT 312.635 -114.405 312.965 -114.075 ;
        RECT 312.635 -115.765 312.965 -115.435 ;
        RECT 312.635 -117.125 312.965 -116.795 ;
        RECT 312.635 -118.485 312.965 -118.155 ;
        RECT 312.635 -119.845 312.965 -119.515 ;
        RECT 312.635 -121.205 312.965 -120.875 ;
        RECT 312.635 -122.565 312.965 -122.235 ;
        RECT 312.635 -123.925 312.965 -123.595 ;
        RECT 312.635 -125.285 312.965 -124.955 ;
        RECT 312.635 -126.645 312.965 -126.315 ;
        RECT 312.635 -128.005 312.965 -127.675 ;
        RECT 312.635 -129.365 312.965 -129.035 ;
        RECT 312.635 -130.725 312.965 -130.395 ;
        RECT 312.635 -132.085 312.965 -131.755 ;
        RECT 312.635 -133.445 312.965 -133.115 ;
        RECT 312.635 -134.805 312.965 -134.475 ;
        RECT 312.635 -136.165 312.965 -135.835 ;
        RECT 312.635 -137.525 312.965 -137.195 ;
        RECT 312.635 -138.885 312.965 -138.555 ;
        RECT 312.635 -140.245 312.965 -139.915 ;
        RECT 312.635 -141.605 312.965 -141.275 ;
        RECT 312.635 -142.965 312.965 -142.635 ;
        RECT 312.635 -144.325 312.965 -143.995 ;
        RECT 312.635 -145.685 312.965 -145.355 ;
        RECT 312.635 -147.045 312.965 -146.715 ;
        RECT 312.635 -148.405 312.965 -148.075 ;
        RECT 312.635 -149.765 312.965 -149.435 ;
        RECT 312.635 -151.125 312.965 -150.795 ;
        RECT 312.635 -152.485 312.965 -152.155 ;
        RECT 312.635 -153.845 312.965 -153.515 ;
        RECT 312.635 -155.205 312.965 -154.875 ;
        RECT 312.635 -156.565 312.965 -156.235 ;
        RECT 312.635 -157.925 312.965 -157.595 ;
        RECT 312.635 -159.285 312.965 -158.955 ;
        RECT 312.635 -160.645 312.965 -160.315 ;
        RECT 312.635 -162.005 312.965 -161.675 ;
        RECT 312.635 -163.365 312.965 -163.035 ;
        RECT 312.635 -164.725 312.965 -164.395 ;
        RECT 312.635 -166.085 312.965 -165.755 ;
        RECT 312.635 -167.445 312.965 -167.115 ;
        RECT 312.635 -168.805 312.965 -168.475 ;
        RECT 312.635 -170.165 312.965 -169.835 ;
        RECT 312.635 -171.525 312.965 -171.195 ;
        RECT 312.635 -172.885 312.965 -172.555 ;
        RECT 312.635 -174.245 312.965 -173.915 ;
        RECT 312.635 -175.605 312.965 -175.275 ;
        RECT 312.635 -176.965 312.965 -176.635 ;
        RECT 312.635 -178.325 312.965 -177.995 ;
        RECT 312.635 -180.57 312.965 -179.44 ;
        RECT 312.64 -180.685 312.96 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 313.995 241.32 314.325 242.45 ;
        RECT 313.995 239.195 314.325 239.525 ;
        RECT 313.995 237.835 314.325 238.165 ;
        RECT 314 237.16 314.32 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 313.995 -95.365 314.325 -95.035 ;
        RECT 313.995 -96.725 314.325 -96.395 ;
        RECT 313.995 -98.085 314.325 -97.755 ;
        RECT 313.995 -99.445 314.325 -99.115 ;
        RECT 313.995 -100.805 314.325 -100.475 ;
        RECT 313.995 -102.165 314.325 -101.835 ;
        RECT 313.995 -103.525 314.325 -103.195 ;
        RECT 313.995 -104.885 314.325 -104.555 ;
        RECT 313.995 -106.245 314.325 -105.915 ;
        RECT 313.995 -107.605 314.325 -107.275 ;
        RECT 313.995 -108.965 314.325 -108.635 ;
        RECT 313.995 -110.325 314.325 -109.995 ;
        RECT 313.995 -111.685 314.325 -111.355 ;
        RECT 313.995 -113.045 314.325 -112.715 ;
        RECT 313.995 -114.405 314.325 -114.075 ;
        RECT 313.995 -115.765 314.325 -115.435 ;
        RECT 313.995 -117.125 314.325 -116.795 ;
        RECT 313.995 -118.485 314.325 -118.155 ;
        RECT 313.995 -119.845 314.325 -119.515 ;
        RECT 313.995 -121.205 314.325 -120.875 ;
        RECT 313.995 -122.565 314.325 -122.235 ;
        RECT 313.995 -123.925 314.325 -123.595 ;
        RECT 313.995 -125.285 314.325 -124.955 ;
        RECT 313.995 -126.645 314.325 -126.315 ;
        RECT 313.995 -128.005 314.325 -127.675 ;
        RECT 313.995 -129.365 314.325 -129.035 ;
        RECT 313.995 -130.725 314.325 -130.395 ;
        RECT 313.995 -132.085 314.325 -131.755 ;
        RECT 313.995 -133.445 314.325 -133.115 ;
        RECT 313.995 -134.805 314.325 -134.475 ;
        RECT 313.995 -136.165 314.325 -135.835 ;
        RECT 313.995 -137.525 314.325 -137.195 ;
        RECT 313.995 -138.885 314.325 -138.555 ;
        RECT 313.995 -140.245 314.325 -139.915 ;
        RECT 313.995 -141.605 314.325 -141.275 ;
        RECT 313.995 -142.965 314.325 -142.635 ;
        RECT 313.995 -144.325 314.325 -143.995 ;
        RECT 313.995 -145.685 314.325 -145.355 ;
        RECT 313.995 -147.045 314.325 -146.715 ;
        RECT 313.995 -148.405 314.325 -148.075 ;
        RECT 313.995 -149.765 314.325 -149.435 ;
        RECT 313.995 -151.125 314.325 -150.795 ;
        RECT 313.995 -152.485 314.325 -152.155 ;
        RECT 313.995 -153.845 314.325 -153.515 ;
        RECT 313.995 -155.205 314.325 -154.875 ;
        RECT 313.995 -156.565 314.325 -156.235 ;
        RECT 313.995 -157.925 314.325 -157.595 ;
        RECT 313.995 -159.285 314.325 -158.955 ;
        RECT 313.995 -160.645 314.325 -160.315 ;
        RECT 313.995 -162.005 314.325 -161.675 ;
        RECT 313.995 -163.365 314.325 -163.035 ;
        RECT 313.995 -164.725 314.325 -164.395 ;
        RECT 313.995 -166.085 314.325 -165.755 ;
        RECT 313.995 -167.445 314.325 -167.115 ;
        RECT 313.995 -168.805 314.325 -168.475 ;
        RECT 313.995 -170.165 314.325 -169.835 ;
        RECT 313.995 -171.525 314.325 -171.195 ;
        RECT 313.995 -172.885 314.325 -172.555 ;
        RECT 313.995 -174.245 314.325 -173.915 ;
        RECT 313.995 -175.605 314.325 -175.275 ;
        RECT 313.995 -176.965 314.325 -176.635 ;
        RECT 313.995 -178.325 314.325 -177.995 ;
        RECT 313.995 -180.57 314.325 -179.44 ;
        RECT 314 -180.685 314.32 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 314.41 -94.075 314.74 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 315.355 241.32 315.685 242.45 ;
        RECT 315.355 239.195 315.685 239.525 ;
        RECT 315.355 237.835 315.685 238.165 ;
        RECT 315.36 237.16 315.68 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 315.355 -1.525 315.685 -1.195 ;
        RECT 315.355 -2.885 315.685 -2.555 ;
        RECT 315.36 -3.56 315.68 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 316.715 241.32 317.045 242.45 ;
        RECT 316.715 239.195 317.045 239.525 ;
        RECT 316.715 237.835 317.045 238.165 ;
        RECT 316.72 237.16 317.04 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 316.715 -1.525 317.045 -1.195 ;
        RECT 316.715 -2.885 317.045 -2.555 ;
        RECT 316.72 -3.56 317.04 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 318.075 241.32 318.405 242.45 ;
        RECT 318.075 239.195 318.405 239.525 ;
        RECT 318.075 237.835 318.405 238.165 ;
        RECT 318.08 237.16 318.4 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 318.075 -1.525 318.405 -1.195 ;
        RECT 318.075 -2.885 318.405 -2.555 ;
        RECT 318.08 -3.56 318.4 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 318.075 -91.285 318.405 -90.955 ;
        RECT 318.075 -92.645 318.405 -92.315 ;
        RECT 318.075 -94.005 318.405 -93.675 ;
        RECT 318.075 -95.365 318.405 -95.035 ;
        RECT 318.075 -96.725 318.405 -96.395 ;
        RECT 318.075 -98.085 318.405 -97.755 ;
        RECT 318.075 -99.445 318.405 -99.115 ;
        RECT 318.075 -100.805 318.405 -100.475 ;
        RECT 318.075 -102.165 318.405 -101.835 ;
        RECT 318.075 -103.525 318.405 -103.195 ;
        RECT 318.075 -104.885 318.405 -104.555 ;
        RECT 318.075 -106.245 318.405 -105.915 ;
        RECT 318.075 -107.605 318.405 -107.275 ;
        RECT 318.075 -108.965 318.405 -108.635 ;
        RECT 318.075 -110.325 318.405 -109.995 ;
        RECT 318.075 -111.685 318.405 -111.355 ;
        RECT 318.075 -113.045 318.405 -112.715 ;
        RECT 318.075 -114.405 318.405 -114.075 ;
        RECT 318.075 -115.765 318.405 -115.435 ;
        RECT 318.075 -117.125 318.405 -116.795 ;
        RECT 318.075 -118.485 318.405 -118.155 ;
        RECT 318.075 -119.845 318.405 -119.515 ;
        RECT 318.075 -121.205 318.405 -120.875 ;
        RECT 318.075 -122.565 318.405 -122.235 ;
        RECT 318.075 -123.925 318.405 -123.595 ;
        RECT 318.075 -125.285 318.405 -124.955 ;
        RECT 318.075 -126.645 318.405 -126.315 ;
        RECT 318.075 -128.005 318.405 -127.675 ;
        RECT 318.075 -129.365 318.405 -129.035 ;
        RECT 318.075 -130.725 318.405 -130.395 ;
        RECT 318.075 -132.085 318.405 -131.755 ;
        RECT 318.075 -133.445 318.405 -133.115 ;
        RECT 318.075 -134.805 318.405 -134.475 ;
        RECT 318.075 -136.165 318.405 -135.835 ;
        RECT 318.075 -137.525 318.405 -137.195 ;
        RECT 318.075 -138.885 318.405 -138.555 ;
        RECT 318.075 -140.245 318.405 -139.915 ;
        RECT 318.075 -141.605 318.405 -141.275 ;
        RECT 318.075 -142.965 318.405 -142.635 ;
        RECT 318.075 -144.325 318.405 -143.995 ;
        RECT 318.075 -145.685 318.405 -145.355 ;
        RECT 318.075 -147.045 318.405 -146.715 ;
        RECT 318.075 -148.405 318.405 -148.075 ;
        RECT 318.075 -149.765 318.405 -149.435 ;
        RECT 318.075 -151.125 318.405 -150.795 ;
        RECT 318.075 -152.485 318.405 -152.155 ;
        RECT 318.075 -153.845 318.405 -153.515 ;
        RECT 318.075 -155.205 318.405 -154.875 ;
        RECT 318.075 -156.565 318.405 -156.235 ;
        RECT 318.075 -157.925 318.405 -157.595 ;
        RECT 318.075 -159.285 318.405 -158.955 ;
        RECT 318.075 -160.645 318.405 -160.315 ;
        RECT 318.075 -162.005 318.405 -161.675 ;
        RECT 318.075 -163.365 318.405 -163.035 ;
        RECT 318.075 -164.725 318.405 -164.395 ;
        RECT 318.075 -166.085 318.405 -165.755 ;
        RECT 318.075 -167.445 318.405 -167.115 ;
        RECT 318.075 -168.805 318.405 -168.475 ;
        RECT 318.075 -170.165 318.405 -169.835 ;
        RECT 318.075 -171.525 318.405 -171.195 ;
        RECT 318.075 -172.885 318.405 -172.555 ;
        RECT 318.075 -174.245 318.405 -173.915 ;
        RECT 318.075 -175.605 318.405 -175.275 ;
        RECT 318.075 -176.965 318.405 -176.635 ;
        RECT 318.075 -178.325 318.405 -177.995 ;
        RECT 318.075 -180.57 318.405 -179.44 ;
        RECT 318.08 -180.685 318.4 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 319.435 241.32 319.765 242.45 ;
        RECT 319.435 239.195 319.765 239.525 ;
        RECT 319.435 237.835 319.765 238.165 ;
        RECT 319.44 237.16 319.76 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 319.435 -95.365 319.765 -95.035 ;
        RECT 319.435 -96.725 319.765 -96.395 ;
        RECT 319.435 -98.085 319.765 -97.755 ;
        RECT 319.435 -99.445 319.765 -99.115 ;
        RECT 319.435 -100.805 319.765 -100.475 ;
        RECT 319.435 -102.165 319.765 -101.835 ;
        RECT 319.435 -103.525 319.765 -103.195 ;
        RECT 319.435 -104.885 319.765 -104.555 ;
        RECT 319.435 -106.245 319.765 -105.915 ;
        RECT 319.435 -107.605 319.765 -107.275 ;
        RECT 319.435 -108.965 319.765 -108.635 ;
        RECT 319.435 -110.325 319.765 -109.995 ;
        RECT 319.435 -111.685 319.765 -111.355 ;
        RECT 319.435 -113.045 319.765 -112.715 ;
        RECT 319.435 -114.405 319.765 -114.075 ;
        RECT 319.435 -115.765 319.765 -115.435 ;
        RECT 319.435 -117.125 319.765 -116.795 ;
        RECT 319.435 -118.485 319.765 -118.155 ;
        RECT 319.435 -119.845 319.765 -119.515 ;
        RECT 319.435 -121.205 319.765 -120.875 ;
        RECT 319.435 -122.565 319.765 -122.235 ;
        RECT 319.435 -123.925 319.765 -123.595 ;
        RECT 319.435 -125.285 319.765 -124.955 ;
        RECT 319.435 -126.645 319.765 -126.315 ;
        RECT 319.435 -128.005 319.765 -127.675 ;
        RECT 319.435 -129.365 319.765 -129.035 ;
        RECT 319.435 -130.725 319.765 -130.395 ;
        RECT 319.435 -132.085 319.765 -131.755 ;
        RECT 319.435 -133.445 319.765 -133.115 ;
        RECT 319.435 -134.805 319.765 -134.475 ;
        RECT 319.435 -136.165 319.765 -135.835 ;
        RECT 319.435 -137.525 319.765 -137.195 ;
        RECT 319.435 -138.885 319.765 -138.555 ;
        RECT 319.435 -140.245 319.765 -139.915 ;
        RECT 319.435 -141.605 319.765 -141.275 ;
        RECT 319.435 -142.965 319.765 -142.635 ;
        RECT 319.435 -144.325 319.765 -143.995 ;
        RECT 319.435 -145.685 319.765 -145.355 ;
        RECT 319.435 -147.045 319.765 -146.715 ;
        RECT 319.435 -148.405 319.765 -148.075 ;
        RECT 319.435 -149.765 319.765 -149.435 ;
        RECT 319.435 -151.125 319.765 -150.795 ;
        RECT 319.435 -152.485 319.765 -152.155 ;
        RECT 319.435 -153.845 319.765 -153.515 ;
        RECT 319.435 -155.205 319.765 -154.875 ;
        RECT 319.435 -156.565 319.765 -156.235 ;
        RECT 319.435 -157.925 319.765 -157.595 ;
        RECT 319.435 -159.285 319.765 -158.955 ;
        RECT 319.435 -160.645 319.765 -160.315 ;
        RECT 319.435 -162.005 319.765 -161.675 ;
        RECT 319.435 -163.365 319.765 -163.035 ;
        RECT 319.435 -164.725 319.765 -164.395 ;
        RECT 319.435 -166.085 319.765 -165.755 ;
        RECT 319.435 -167.445 319.765 -167.115 ;
        RECT 319.435 -168.805 319.765 -168.475 ;
        RECT 319.435 -170.165 319.765 -169.835 ;
        RECT 319.435 -171.525 319.765 -171.195 ;
        RECT 319.435 -172.885 319.765 -172.555 ;
        RECT 319.435 -174.245 319.765 -173.915 ;
        RECT 319.435 -175.605 319.765 -175.275 ;
        RECT 319.435 -176.965 319.765 -176.635 ;
        RECT 319.435 -178.325 319.765 -177.995 ;
        RECT 319.435 -180.57 319.765 -179.44 ;
        RECT 319.44 -180.685 319.76 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 320.51 -94.075 320.84 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 320.795 241.32 321.125 242.45 ;
        RECT 320.795 239.195 321.125 239.525 ;
        RECT 320.795 237.835 321.125 238.165 ;
        RECT 320.8 237.16 321.12 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 322.155 241.32 322.485 242.45 ;
        RECT 322.155 239.195 322.485 239.525 ;
        RECT 322.155 237.835 322.485 238.165 ;
        RECT 322.16 237.16 322.48 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 322.155 -1.525 322.485 -1.195 ;
        RECT 322.155 -2.885 322.485 -2.555 ;
        RECT 322.16 -3.56 322.48 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 323.515 241.32 323.845 242.45 ;
        RECT 323.515 239.195 323.845 239.525 ;
        RECT 323.515 237.835 323.845 238.165 ;
        RECT 323.52 237.16 323.84 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 323.515 -1.525 323.845 -1.195 ;
        RECT 323.515 -2.885 323.845 -2.555 ;
        RECT 323.52 -3.56 323.84 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 324.875 241.32 325.205 242.45 ;
        RECT 324.875 239.195 325.205 239.525 ;
        RECT 324.875 237.835 325.205 238.165 ;
        RECT 324.88 237.16 325.2 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 324.875 -1.525 325.205 -1.195 ;
        RECT 324.875 -2.885 325.205 -2.555 ;
        RECT 324.88 -3.56 325.2 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 324.875 -91.285 325.205 -90.955 ;
        RECT 324.875 -92.645 325.205 -92.315 ;
        RECT 324.875 -94.005 325.205 -93.675 ;
        RECT 324.875 -95.365 325.205 -95.035 ;
        RECT 324.875 -96.725 325.205 -96.395 ;
        RECT 324.875 -98.085 325.205 -97.755 ;
        RECT 324.875 -99.445 325.205 -99.115 ;
        RECT 324.875 -100.805 325.205 -100.475 ;
        RECT 324.875 -102.165 325.205 -101.835 ;
        RECT 324.875 -103.525 325.205 -103.195 ;
        RECT 324.875 -104.885 325.205 -104.555 ;
        RECT 324.875 -106.245 325.205 -105.915 ;
        RECT 324.875 -107.605 325.205 -107.275 ;
        RECT 324.875 -108.965 325.205 -108.635 ;
        RECT 324.875 -110.325 325.205 -109.995 ;
        RECT 324.875 -111.685 325.205 -111.355 ;
        RECT 324.875 -113.045 325.205 -112.715 ;
        RECT 324.875 -114.405 325.205 -114.075 ;
        RECT 324.875 -115.765 325.205 -115.435 ;
        RECT 324.875 -117.125 325.205 -116.795 ;
        RECT 324.875 -118.485 325.205 -118.155 ;
        RECT 324.875 -119.845 325.205 -119.515 ;
        RECT 324.875 -121.205 325.205 -120.875 ;
        RECT 324.875 -122.565 325.205 -122.235 ;
        RECT 324.875 -123.925 325.205 -123.595 ;
        RECT 324.875 -125.285 325.205 -124.955 ;
        RECT 324.875 -126.645 325.205 -126.315 ;
        RECT 324.875 -128.005 325.205 -127.675 ;
        RECT 324.875 -129.365 325.205 -129.035 ;
        RECT 324.875 -130.725 325.205 -130.395 ;
        RECT 324.875 -132.085 325.205 -131.755 ;
        RECT 324.875 -133.445 325.205 -133.115 ;
        RECT 324.875 -134.805 325.205 -134.475 ;
        RECT 324.875 -136.165 325.205 -135.835 ;
        RECT 324.875 -137.525 325.205 -137.195 ;
        RECT 324.875 -138.885 325.205 -138.555 ;
        RECT 324.875 -140.245 325.205 -139.915 ;
        RECT 324.875 -141.605 325.205 -141.275 ;
        RECT 324.875 -142.965 325.205 -142.635 ;
        RECT 324.875 -144.325 325.205 -143.995 ;
        RECT 324.875 -145.685 325.205 -145.355 ;
        RECT 324.875 -147.045 325.205 -146.715 ;
        RECT 324.875 -148.405 325.205 -148.075 ;
        RECT 324.875 -149.765 325.205 -149.435 ;
        RECT 324.875 -151.125 325.205 -150.795 ;
        RECT 324.875 -152.485 325.205 -152.155 ;
        RECT 324.875 -153.845 325.205 -153.515 ;
        RECT 324.875 -155.205 325.205 -154.875 ;
        RECT 324.875 -156.565 325.205 -156.235 ;
        RECT 324.875 -157.925 325.205 -157.595 ;
        RECT 324.875 -159.285 325.205 -158.955 ;
        RECT 324.875 -160.645 325.205 -160.315 ;
        RECT 324.875 -162.005 325.205 -161.675 ;
        RECT 324.875 -163.365 325.205 -163.035 ;
        RECT 324.875 -164.725 325.205 -164.395 ;
        RECT 324.875 -166.085 325.205 -165.755 ;
        RECT 324.875 -167.445 325.205 -167.115 ;
        RECT 324.875 -168.805 325.205 -168.475 ;
        RECT 324.875 -170.165 325.205 -169.835 ;
        RECT 324.875 -171.525 325.205 -171.195 ;
        RECT 324.875 -172.885 325.205 -172.555 ;
        RECT 324.875 -174.245 325.205 -173.915 ;
        RECT 324.875 -175.605 325.205 -175.275 ;
        RECT 324.875 -176.965 325.205 -176.635 ;
        RECT 324.875 -178.325 325.205 -177.995 ;
        RECT 324.875 -180.57 325.205 -179.44 ;
        RECT 324.88 -180.685 325.2 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 326.235 241.32 326.565 242.45 ;
        RECT 326.235 239.195 326.565 239.525 ;
        RECT 326.235 237.835 326.565 238.165 ;
        RECT 326.24 237.16 326.56 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 326.235 -95.365 326.565 -95.035 ;
        RECT 326.235 -96.725 326.565 -96.395 ;
        RECT 326.235 -98.085 326.565 -97.755 ;
        RECT 326.235 -99.445 326.565 -99.115 ;
        RECT 326.235 -100.805 326.565 -100.475 ;
        RECT 326.235 -102.165 326.565 -101.835 ;
        RECT 326.235 -103.525 326.565 -103.195 ;
        RECT 326.235 -104.885 326.565 -104.555 ;
        RECT 326.235 -106.245 326.565 -105.915 ;
        RECT 326.235 -107.605 326.565 -107.275 ;
        RECT 326.235 -108.965 326.565 -108.635 ;
        RECT 326.235 -110.325 326.565 -109.995 ;
        RECT 326.235 -111.685 326.565 -111.355 ;
        RECT 326.235 -113.045 326.565 -112.715 ;
        RECT 326.235 -114.405 326.565 -114.075 ;
        RECT 326.235 -115.765 326.565 -115.435 ;
        RECT 326.235 -117.125 326.565 -116.795 ;
        RECT 326.235 -118.485 326.565 -118.155 ;
        RECT 326.235 -119.845 326.565 -119.515 ;
        RECT 326.235 -121.205 326.565 -120.875 ;
        RECT 326.235 -122.565 326.565 -122.235 ;
        RECT 326.235 -123.925 326.565 -123.595 ;
        RECT 326.235 -125.285 326.565 -124.955 ;
        RECT 326.235 -126.645 326.565 -126.315 ;
        RECT 326.235 -128.005 326.565 -127.675 ;
        RECT 326.235 -129.365 326.565 -129.035 ;
        RECT 326.235 -130.725 326.565 -130.395 ;
        RECT 326.235 -132.085 326.565 -131.755 ;
        RECT 326.235 -133.445 326.565 -133.115 ;
        RECT 326.235 -134.805 326.565 -134.475 ;
        RECT 326.235 -136.165 326.565 -135.835 ;
        RECT 326.235 -137.525 326.565 -137.195 ;
        RECT 326.235 -138.885 326.565 -138.555 ;
        RECT 326.235 -140.245 326.565 -139.915 ;
        RECT 326.235 -141.605 326.565 -141.275 ;
        RECT 326.235 -142.965 326.565 -142.635 ;
        RECT 326.235 -144.325 326.565 -143.995 ;
        RECT 326.235 -145.685 326.565 -145.355 ;
        RECT 326.235 -147.045 326.565 -146.715 ;
        RECT 326.235 -148.405 326.565 -148.075 ;
        RECT 326.235 -149.765 326.565 -149.435 ;
        RECT 326.235 -151.125 326.565 -150.795 ;
        RECT 326.235 -152.485 326.565 -152.155 ;
        RECT 326.235 -153.845 326.565 -153.515 ;
        RECT 326.235 -155.205 326.565 -154.875 ;
        RECT 326.235 -156.565 326.565 -156.235 ;
        RECT 326.235 -157.925 326.565 -157.595 ;
        RECT 326.235 -159.285 326.565 -158.955 ;
        RECT 326.235 -160.645 326.565 -160.315 ;
        RECT 326.235 -162.005 326.565 -161.675 ;
        RECT 326.235 -163.365 326.565 -163.035 ;
        RECT 326.235 -164.725 326.565 -164.395 ;
        RECT 326.235 -166.085 326.565 -165.755 ;
        RECT 326.235 -167.445 326.565 -167.115 ;
        RECT 326.235 -168.805 326.565 -168.475 ;
        RECT 326.235 -170.165 326.565 -169.835 ;
        RECT 326.235 -171.525 326.565 -171.195 ;
        RECT 326.235 -172.885 326.565 -172.555 ;
        RECT 326.235 -174.245 326.565 -173.915 ;
        RECT 326.235 -175.605 326.565 -175.275 ;
        RECT 326.235 -176.965 326.565 -176.635 ;
        RECT 326.235 -178.325 326.565 -177.995 ;
        RECT 326.235 -180.57 326.565 -179.44 ;
        RECT 326.24 -180.685 326.56 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 326.61 -94.075 326.94 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 327.595 241.32 327.925 242.45 ;
        RECT 327.595 239.195 327.925 239.525 ;
        RECT 327.595 237.835 327.925 238.165 ;
        RECT 327.6 237.16 327.92 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 327.595 -1.525 327.925 -1.195 ;
        RECT 327.595 -2.885 327.925 -2.555 ;
        RECT 327.6 -3.56 327.92 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 328.955 241.32 329.285 242.45 ;
        RECT 328.955 239.195 329.285 239.525 ;
        RECT 328.955 237.835 329.285 238.165 ;
        RECT 328.96 237.16 329.28 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 328.955 -1.525 329.285 -1.195 ;
        RECT 328.955 -2.885 329.285 -2.555 ;
        RECT 328.96 -3.56 329.28 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 330.315 241.32 330.645 242.45 ;
        RECT 330.315 239.195 330.645 239.525 ;
        RECT 330.315 237.835 330.645 238.165 ;
        RECT 330.32 237.16 330.64 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 330.315 -1.525 330.645 -1.195 ;
        RECT 330.315 -2.885 330.645 -2.555 ;
        RECT 330.32 -3.56 330.64 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 330.315 -91.285 330.645 -90.955 ;
        RECT 330.315 -92.645 330.645 -92.315 ;
        RECT 330.315 -94.005 330.645 -93.675 ;
        RECT 330.315 -95.365 330.645 -95.035 ;
        RECT 330.315 -96.725 330.645 -96.395 ;
        RECT 330.315 -98.085 330.645 -97.755 ;
        RECT 330.315 -99.445 330.645 -99.115 ;
        RECT 330.315 -100.805 330.645 -100.475 ;
        RECT 330.315 -102.165 330.645 -101.835 ;
        RECT 330.315 -103.525 330.645 -103.195 ;
        RECT 330.315 -104.885 330.645 -104.555 ;
        RECT 330.315 -106.245 330.645 -105.915 ;
        RECT 330.315 -107.605 330.645 -107.275 ;
        RECT 330.315 -108.965 330.645 -108.635 ;
        RECT 330.315 -110.325 330.645 -109.995 ;
        RECT 330.315 -111.685 330.645 -111.355 ;
        RECT 330.315 -113.045 330.645 -112.715 ;
        RECT 330.315 -114.405 330.645 -114.075 ;
        RECT 330.315 -115.765 330.645 -115.435 ;
        RECT 330.315 -117.125 330.645 -116.795 ;
        RECT 330.315 -118.485 330.645 -118.155 ;
        RECT 330.315 -119.845 330.645 -119.515 ;
        RECT 330.315 -121.205 330.645 -120.875 ;
        RECT 330.315 -122.565 330.645 -122.235 ;
        RECT 330.315 -123.925 330.645 -123.595 ;
        RECT 330.315 -125.285 330.645 -124.955 ;
        RECT 330.315 -126.645 330.645 -126.315 ;
        RECT 330.315 -128.005 330.645 -127.675 ;
        RECT 330.315 -129.365 330.645 -129.035 ;
        RECT 330.315 -130.725 330.645 -130.395 ;
        RECT 330.315 -132.085 330.645 -131.755 ;
        RECT 330.315 -133.445 330.645 -133.115 ;
        RECT 330.315 -134.805 330.645 -134.475 ;
        RECT 330.315 -136.165 330.645 -135.835 ;
        RECT 330.315 -137.525 330.645 -137.195 ;
        RECT 330.315 -138.885 330.645 -138.555 ;
        RECT 330.315 -140.245 330.645 -139.915 ;
        RECT 330.315 -141.605 330.645 -141.275 ;
        RECT 330.315 -142.965 330.645 -142.635 ;
        RECT 330.315 -144.325 330.645 -143.995 ;
        RECT 330.315 -145.685 330.645 -145.355 ;
        RECT 330.315 -147.045 330.645 -146.715 ;
        RECT 330.315 -148.405 330.645 -148.075 ;
        RECT 330.315 -149.765 330.645 -149.435 ;
        RECT 330.315 -151.125 330.645 -150.795 ;
        RECT 330.315 -152.485 330.645 -152.155 ;
        RECT 330.315 -153.845 330.645 -153.515 ;
        RECT 330.315 -155.205 330.645 -154.875 ;
        RECT 330.315 -156.565 330.645 -156.235 ;
        RECT 330.315 -157.925 330.645 -157.595 ;
        RECT 330.315 -159.285 330.645 -158.955 ;
        RECT 330.315 -160.645 330.645 -160.315 ;
        RECT 330.315 -162.005 330.645 -161.675 ;
        RECT 330.315 -163.365 330.645 -163.035 ;
        RECT 330.315 -164.725 330.645 -164.395 ;
        RECT 330.315 -166.085 330.645 -165.755 ;
        RECT 330.315 -167.445 330.645 -167.115 ;
        RECT 330.315 -168.805 330.645 -168.475 ;
        RECT 330.315 -170.165 330.645 -169.835 ;
        RECT 330.315 -171.525 330.645 -171.195 ;
        RECT 330.315 -172.885 330.645 -172.555 ;
        RECT 330.315 -174.245 330.645 -173.915 ;
        RECT 330.315 -175.605 330.645 -175.275 ;
        RECT 330.315 -176.965 330.645 -176.635 ;
        RECT 330.315 -178.325 330.645 -177.995 ;
        RECT 330.315 -180.57 330.645 -179.44 ;
        RECT 330.32 -180.685 330.64 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 331.675 241.32 332.005 242.45 ;
        RECT 331.675 239.195 332.005 239.525 ;
        RECT 331.675 237.835 332.005 238.165 ;
        RECT 331.68 237.16 332 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 331.675 -95.365 332.005 -95.035 ;
        RECT 331.675 -96.725 332.005 -96.395 ;
        RECT 331.675 -98.085 332.005 -97.755 ;
        RECT 331.675 -99.445 332.005 -99.115 ;
        RECT 331.675 -100.805 332.005 -100.475 ;
        RECT 331.675 -102.165 332.005 -101.835 ;
        RECT 331.675 -103.525 332.005 -103.195 ;
        RECT 331.675 -104.885 332.005 -104.555 ;
        RECT 331.675 -106.245 332.005 -105.915 ;
        RECT 331.675 -107.605 332.005 -107.275 ;
        RECT 331.675 -108.965 332.005 -108.635 ;
        RECT 331.675 -110.325 332.005 -109.995 ;
        RECT 331.675 -111.685 332.005 -111.355 ;
        RECT 331.675 -113.045 332.005 -112.715 ;
        RECT 331.675 -114.405 332.005 -114.075 ;
        RECT 331.675 -115.765 332.005 -115.435 ;
        RECT 331.675 -117.125 332.005 -116.795 ;
        RECT 331.675 -118.485 332.005 -118.155 ;
        RECT 331.675 -119.845 332.005 -119.515 ;
        RECT 331.675 -121.205 332.005 -120.875 ;
        RECT 331.675 -122.565 332.005 -122.235 ;
        RECT 331.675 -123.925 332.005 -123.595 ;
        RECT 331.675 -125.285 332.005 -124.955 ;
        RECT 331.675 -126.645 332.005 -126.315 ;
        RECT 331.675 -128.005 332.005 -127.675 ;
        RECT 331.675 -129.365 332.005 -129.035 ;
        RECT 331.675 -130.725 332.005 -130.395 ;
        RECT 331.675 -132.085 332.005 -131.755 ;
        RECT 331.675 -133.445 332.005 -133.115 ;
        RECT 331.675 -134.805 332.005 -134.475 ;
        RECT 331.675 -136.165 332.005 -135.835 ;
        RECT 331.675 -137.525 332.005 -137.195 ;
        RECT 331.675 -138.885 332.005 -138.555 ;
        RECT 331.675 -140.245 332.005 -139.915 ;
        RECT 331.675 -141.605 332.005 -141.275 ;
        RECT 331.675 -142.965 332.005 -142.635 ;
        RECT 331.675 -144.325 332.005 -143.995 ;
        RECT 331.675 -145.685 332.005 -145.355 ;
        RECT 331.675 -147.045 332.005 -146.715 ;
        RECT 331.675 -148.405 332.005 -148.075 ;
        RECT 331.675 -149.765 332.005 -149.435 ;
        RECT 331.675 -151.125 332.005 -150.795 ;
        RECT 331.675 -152.485 332.005 -152.155 ;
        RECT 331.675 -153.845 332.005 -153.515 ;
        RECT 331.675 -155.205 332.005 -154.875 ;
        RECT 331.675 -156.565 332.005 -156.235 ;
        RECT 331.675 -157.925 332.005 -157.595 ;
        RECT 331.675 -159.285 332.005 -158.955 ;
        RECT 331.675 -160.645 332.005 -160.315 ;
        RECT 331.675 -162.005 332.005 -161.675 ;
        RECT 331.675 -163.365 332.005 -163.035 ;
        RECT 331.675 -164.725 332.005 -164.395 ;
        RECT 331.675 -166.085 332.005 -165.755 ;
        RECT 331.675 -167.445 332.005 -167.115 ;
        RECT 331.675 -168.805 332.005 -168.475 ;
        RECT 331.675 -170.165 332.005 -169.835 ;
        RECT 331.675 -171.525 332.005 -171.195 ;
        RECT 331.675 -172.885 332.005 -172.555 ;
        RECT 331.675 -174.245 332.005 -173.915 ;
        RECT 331.675 -175.605 332.005 -175.275 ;
        RECT 331.675 -176.965 332.005 -176.635 ;
        RECT 331.675 -178.325 332.005 -177.995 ;
        RECT 331.675 -180.57 332.005 -179.44 ;
        RECT 331.68 -180.685 332 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 332.71 -94.075 333.04 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 333.035 241.32 333.365 242.45 ;
        RECT 333.035 239.195 333.365 239.525 ;
        RECT 333.035 237.835 333.365 238.165 ;
        RECT 333.04 237.16 333.36 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 334.395 241.32 334.725 242.45 ;
        RECT 334.395 239.195 334.725 239.525 ;
        RECT 334.395 237.835 334.725 238.165 ;
        RECT 334.4 237.16 334.72 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 334.395 -1.525 334.725 -1.195 ;
        RECT 334.395 -2.885 334.725 -2.555 ;
        RECT 334.4 -3.56 334.72 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 335.755 241.32 336.085 242.45 ;
        RECT 335.755 239.195 336.085 239.525 ;
        RECT 335.755 237.835 336.085 238.165 ;
        RECT 335.76 237.16 336.08 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 335.755 -1.525 336.085 -1.195 ;
        RECT 335.755 -2.885 336.085 -2.555 ;
        RECT 335.76 -3.56 336.08 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 335.755 -118.485 336.085 -118.155 ;
        RECT 335.755 -119.845 336.085 -119.515 ;
        RECT 335.755 -121.205 336.085 -120.875 ;
        RECT 335.755 -122.565 336.085 -122.235 ;
        RECT 335.755 -123.925 336.085 -123.595 ;
        RECT 335.755 -125.285 336.085 -124.955 ;
        RECT 335.755 -126.645 336.085 -126.315 ;
        RECT 335.755 -128.005 336.085 -127.675 ;
        RECT 335.755 -129.365 336.085 -129.035 ;
        RECT 335.755 -130.725 336.085 -130.395 ;
        RECT 335.755 -132.085 336.085 -131.755 ;
        RECT 335.755 -133.445 336.085 -133.115 ;
        RECT 335.755 -134.805 336.085 -134.475 ;
        RECT 335.755 -136.165 336.085 -135.835 ;
        RECT 335.755 -137.525 336.085 -137.195 ;
        RECT 335.755 -138.885 336.085 -138.555 ;
        RECT 335.755 -140.245 336.085 -139.915 ;
        RECT 335.755 -141.605 336.085 -141.275 ;
        RECT 335.755 -142.965 336.085 -142.635 ;
        RECT 335.755 -144.325 336.085 -143.995 ;
        RECT 335.755 -145.685 336.085 -145.355 ;
        RECT 335.755 -147.045 336.085 -146.715 ;
        RECT 335.755 -148.405 336.085 -148.075 ;
        RECT 335.755 -149.765 336.085 -149.435 ;
        RECT 335.755 -151.125 336.085 -150.795 ;
        RECT 335.755 -152.485 336.085 -152.155 ;
        RECT 335.755 -153.845 336.085 -153.515 ;
        RECT 335.755 -155.205 336.085 -154.875 ;
        RECT 335.755 -156.565 336.085 -156.235 ;
        RECT 335.755 -157.925 336.085 -157.595 ;
        RECT 335.755 -159.285 336.085 -158.955 ;
        RECT 335.755 -160.645 336.085 -160.315 ;
        RECT 335.755 -162.005 336.085 -161.675 ;
        RECT 335.755 -163.365 336.085 -163.035 ;
        RECT 335.755 -164.725 336.085 -164.395 ;
        RECT 335.755 -166.085 336.085 -165.755 ;
        RECT 335.755 -167.445 336.085 -167.115 ;
        RECT 335.755 -168.805 336.085 -168.475 ;
        RECT 335.755 -170.165 336.085 -169.835 ;
        RECT 335.755 -171.525 336.085 -171.195 ;
        RECT 335.755 -172.885 336.085 -172.555 ;
        RECT 335.755 -174.245 336.085 -173.915 ;
        RECT 335.755 -175.605 336.085 -175.275 ;
        RECT 335.755 -176.965 336.085 -176.635 ;
        RECT 335.755 -178.325 336.085 -177.995 ;
        RECT 335.755 -180.57 336.085 -179.44 ;
        RECT 335.76 -180.685 336.08 -90.955 ;
        RECT 335.755 -91.285 336.085 -90.955 ;
        RECT 335.755 -92.645 336.085 -92.315 ;
        RECT 335.755 -94.005 336.085 -93.675 ;
        RECT 335.755 -95.365 336.085 -95.035 ;
        RECT 335.755 -96.725 336.085 -96.395 ;
        RECT 335.755 -98.085 336.085 -97.755 ;
        RECT 335.755 -99.445 336.085 -99.115 ;
        RECT 335.755 -100.805 336.085 -100.475 ;
        RECT 335.755 -102.165 336.085 -101.835 ;
        RECT 335.755 -103.525 336.085 -103.195 ;
        RECT 335.755 -104.885 336.085 -104.555 ;
        RECT 335.755 -106.245 336.085 -105.915 ;
        RECT 335.755 -107.605 336.085 -107.275 ;
        RECT 335.755 -108.965 336.085 -108.635 ;
        RECT 335.755 -110.325 336.085 -109.995 ;
        RECT 335.755 -111.685 336.085 -111.355 ;
        RECT 335.755 -113.045 336.085 -112.715 ;
        RECT 335.755 -114.405 336.085 -114.075 ;
        RECT 335.755 -115.765 336.085 -115.435 ;
        RECT 335.755 -117.125 336.085 -116.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 270.475 241.32 270.805 242.45 ;
        RECT 270.475 239.195 270.805 239.525 ;
        RECT 270.475 237.835 270.805 238.165 ;
        RECT 270.48 237.16 270.8 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 270.475 -95.365 270.805 -95.035 ;
        RECT 270.475 -96.725 270.805 -96.395 ;
        RECT 270.475 -98.085 270.805 -97.755 ;
        RECT 270.475 -99.445 270.805 -99.115 ;
        RECT 270.475 -100.805 270.805 -100.475 ;
        RECT 270.475 -102.165 270.805 -101.835 ;
        RECT 270.475 -103.525 270.805 -103.195 ;
        RECT 270.475 -104.885 270.805 -104.555 ;
        RECT 270.475 -106.245 270.805 -105.915 ;
        RECT 270.475 -107.605 270.805 -107.275 ;
        RECT 270.475 -108.965 270.805 -108.635 ;
        RECT 270.475 -110.325 270.805 -109.995 ;
        RECT 270.475 -111.685 270.805 -111.355 ;
        RECT 270.475 -113.045 270.805 -112.715 ;
        RECT 270.475 -114.405 270.805 -114.075 ;
        RECT 270.475 -115.765 270.805 -115.435 ;
        RECT 270.475 -117.125 270.805 -116.795 ;
        RECT 270.475 -118.485 270.805 -118.155 ;
        RECT 270.475 -119.845 270.805 -119.515 ;
        RECT 270.475 -121.205 270.805 -120.875 ;
        RECT 270.475 -122.565 270.805 -122.235 ;
        RECT 270.475 -123.925 270.805 -123.595 ;
        RECT 270.475 -125.285 270.805 -124.955 ;
        RECT 270.475 -126.645 270.805 -126.315 ;
        RECT 270.475 -128.005 270.805 -127.675 ;
        RECT 270.475 -129.365 270.805 -129.035 ;
        RECT 270.475 -130.725 270.805 -130.395 ;
        RECT 270.475 -132.085 270.805 -131.755 ;
        RECT 270.475 -133.445 270.805 -133.115 ;
        RECT 270.475 -134.805 270.805 -134.475 ;
        RECT 270.475 -136.165 270.805 -135.835 ;
        RECT 270.475 -137.525 270.805 -137.195 ;
        RECT 270.475 -138.885 270.805 -138.555 ;
        RECT 270.475 -140.245 270.805 -139.915 ;
        RECT 270.475 -141.605 270.805 -141.275 ;
        RECT 270.475 -142.965 270.805 -142.635 ;
        RECT 270.475 -144.325 270.805 -143.995 ;
        RECT 270.475 -145.685 270.805 -145.355 ;
        RECT 270.475 -147.045 270.805 -146.715 ;
        RECT 270.475 -148.405 270.805 -148.075 ;
        RECT 270.475 -149.765 270.805 -149.435 ;
        RECT 270.475 -151.125 270.805 -150.795 ;
        RECT 270.475 -152.485 270.805 -152.155 ;
        RECT 270.475 -153.845 270.805 -153.515 ;
        RECT 270.475 -155.205 270.805 -154.875 ;
        RECT 270.475 -156.565 270.805 -156.235 ;
        RECT 270.475 -157.925 270.805 -157.595 ;
        RECT 270.475 -159.285 270.805 -158.955 ;
        RECT 270.475 -160.645 270.805 -160.315 ;
        RECT 270.475 -162.005 270.805 -161.675 ;
        RECT 270.475 -163.365 270.805 -163.035 ;
        RECT 270.475 -164.725 270.805 -164.395 ;
        RECT 270.475 -166.085 270.805 -165.755 ;
        RECT 270.475 -167.445 270.805 -167.115 ;
        RECT 270.475 -168.805 270.805 -168.475 ;
        RECT 270.475 -170.165 270.805 -169.835 ;
        RECT 270.475 -171.525 270.805 -171.195 ;
        RECT 270.475 -172.885 270.805 -172.555 ;
        RECT 270.475 -174.245 270.805 -173.915 ;
        RECT 270.475 -175.605 270.805 -175.275 ;
        RECT 270.475 -176.965 270.805 -176.635 ;
        RECT 270.475 -178.325 270.805 -177.995 ;
        RECT 270.475 -180.57 270.805 -179.44 ;
        RECT 270.48 -180.685 270.8 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 271.71 -94.075 272.04 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 271.835 241.32 272.165 242.45 ;
        RECT 271.835 239.195 272.165 239.525 ;
        RECT 271.835 237.835 272.165 238.165 ;
        RECT 271.84 237.16 272.16 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 273.195 241.32 273.525 242.45 ;
        RECT 273.195 239.195 273.525 239.525 ;
        RECT 273.195 237.835 273.525 238.165 ;
        RECT 273.2 237.16 273.52 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 273.195 -1.525 273.525 -1.195 ;
        RECT 273.195 -2.885 273.525 -2.555 ;
        RECT 273.2 -3.56 273.52 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 273.195 -91.285 273.525 -90.955 ;
        RECT 273.195 -92.645 273.525 -92.315 ;
        RECT 273.195 -94.005 273.525 -93.675 ;
        RECT 273.195 -95.365 273.525 -95.035 ;
        RECT 273.195 -96.725 273.525 -96.395 ;
        RECT 273.195 -98.085 273.525 -97.755 ;
        RECT 273.195 -99.445 273.525 -99.115 ;
        RECT 273.195 -100.805 273.525 -100.475 ;
        RECT 273.195 -102.165 273.525 -101.835 ;
        RECT 273.195 -103.525 273.525 -103.195 ;
        RECT 273.195 -104.885 273.525 -104.555 ;
        RECT 273.195 -106.245 273.525 -105.915 ;
        RECT 273.195 -107.605 273.525 -107.275 ;
        RECT 273.195 -108.965 273.525 -108.635 ;
        RECT 273.195 -110.325 273.525 -109.995 ;
        RECT 273.195 -111.685 273.525 -111.355 ;
        RECT 273.195 -113.045 273.525 -112.715 ;
        RECT 273.195 -114.405 273.525 -114.075 ;
        RECT 273.195 -115.765 273.525 -115.435 ;
        RECT 273.195 -117.125 273.525 -116.795 ;
        RECT 273.195 -118.485 273.525 -118.155 ;
        RECT 273.195 -119.845 273.525 -119.515 ;
        RECT 273.195 -121.205 273.525 -120.875 ;
        RECT 273.195 -122.565 273.525 -122.235 ;
        RECT 273.195 -123.925 273.525 -123.595 ;
        RECT 273.195 -125.285 273.525 -124.955 ;
        RECT 273.195 -126.645 273.525 -126.315 ;
        RECT 273.195 -128.005 273.525 -127.675 ;
        RECT 273.195 -129.365 273.525 -129.035 ;
        RECT 273.195 -130.725 273.525 -130.395 ;
        RECT 273.195 -132.085 273.525 -131.755 ;
        RECT 273.195 -133.445 273.525 -133.115 ;
        RECT 273.195 -134.805 273.525 -134.475 ;
        RECT 273.195 -136.165 273.525 -135.835 ;
        RECT 273.195 -137.525 273.525 -137.195 ;
        RECT 273.195 -138.885 273.525 -138.555 ;
        RECT 273.195 -140.245 273.525 -139.915 ;
        RECT 273.195 -141.605 273.525 -141.275 ;
        RECT 273.195 -142.965 273.525 -142.635 ;
        RECT 273.195 -144.325 273.525 -143.995 ;
        RECT 273.195 -145.685 273.525 -145.355 ;
        RECT 273.195 -147.045 273.525 -146.715 ;
        RECT 273.195 -148.405 273.525 -148.075 ;
        RECT 273.195 -149.765 273.525 -149.435 ;
        RECT 273.195 -151.125 273.525 -150.795 ;
        RECT 273.195 -152.485 273.525 -152.155 ;
        RECT 273.195 -153.845 273.525 -153.515 ;
        RECT 273.195 -155.205 273.525 -154.875 ;
        RECT 273.195 -156.565 273.525 -156.235 ;
        RECT 273.195 -157.925 273.525 -157.595 ;
        RECT 273.195 -159.285 273.525 -158.955 ;
        RECT 273.195 -160.645 273.525 -160.315 ;
        RECT 273.195 -162.005 273.525 -161.675 ;
        RECT 273.195 -163.365 273.525 -163.035 ;
        RECT 273.195 -164.725 273.525 -164.395 ;
        RECT 273.195 -166.085 273.525 -165.755 ;
        RECT 273.195 -167.445 273.525 -167.115 ;
        RECT 273.195 -168.805 273.525 -168.475 ;
        RECT 273.195 -170.165 273.525 -169.835 ;
        RECT 273.195 -171.525 273.525 -171.195 ;
        RECT 273.195 -172.885 273.525 -172.555 ;
        RECT 273.195 -174.245 273.525 -173.915 ;
        RECT 273.195 -175.605 273.525 -175.275 ;
        RECT 273.195 -176.965 273.525 -176.635 ;
        RECT 273.195 -178.325 273.525 -177.995 ;
        RECT 273.195 -180.57 273.525 -179.44 ;
        RECT 273.2 -180.685 273.52 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 274.555 241.32 274.885 242.45 ;
        RECT 274.555 239.195 274.885 239.525 ;
        RECT 274.555 237.835 274.885 238.165 ;
        RECT 274.56 237.16 274.88 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 274.555 -1.525 274.885 -1.195 ;
        RECT 274.555 -2.885 274.885 -2.555 ;
        RECT 274.56 -3.56 274.88 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 275.915 241.32 276.245 242.45 ;
        RECT 275.915 239.195 276.245 239.525 ;
        RECT 275.915 237.835 276.245 238.165 ;
        RECT 275.92 237.16 276.24 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 275.915 -1.525 276.245 -1.195 ;
        RECT 275.915 -2.885 276.245 -2.555 ;
        RECT 275.92 -3.56 276.24 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 275.915 -91.285 276.245 -90.955 ;
        RECT 275.915 -92.645 276.245 -92.315 ;
        RECT 275.915 -94.005 276.245 -93.675 ;
        RECT 275.915 -95.365 276.245 -95.035 ;
        RECT 275.915 -96.725 276.245 -96.395 ;
        RECT 275.915 -98.085 276.245 -97.755 ;
        RECT 275.915 -99.445 276.245 -99.115 ;
        RECT 275.915 -100.805 276.245 -100.475 ;
        RECT 275.915 -102.165 276.245 -101.835 ;
        RECT 275.915 -103.525 276.245 -103.195 ;
        RECT 275.915 -104.885 276.245 -104.555 ;
        RECT 275.915 -106.245 276.245 -105.915 ;
        RECT 275.915 -107.605 276.245 -107.275 ;
        RECT 275.915 -108.965 276.245 -108.635 ;
        RECT 275.915 -110.325 276.245 -109.995 ;
        RECT 275.915 -111.685 276.245 -111.355 ;
        RECT 275.915 -113.045 276.245 -112.715 ;
        RECT 275.915 -114.405 276.245 -114.075 ;
        RECT 275.915 -115.765 276.245 -115.435 ;
        RECT 275.915 -117.125 276.245 -116.795 ;
        RECT 275.915 -118.485 276.245 -118.155 ;
        RECT 275.915 -119.845 276.245 -119.515 ;
        RECT 275.915 -121.205 276.245 -120.875 ;
        RECT 275.915 -122.565 276.245 -122.235 ;
        RECT 275.915 -123.925 276.245 -123.595 ;
        RECT 275.915 -125.285 276.245 -124.955 ;
        RECT 275.915 -126.645 276.245 -126.315 ;
        RECT 275.915 -128.005 276.245 -127.675 ;
        RECT 275.915 -129.365 276.245 -129.035 ;
        RECT 275.915 -130.725 276.245 -130.395 ;
        RECT 275.915 -132.085 276.245 -131.755 ;
        RECT 275.915 -133.445 276.245 -133.115 ;
        RECT 275.915 -134.805 276.245 -134.475 ;
        RECT 275.915 -136.165 276.245 -135.835 ;
        RECT 275.915 -137.525 276.245 -137.195 ;
        RECT 275.915 -138.885 276.245 -138.555 ;
        RECT 275.915 -140.245 276.245 -139.915 ;
        RECT 275.915 -141.605 276.245 -141.275 ;
        RECT 275.915 -142.965 276.245 -142.635 ;
        RECT 275.915 -144.325 276.245 -143.995 ;
        RECT 275.915 -145.685 276.245 -145.355 ;
        RECT 275.915 -147.045 276.245 -146.715 ;
        RECT 275.915 -148.405 276.245 -148.075 ;
        RECT 275.915 -149.765 276.245 -149.435 ;
        RECT 275.915 -151.125 276.245 -150.795 ;
        RECT 275.915 -152.485 276.245 -152.155 ;
        RECT 275.915 -153.845 276.245 -153.515 ;
        RECT 275.915 -155.205 276.245 -154.875 ;
        RECT 275.915 -156.565 276.245 -156.235 ;
        RECT 275.915 -157.925 276.245 -157.595 ;
        RECT 275.915 -159.285 276.245 -158.955 ;
        RECT 275.915 -160.645 276.245 -160.315 ;
        RECT 275.915 -162.005 276.245 -161.675 ;
        RECT 275.915 -163.365 276.245 -163.035 ;
        RECT 275.915 -164.725 276.245 -164.395 ;
        RECT 275.915 -166.085 276.245 -165.755 ;
        RECT 275.915 -167.445 276.245 -167.115 ;
        RECT 275.915 -168.805 276.245 -168.475 ;
        RECT 275.915 -170.165 276.245 -169.835 ;
        RECT 275.915 -171.525 276.245 -171.195 ;
        RECT 275.915 -172.885 276.245 -172.555 ;
        RECT 275.915 -174.245 276.245 -173.915 ;
        RECT 275.915 -175.605 276.245 -175.275 ;
        RECT 275.915 -176.965 276.245 -176.635 ;
        RECT 275.915 -178.325 276.245 -177.995 ;
        RECT 275.915 -180.57 276.245 -179.44 ;
        RECT 275.92 -180.685 276.24 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 277.275 241.32 277.605 242.45 ;
        RECT 277.275 239.195 277.605 239.525 ;
        RECT 277.275 237.835 277.605 238.165 ;
        RECT 277.28 237.16 277.6 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 277.275 -95.365 277.605 -95.035 ;
        RECT 277.275 -96.725 277.605 -96.395 ;
        RECT 277.275 -98.085 277.605 -97.755 ;
        RECT 277.275 -99.445 277.605 -99.115 ;
        RECT 277.275 -100.805 277.605 -100.475 ;
        RECT 277.275 -102.165 277.605 -101.835 ;
        RECT 277.275 -103.525 277.605 -103.195 ;
        RECT 277.275 -104.885 277.605 -104.555 ;
        RECT 277.275 -106.245 277.605 -105.915 ;
        RECT 277.275 -107.605 277.605 -107.275 ;
        RECT 277.275 -108.965 277.605 -108.635 ;
        RECT 277.275 -110.325 277.605 -109.995 ;
        RECT 277.275 -111.685 277.605 -111.355 ;
        RECT 277.275 -113.045 277.605 -112.715 ;
        RECT 277.275 -114.405 277.605 -114.075 ;
        RECT 277.275 -115.765 277.605 -115.435 ;
        RECT 277.275 -117.125 277.605 -116.795 ;
        RECT 277.275 -118.485 277.605 -118.155 ;
        RECT 277.275 -119.845 277.605 -119.515 ;
        RECT 277.275 -121.205 277.605 -120.875 ;
        RECT 277.275 -122.565 277.605 -122.235 ;
        RECT 277.275 -123.925 277.605 -123.595 ;
        RECT 277.275 -125.285 277.605 -124.955 ;
        RECT 277.275 -126.645 277.605 -126.315 ;
        RECT 277.275 -128.005 277.605 -127.675 ;
        RECT 277.275 -129.365 277.605 -129.035 ;
        RECT 277.275 -130.725 277.605 -130.395 ;
        RECT 277.275 -132.085 277.605 -131.755 ;
        RECT 277.275 -133.445 277.605 -133.115 ;
        RECT 277.275 -134.805 277.605 -134.475 ;
        RECT 277.275 -136.165 277.605 -135.835 ;
        RECT 277.275 -137.525 277.605 -137.195 ;
        RECT 277.275 -138.885 277.605 -138.555 ;
        RECT 277.275 -140.245 277.605 -139.915 ;
        RECT 277.275 -141.605 277.605 -141.275 ;
        RECT 277.275 -142.965 277.605 -142.635 ;
        RECT 277.275 -144.325 277.605 -143.995 ;
        RECT 277.275 -145.685 277.605 -145.355 ;
        RECT 277.275 -147.045 277.605 -146.715 ;
        RECT 277.275 -148.405 277.605 -148.075 ;
        RECT 277.275 -149.765 277.605 -149.435 ;
        RECT 277.275 -151.125 277.605 -150.795 ;
        RECT 277.275 -152.485 277.605 -152.155 ;
        RECT 277.275 -153.845 277.605 -153.515 ;
        RECT 277.275 -155.205 277.605 -154.875 ;
        RECT 277.275 -156.565 277.605 -156.235 ;
        RECT 277.275 -157.925 277.605 -157.595 ;
        RECT 277.275 -159.285 277.605 -158.955 ;
        RECT 277.275 -160.645 277.605 -160.315 ;
        RECT 277.275 -162.005 277.605 -161.675 ;
        RECT 277.275 -163.365 277.605 -163.035 ;
        RECT 277.275 -164.725 277.605 -164.395 ;
        RECT 277.275 -166.085 277.605 -165.755 ;
        RECT 277.275 -167.445 277.605 -167.115 ;
        RECT 277.275 -168.805 277.605 -168.475 ;
        RECT 277.275 -170.165 277.605 -169.835 ;
        RECT 277.275 -171.525 277.605 -171.195 ;
        RECT 277.275 -172.885 277.605 -172.555 ;
        RECT 277.275 -174.245 277.605 -173.915 ;
        RECT 277.275 -175.605 277.605 -175.275 ;
        RECT 277.275 -176.965 277.605 -176.635 ;
        RECT 277.275 -178.325 277.605 -177.995 ;
        RECT 277.275 -180.57 277.605 -179.44 ;
        RECT 277.28 -180.685 277.6 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 277.81 -94.075 278.14 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 278.635 241.32 278.965 242.45 ;
        RECT 278.635 239.195 278.965 239.525 ;
        RECT 278.635 237.835 278.965 238.165 ;
        RECT 278.64 237.16 278.96 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 278.635 -1.525 278.965 -1.195 ;
        RECT 278.635 -2.885 278.965 -2.555 ;
        RECT 278.64 -3.56 278.96 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 279.995 241.32 280.325 242.45 ;
        RECT 279.995 239.195 280.325 239.525 ;
        RECT 279.995 237.835 280.325 238.165 ;
        RECT 280 237.16 280.32 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 279.995 -1.525 280.325 -1.195 ;
        RECT 279.995 -2.885 280.325 -2.555 ;
        RECT 280 -3.56 280.32 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 281.355 241.32 281.685 242.45 ;
        RECT 281.355 239.195 281.685 239.525 ;
        RECT 281.355 237.835 281.685 238.165 ;
        RECT 281.36 237.16 281.68 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 281.355 -1.525 281.685 -1.195 ;
        RECT 281.355 -2.885 281.685 -2.555 ;
        RECT 281.36 -3.56 281.68 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 281.355 -91.285 281.685 -90.955 ;
        RECT 281.355 -92.645 281.685 -92.315 ;
        RECT 281.355 -94.005 281.685 -93.675 ;
        RECT 281.355 -95.365 281.685 -95.035 ;
        RECT 281.355 -96.725 281.685 -96.395 ;
        RECT 281.355 -98.085 281.685 -97.755 ;
        RECT 281.355 -99.445 281.685 -99.115 ;
        RECT 281.355 -100.805 281.685 -100.475 ;
        RECT 281.355 -102.165 281.685 -101.835 ;
        RECT 281.355 -103.525 281.685 -103.195 ;
        RECT 281.355 -104.885 281.685 -104.555 ;
        RECT 281.355 -106.245 281.685 -105.915 ;
        RECT 281.355 -107.605 281.685 -107.275 ;
        RECT 281.355 -108.965 281.685 -108.635 ;
        RECT 281.355 -110.325 281.685 -109.995 ;
        RECT 281.355 -111.685 281.685 -111.355 ;
        RECT 281.355 -113.045 281.685 -112.715 ;
        RECT 281.355 -114.405 281.685 -114.075 ;
        RECT 281.355 -115.765 281.685 -115.435 ;
        RECT 281.355 -117.125 281.685 -116.795 ;
        RECT 281.355 -118.485 281.685 -118.155 ;
        RECT 281.355 -119.845 281.685 -119.515 ;
        RECT 281.355 -121.205 281.685 -120.875 ;
        RECT 281.355 -122.565 281.685 -122.235 ;
        RECT 281.355 -123.925 281.685 -123.595 ;
        RECT 281.355 -125.285 281.685 -124.955 ;
        RECT 281.355 -126.645 281.685 -126.315 ;
        RECT 281.355 -128.005 281.685 -127.675 ;
        RECT 281.355 -129.365 281.685 -129.035 ;
        RECT 281.355 -130.725 281.685 -130.395 ;
        RECT 281.355 -132.085 281.685 -131.755 ;
        RECT 281.355 -133.445 281.685 -133.115 ;
        RECT 281.355 -134.805 281.685 -134.475 ;
        RECT 281.355 -136.165 281.685 -135.835 ;
        RECT 281.355 -137.525 281.685 -137.195 ;
        RECT 281.355 -138.885 281.685 -138.555 ;
        RECT 281.355 -140.245 281.685 -139.915 ;
        RECT 281.355 -141.605 281.685 -141.275 ;
        RECT 281.355 -142.965 281.685 -142.635 ;
        RECT 281.355 -144.325 281.685 -143.995 ;
        RECT 281.355 -145.685 281.685 -145.355 ;
        RECT 281.355 -147.045 281.685 -146.715 ;
        RECT 281.355 -148.405 281.685 -148.075 ;
        RECT 281.355 -149.765 281.685 -149.435 ;
        RECT 281.355 -151.125 281.685 -150.795 ;
        RECT 281.355 -152.485 281.685 -152.155 ;
        RECT 281.355 -153.845 281.685 -153.515 ;
        RECT 281.355 -155.205 281.685 -154.875 ;
        RECT 281.355 -156.565 281.685 -156.235 ;
        RECT 281.355 -157.925 281.685 -157.595 ;
        RECT 281.355 -159.285 281.685 -158.955 ;
        RECT 281.355 -160.645 281.685 -160.315 ;
        RECT 281.355 -162.005 281.685 -161.675 ;
        RECT 281.355 -163.365 281.685 -163.035 ;
        RECT 281.355 -164.725 281.685 -164.395 ;
        RECT 281.355 -166.085 281.685 -165.755 ;
        RECT 281.355 -167.445 281.685 -167.115 ;
        RECT 281.355 -168.805 281.685 -168.475 ;
        RECT 281.355 -170.165 281.685 -169.835 ;
        RECT 281.355 -171.525 281.685 -171.195 ;
        RECT 281.355 -172.885 281.685 -172.555 ;
        RECT 281.355 -174.245 281.685 -173.915 ;
        RECT 281.355 -175.605 281.685 -175.275 ;
        RECT 281.355 -176.965 281.685 -176.635 ;
        RECT 281.355 -178.325 281.685 -177.995 ;
        RECT 281.355 -180.57 281.685 -179.44 ;
        RECT 281.36 -180.685 281.68 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 282.715 241.32 283.045 242.45 ;
        RECT 282.715 239.195 283.045 239.525 ;
        RECT 282.715 237.835 283.045 238.165 ;
        RECT 282.72 237.16 283.04 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 282.715 -95.365 283.045 -95.035 ;
        RECT 282.715 -96.725 283.045 -96.395 ;
        RECT 282.715 -98.085 283.045 -97.755 ;
        RECT 282.715 -99.445 283.045 -99.115 ;
        RECT 282.715 -100.805 283.045 -100.475 ;
        RECT 282.715 -102.165 283.045 -101.835 ;
        RECT 282.715 -103.525 283.045 -103.195 ;
        RECT 282.715 -104.885 283.045 -104.555 ;
        RECT 282.715 -106.245 283.045 -105.915 ;
        RECT 282.715 -107.605 283.045 -107.275 ;
        RECT 282.715 -108.965 283.045 -108.635 ;
        RECT 282.715 -110.325 283.045 -109.995 ;
        RECT 282.715 -111.685 283.045 -111.355 ;
        RECT 282.715 -113.045 283.045 -112.715 ;
        RECT 282.715 -114.405 283.045 -114.075 ;
        RECT 282.715 -115.765 283.045 -115.435 ;
        RECT 282.715 -117.125 283.045 -116.795 ;
        RECT 282.715 -118.485 283.045 -118.155 ;
        RECT 282.715 -119.845 283.045 -119.515 ;
        RECT 282.715 -121.205 283.045 -120.875 ;
        RECT 282.715 -122.565 283.045 -122.235 ;
        RECT 282.715 -123.925 283.045 -123.595 ;
        RECT 282.715 -125.285 283.045 -124.955 ;
        RECT 282.715 -126.645 283.045 -126.315 ;
        RECT 282.715 -128.005 283.045 -127.675 ;
        RECT 282.715 -129.365 283.045 -129.035 ;
        RECT 282.715 -130.725 283.045 -130.395 ;
        RECT 282.715 -132.085 283.045 -131.755 ;
        RECT 282.715 -133.445 283.045 -133.115 ;
        RECT 282.715 -134.805 283.045 -134.475 ;
        RECT 282.715 -136.165 283.045 -135.835 ;
        RECT 282.715 -137.525 283.045 -137.195 ;
        RECT 282.715 -138.885 283.045 -138.555 ;
        RECT 282.715 -140.245 283.045 -139.915 ;
        RECT 282.715 -141.605 283.045 -141.275 ;
        RECT 282.715 -142.965 283.045 -142.635 ;
        RECT 282.715 -144.325 283.045 -143.995 ;
        RECT 282.715 -145.685 283.045 -145.355 ;
        RECT 282.715 -147.045 283.045 -146.715 ;
        RECT 282.715 -148.405 283.045 -148.075 ;
        RECT 282.715 -149.765 283.045 -149.435 ;
        RECT 282.715 -151.125 283.045 -150.795 ;
        RECT 282.715 -152.485 283.045 -152.155 ;
        RECT 282.715 -153.845 283.045 -153.515 ;
        RECT 282.715 -155.205 283.045 -154.875 ;
        RECT 282.715 -156.565 283.045 -156.235 ;
        RECT 282.715 -157.925 283.045 -157.595 ;
        RECT 282.715 -159.285 283.045 -158.955 ;
        RECT 282.715 -160.645 283.045 -160.315 ;
        RECT 282.715 -162.005 283.045 -161.675 ;
        RECT 282.715 -163.365 283.045 -163.035 ;
        RECT 282.715 -164.725 283.045 -164.395 ;
        RECT 282.715 -166.085 283.045 -165.755 ;
        RECT 282.715 -167.445 283.045 -167.115 ;
        RECT 282.715 -168.805 283.045 -168.475 ;
        RECT 282.715 -170.165 283.045 -169.835 ;
        RECT 282.715 -171.525 283.045 -171.195 ;
        RECT 282.715 -172.885 283.045 -172.555 ;
        RECT 282.715 -174.245 283.045 -173.915 ;
        RECT 282.715 -175.605 283.045 -175.275 ;
        RECT 282.715 -176.965 283.045 -176.635 ;
        RECT 282.715 -178.325 283.045 -177.995 ;
        RECT 282.715 -180.57 283.045 -179.44 ;
        RECT 282.72 -180.685 283.04 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 283.91 -94.075 284.24 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 284.075 241.32 284.405 242.45 ;
        RECT 284.075 239.195 284.405 239.525 ;
        RECT 284.075 237.835 284.405 238.165 ;
        RECT 284.08 237.16 284.4 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 285.435 241.32 285.765 242.45 ;
        RECT 285.435 239.195 285.765 239.525 ;
        RECT 285.435 237.835 285.765 238.165 ;
        RECT 285.44 237.16 285.76 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 285.435 -1.525 285.765 -1.195 ;
        RECT 285.435 -2.885 285.765 -2.555 ;
        RECT 285.44 -3.56 285.76 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 285.435 -91.285 285.765 -90.955 ;
        RECT 285.435 -92.645 285.765 -92.315 ;
        RECT 285.435 -94.005 285.765 -93.675 ;
        RECT 285.435 -95.365 285.765 -95.035 ;
        RECT 285.435 -96.725 285.765 -96.395 ;
        RECT 285.435 -98.085 285.765 -97.755 ;
        RECT 285.435 -99.445 285.765 -99.115 ;
        RECT 285.435 -100.805 285.765 -100.475 ;
        RECT 285.435 -102.165 285.765 -101.835 ;
        RECT 285.435 -103.525 285.765 -103.195 ;
        RECT 285.435 -104.885 285.765 -104.555 ;
        RECT 285.435 -106.245 285.765 -105.915 ;
        RECT 285.435 -107.605 285.765 -107.275 ;
        RECT 285.435 -108.965 285.765 -108.635 ;
        RECT 285.435 -110.325 285.765 -109.995 ;
        RECT 285.435 -111.685 285.765 -111.355 ;
        RECT 285.435 -113.045 285.765 -112.715 ;
        RECT 285.435 -114.405 285.765 -114.075 ;
        RECT 285.435 -115.765 285.765 -115.435 ;
        RECT 285.435 -117.125 285.765 -116.795 ;
        RECT 285.435 -118.485 285.765 -118.155 ;
        RECT 285.435 -119.845 285.765 -119.515 ;
        RECT 285.435 -121.205 285.765 -120.875 ;
        RECT 285.435 -122.565 285.765 -122.235 ;
        RECT 285.435 -123.925 285.765 -123.595 ;
        RECT 285.435 -125.285 285.765 -124.955 ;
        RECT 285.435 -126.645 285.765 -126.315 ;
        RECT 285.435 -128.005 285.765 -127.675 ;
        RECT 285.435 -129.365 285.765 -129.035 ;
        RECT 285.435 -130.725 285.765 -130.395 ;
        RECT 285.435 -132.085 285.765 -131.755 ;
        RECT 285.435 -133.445 285.765 -133.115 ;
        RECT 285.435 -134.805 285.765 -134.475 ;
        RECT 285.435 -136.165 285.765 -135.835 ;
        RECT 285.435 -137.525 285.765 -137.195 ;
        RECT 285.435 -138.885 285.765 -138.555 ;
        RECT 285.435 -140.245 285.765 -139.915 ;
        RECT 285.435 -141.605 285.765 -141.275 ;
        RECT 285.435 -142.965 285.765 -142.635 ;
        RECT 285.435 -144.325 285.765 -143.995 ;
        RECT 285.435 -145.685 285.765 -145.355 ;
        RECT 285.435 -147.045 285.765 -146.715 ;
        RECT 285.435 -148.405 285.765 -148.075 ;
        RECT 285.435 -149.765 285.765 -149.435 ;
        RECT 285.435 -151.125 285.765 -150.795 ;
        RECT 285.435 -152.485 285.765 -152.155 ;
        RECT 285.435 -153.845 285.765 -153.515 ;
        RECT 285.435 -155.205 285.765 -154.875 ;
        RECT 285.435 -156.565 285.765 -156.235 ;
        RECT 285.435 -157.925 285.765 -157.595 ;
        RECT 285.435 -159.285 285.765 -158.955 ;
        RECT 285.435 -160.645 285.765 -160.315 ;
        RECT 285.435 -162.005 285.765 -161.675 ;
        RECT 285.435 -163.365 285.765 -163.035 ;
        RECT 285.435 -164.725 285.765 -164.395 ;
        RECT 285.435 -166.085 285.765 -165.755 ;
        RECT 285.435 -167.445 285.765 -167.115 ;
        RECT 285.435 -168.805 285.765 -168.475 ;
        RECT 285.435 -170.165 285.765 -169.835 ;
        RECT 285.435 -171.525 285.765 -171.195 ;
        RECT 285.435 -172.885 285.765 -172.555 ;
        RECT 285.435 -174.245 285.765 -173.915 ;
        RECT 285.435 -175.605 285.765 -175.275 ;
        RECT 285.435 -176.965 285.765 -176.635 ;
        RECT 285.435 -178.325 285.765 -177.995 ;
        RECT 285.435 -180.57 285.765 -179.44 ;
        RECT 285.44 -180.685 285.76 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 286.795 241.32 287.125 242.45 ;
        RECT 286.795 239.195 287.125 239.525 ;
        RECT 286.795 237.835 287.125 238.165 ;
        RECT 286.8 237.16 287.12 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 286.795 -1.525 287.125 -1.195 ;
        RECT 286.795 -2.885 287.125 -2.555 ;
        RECT 286.8 -3.56 287.12 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 288.155 241.32 288.485 242.45 ;
        RECT 288.155 239.195 288.485 239.525 ;
        RECT 288.155 237.835 288.485 238.165 ;
        RECT 288.16 237.16 288.48 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 288.155 -1.525 288.485 -1.195 ;
        RECT 288.155 -2.885 288.485 -2.555 ;
        RECT 288.16 -3.56 288.48 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 288.155 -91.285 288.485 -90.955 ;
        RECT 288.155 -92.645 288.485 -92.315 ;
        RECT 288.155 -94.005 288.485 -93.675 ;
        RECT 288.155 -95.365 288.485 -95.035 ;
        RECT 288.155 -96.725 288.485 -96.395 ;
        RECT 288.155 -98.085 288.485 -97.755 ;
        RECT 288.155 -99.445 288.485 -99.115 ;
        RECT 288.155 -100.805 288.485 -100.475 ;
        RECT 288.155 -102.165 288.485 -101.835 ;
        RECT 288.155 -103.525 288.485 -103.195 ;
        RECT 288.155 -104.885 288.485 -104.555 ;
        RECT 288.155 -106.245 288.485 -105.915 ;
        RECT 288.155 -107.605 288.485 -107.275 ;
        RECT 288.155 -108.965 288.485 -108.635 ;
        RECT 288.155 -110.325 288.485 -109.995 ;
        RECT 288.155 -111.685 288.485 -111.355 ;
        RECT 288.155 -113.045 288.485 -112.715 ;
        RECT 288.155 -114.405 288.485 -114.075 ;
        RECT 288.155 -115.765 288.485 -115.435 ;
        RECT 288.155 -117.125 288.485 -116.795 ;
        RECT 288.155 -118.485 288.485 -118.155 ;
        RECT 288.155 -119.845 288.485 -119.515 ;
        RECT 288.155 -121.205 288.485 -120.875 ;
        RECT 288.155 -122.565 288.485 -122.235 ;
        RECT 288.155 -123.925 288.485 -123.595 ;
        RECT 288.155 -125.285 288.485 -124.955 ;
        RECT 288.155 -126.645 288.485 -126.315 ;
        RECT 288.155 -128.005 288.485 -127.675 ;
        RECT 288.155 -129.365 288.485 -129.035 ;
        RECT 288.155 -130.725 288.485 -130.395 ;
        RECT 288.155 -132.085 288.485 -131.755 ;
        RECT 288.155 -133.445 288.485 -133.115 ;
        RECT 288.155 -134.805 288.485 -134.475 ;
        RECT 288.155 -136.165 288.485 -135.835 ;
        RECT 288.155 -137.525 288.485 -137.195 ;
        RECT 288.155 -138.885 288.485 -138.555 ;
        RECT 288.155 -140.245 288.485 -139.915 ;
        RECT 288.155 -141.605 288.485 -141.275 ;
        RECT 288.155 -142.965 288.485 -142.635 ;
        RECT 288.155 -144.325 288.485 -143.995 ;
        RECT 288.155 -145.685 288.485 -145.355 ;
        RECT 288.155 -147.045 288.485 -146.715 ;
        RECT 288.155 -148.405 288.485 -148.075 ;
        RECT 288.155 -149.765 288.485 -149.435 ;
        RECT 288.155 -151.125 288.485 -150.795 ;
        RECT 288.155 -152.485 288.485 -152.155 ;
        RECT 288.155 -153.845 288.485 -153.515 ;
        RECT 288.155 -155.205 288.485 -154.875 ;
        RECT 288.155 -156.565 288.485 -156.235 ;
        RECT 288.155 -157.925 288.485 -157.595 ;
        RECT 288.155 -159.285 288.485 -158.955 ;
        RECT 288.155 -160.645 288.485 -160.315 ;
        RECT 288.155 -162.005 288.485 -161.675 ;
        RECT 288.155 -163.365 288.485 -163.035 ;
        RECT 288.155 -164.725 288.485 -164.395 ;
        RECT 288.155 -166.085 288.485 -165.755 ;
        RECT 288.155 -167.445 288.485 -167.115 ;
        RECT 288.155 -168.805 288.485 -168.475 ;
        RECT 288.155 -170.165 288.485 -169.835 ;
        RECT 288.155 -171.525 288.485 -171.195 ;
        RECT 288.155 -172.885 288.485 -172.555 ;
        RECT 288.155 -174.245 288.485 -173.915 ;
        RECT 288.155 -175.605 288.485 -175.275 ;
        RECT 288.155 -176.965 288.485 -176.635 ;
        RECT 288.155 -178.325 288.485 -177.995 ;
        RECT 288.155 -180.57 288.485 -179.44 ;
        RECT 288.16 -180.685 288.48 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 289.515 241.32 289.845 242.45 ;
        RECT 289.515 239.195 289.845 239.525 ;
        RECT 289.515 237.835 289.845 238.165 ;
        RECT 289.52 237.16 289.84 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 289.515 -95.365 289.845 -95.035 ;
        RECT 289.515 -96.725 289.845 -96.395 ;
        RECT 289.515 -98.085 289.845 -97.755 ;
        RECT 289.515 -99.445 289.845 -99.115 ;
        RECT 289.515 -100.805 289.845 -100.475 ;
        RECT 289.515 -102.165 289.845 -101.835 ;
        RECT 289.515 -103.525 289.845 -103.195 ;
        RECT 289.515 -104.885 289.845 -104.555 ;
        RECT 289.515 -106.245 289.845 -105.915 ;
        RECT 289.515 -107.605 289.845 -107.275 ;
        RECT 289.515 -108.965 289.845 -108.635 ;
        RECT 289.515 -110.325 289.845 -109.995 ;
        RECT 289.515 -111.685 289.845 -111.355 ;
        RECT 289.515 -113.045 289.845 -112.715 ;
        RECT 289.515 -114.405 289.845 -114.075 ;
        RECT 289.515 -115.765 289.845 -115.435 ;
        RECT 289.515 -117.125 289.845 -116.795 ;
        RECT 289.515 -118.485 289.845 -118.155 ;
        RECT 289.515 -119.845 289.845 -119.515 ;
        RECT 289.515 -121.205 289.845 -120.875 ;
        RECT 289.515 -122.565 289.845 -122.235 ;
        RECT 289.515 -123.925 289.845 -123.595 ;
        RECT 289.515 -125.285 289.845 -124.955 ;
        RECT 289.515 -126.645 289.845 -126.315 ;
        RECT 289.515 -128.005 289.845 -127.675 ;
        RECT 289.515 -129.365 289.845 -129.035 ;
        RECT 289.515 -130.725 289.845 -130.395 ;
        RECT 289.515 -132.085 289.845 -131.755 ;
        RECT 289.515 -133.445 289.845 -133.115 ;
        RECT 289.515 -134.805 289.845 -134.475 ;
        RECT 289.515 -136.165 289.845 -135.835 ;
        RECT 289.515 -137.525 289.845 -137.195 ;
        RECT 289.515 -138.885 289.845 -138.555 ;
        RECT 289.515 -140.245 289.845 -139.915 ;
        RECT 289.515 -141.605 289.845 -141.275 ;
        RECT 289.515 -142.965 289.845 -142.635 ;
        RECT 289.515 -144.325 289.845 -143.995 ;
        RECT 289.515 -145.685 289.845 -145.355 ;
        RECT 289.515 -147.045 289.845 -146.715 ;
        RECT 289.515 -148.405 289.845 -148.075 ;
        RECT 289.515 -149.765 289.845 -149.435 ;
        RECT 289.515 -151.125 289.845 -150.795 ;
        RECT 289.515 -152.485 289.845 -152.155 ;
        RECT 289.515 -153.845 289.845 -153.515 ;
        RECT 289.515 -155.205 289.845 -154.875 ;
        RECT 289.515 -156.565 289.845 -156.235 ;
        RECT 289.515 -157.925 289.845 -157.595 ;
        RECT 289.515 -159.285 289.845 -158.955 ;
        RECT 289.515 -160.645 289.845 -160.315 ;
        RECT 289.515 -162.005 289.845 -161.675 ;
        RECT 289.515 -163.365 289.845 -163.035 ;
        RECT 289.515 -164.725 289.845 -164.395 ;
        RECT 289.515 -166.085 289.845 -165.755 ;
        RECT 289.515 -167.445 289.845 -167.115 ;
        RECT 289.515 -168.805 289.845 -168.475 ;
        RECT 289.515 -170.165 289.845 -169.835 ;
        RECT 289.515 -171.525 289.845 -171.195 ;
        RECT 289.515 -172.885 289.845 -172.555 ;
        RECT 289.515 -174.245 289.845 -173.915 ;
        RECT 289.515 -175.605 289.845 -175.275 ;
        RECT 289.515 -176.965 289.845 -176.635 ;
        RECT 289.515 -178.325 289.845 -177.995 ;
        RECT 289.515 -180.57 289.845 -179.44 ;
        RECT 289.52 -180.685 289.84 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 290.01 -94.075 290.34 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 290.875 241.32 291.205 242.45 ;
        RECT 290.875 239.195 291.205 239.525 ;
        RECT 290.875 237.835 291.205 238.165 ;
        RECT 290.88 237.16 291.2 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 290.875 -1.525 291.205 -1.195 ;
        RECT 290.875 -2.885 291.205 -2.555 ;
        RECT 290.88 -3.56 291.2 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 292.235 241.32 292.565 242.45 ;
        RECT 292.235 239.195 292.565 239.525 ;
        RECT 292.235 237.835 292.565 238.165 ;
        RECT 292.24 237.16 292.56 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 292.235 -1.525 292.565 -1.195 ;
        RECT 292.235 -2.885 292.565 -2.555 ;
        RECT 292.24 -3.56 292.56 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 293.595 241.32 293.925 242.45 ;
        RECT 293.595 239.195 293.925 239.525 ;
        RECT 293.595 237.835 293.925 238.165 ;
        RECT 293.6 237.16 293.92 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 293.595 -1.525 293.925 -1.195 ;
        RECT 293.595 -2.885 293.925 -2.555 ;
        RECT 293.6 -3.56 293.92 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 293.595 -91.285 293.925 -90.955 ;
        RECT 293.595 -92.645 293.925 -92.315 ;
        RECT 293.595 -94.005 293.925 -93.675 ;
        RECT 293.595 -95.365 293.925 -95.035 ;
        RECT 293.595 -96.725 293.925 -96.395 ;
        RECT 293.595 -98.085 293.925 -97.755 ;
        RECT 293.595 -99.445 293.925 -99.115 ;
        RECT 293.595 -100.805 293.925 -100.475 ;
        RECT 293.595 -102.165 293.925 -101.835 ;
        RECT 293.595 -103.525 293.925 -103.195 ;
        RECT 293.595 -104.885 293.925 -104.555 ;
        RECT 293.595 -106.245 293.925 -105.915 ;
        RECT 293.595 -107.605 293.925 -107.275 ;
        RECT 293.595 -108.965 293.925 -108.635 ;
        RECT 293.595 -110.325 293.925 -109.995 ;
        RECT 293.595 -111.685 293.925 -111.355 ;
        RECT 293.595 -113.045 293.925 -112.715 ;
        RECT 293.595 -114.405 293.925 -114.075 ;
        RECT 293.595 -115.765 293.925 -115.435 ;
        RECT 293.595 -117.125 293.925 -116.795 ;
        RECT 293.595 -118.485 293.925 -118.155 ;
        RECT 293.595 -119.845 293.925 -119.515 ;
        RECT 293.595 -121.205 293.925 -120.875 ;
        RECT 293.595 -122.565 293.925 -122.235 ;
        RECT 293.595 -123.925 293.925 -123.595 ;
        RECT 293.595 -125.285 293.925 -124.955 ;
        RECT 293.595 -126.645 293.925 -126.315 ;
        RECT 293.595 -128.005 293.925 -127.675 ;
        RECT 293.595 -129.365 293.925 -129.035 ;
        RECT 293.595 -130.725 293.925 -130.395 ;
        RECT 293.595 -132.085 293.925 -131.755 ;
        RECT 293.595 -133.445 293.925 -133.115 ;
        RECT 293.595 -134.805 293.925 -134.475 ;
        RECT 293.595 -136.165 293.925 -135.835 ;
        RECT 293.595 -137.525 293.925 -137.195 ;
        RECT 293.595 -138.885 293.925 -138.555 ;
        RECT 293.595 -140.245 293.925 -139.915 ;
        RECT 293.595 -141.605 293.925 -141.275 ;
        RECT 293.595 -142.965 293.925 -142.635 ;
        RECT 293.595 -144.325 293.925 -143.995 ;
        RECT 293.595 -145.685 293.925 -145.355 ;
        RECT 293.595 -147.045 293.925 -146.715 ;
        RECT 293.595 -148.405 293.925 -148.075 ;
        RECT 293.595 -149.765 293.925 -149.435 ;
        RECT 293.595 -151.125 293.925 -150.795 ;
        RECT 293.595 -152.485 293.925 -152.155 ;
        RECT 293.595 -153.845 293.925 -153.515 ;
        RECT 293.595 -155.205 293.925 -154.875 ;
        RECT 293.595 -156.565 293.925 -156.235 ;
        RECT 293.595 -157.925 293.925 -157.595 ;
        RECT 293.595 -159.285 293.925 -158.955 ;
        RECT 293.595 -160.645 293.925 -160.315 ;
        RECT 293.595 -162.005 293.925 -161.675 ;
        RECT 293.595 -163.365 293.925 -163.035 ;
        RECT 293.595 -164.725 293.925 -164.395 ;
        RECT 293.595 -166.085 293.925 -165.755 ;
        RECT 293.595 -167.445 293.925 -167.115 ;
        RECT 293.595 -168.805 293.925 -168.475 ;
        RECT 293.595 -170.165 293.925 -169.835 ;
        RECT 293.595 -171.525 293.925 -171.195 ;
        RECT 293.595 -172.885 293.925 -172.555 ;
        RECT 293.595 -174.245 293.925 -173.915 ;
        RECT 293.595 -175.605 293.925 -175.275 ;
        RECT 293.595 -176.965 293.925 -176.635 ;
        RECT 293.595 -178.325 293.925 -177.995 ;
        RECT 293.595 -180.57 293.925 -179.44 ;
        RECT 293.6 -180.685 293.92 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 294.955 241.32 295.285 242.45 ;
        RECT 294.955 239.195 295.285 239.525 ;
        RECT 294.955 237.835 295.285 238.165 ;
        RECT 294.96 237.16 295.28 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 294.955 -95.365 295.285 -95.035 ;
        RECT 294.955 -96.725 295.285 -96.395 ;
        RECT 294.955 -98.085 295.285 -97.755 ;
        RECT 294.955 -99.445 295.285 -99.115 ;
        RECT 294.955 -100.805 295.285 -100.475 ;
        RECT 294.955 -102.165 295.285 -101.835 ;
        RECT 294.955 -103.525 295.285 -103.195 ;
        RECT 294.955 -104.885 295.285 -104.555 ;
        RECT 294.955 -106.245 295.285 -105.915 ;
        RECT 294.955 -107.605 295.285 -107.275 ;
        RECT 294.955 -108.965 295.285 -108.635 ;
        RECT 294.955 -110.325 295.285 -109.995 ;
        RECT 294.955 -111.685 295.285 -111.355 ;
        RECT 294.955 -113.045 295.285 -112.715 ;
        RECT 294.955 -114.405 295.285 -114.075 ;
        RECT 294.955 -115.765 295.285 -115.435 ;
        RECT 294.955 -117.125 295.285 -116.795 ;
        RECT 294.955 -118.485 295.285 -118.155 ;
        RECT 294.955 -119.845 295.285 -119.515 ;
        RECT 294.955 -121.205 295.285 -120.875 ;
        RECT 294.955 -122.565 295.285 -122.235 ;
        RECT 294.955 -123.925 295.285 -123.595 ;
        RECT 294.955 -125.285 295.285 -124.955 ;
        RECT 294.955 -126.645 295.285 -126.315 ;
        RECT 294.955 -128.005 295.285 -127.675 ;
        RECT 294.955 -129.365 295.285 -129.035 ;
        RECT 294.955 -130.725 295.285 -130.395 ;
        RECT 294.955 -132.085 295.285 -131.755 ;
        RECT 294.955 -133.445 295.285 -133.115 ;
        RECT 294.955 -134.805 295.285 -134.475 ;
        RECT 294.955 -136.165 295.285 -135.835 ;
        RECT 294.955 -137.525 295.285 -137.195 ;
        RECT 294.955 -138.885 295.285 -138.555 ;
        RECT 294.955 -140.245 295.285 -139.915 ;
        RECT 294.955 -141.605 295.285 -141.275 ;
        RECT 294.955 -142.965 295.285 -142.635 ;
        RECT 294.955 -144.325 295.285 -143.995 ;
        RECT 294.955 -145.685 295.285 -145.355 ;
        RECT 294.955 -147.045 295.285 -146.715 ;
        RECT 294.955 -148.405 295.285 -148.075 ;
        RECT 294.955 -149.765 295.285 -149.435 ;
        RECT 294.955 -151.125 295.285 -150.795 ;
        RECT 294.955 -152.485 295.285 -152.155 ;
        RECT 294.955 -153.845 295.285 -153.515 ;
        RECT 294.955 -155.205 295.285 -154.875 ;
        RECT 294.955 -156.565 295.285 -156.235 ;
        RECT 294.955 -157.925 295.285 -157.595 ;
        RECT 294.955 -159.285 295.285 -158.955 ;
        RECT 294.955 -160.645 295.285 -160.315 ;
        RECT 294.955 -162.005 295.285 -161.675 ;
        RECT 294.955 -163.365 295.285 -163.035 ;
        RECT 294.955 -164.725 295.285 -164.395 ;
        RECT 294.955 -166.085 295.285 -165.755 ;
        RECT 294.955 -167.445 295.285 -167.115 ;
        RECT 294.955 -168.805 295.285 -168.475 ;
        RECT 294.955 -170.165 295.285 -169.835 ;
        RECT 294.955 -171.525 295.285 -171.195 ;
        RECT 294.955 -172.885 295.285 -172.555 ;
        RECT 294.955 -174.245 295.285 -173.915 ;
        RECT 294.955 -175.605 295.285 -175.275 ;
        RECT 294.955 -176.965 295.285 -176.635 ;
        RECT 294.955 -178.325 295.285 -177.995 ;
        RECT 294.955 -180.57 295.285 -179.44 ;
        RECT 294.96 -180.685 295.28 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 296.11 -94.075 296.44 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 296.315 241.32 296.645 242.45 ;
        RECT 296.315 239.195 296.645 239.525 ;
        RECT 296.315 237.835 296.645 238.165 ;
        RECT 296.32 237.16 296.64 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 297.675 241.32 298.005 242.45 ;
        RECT 297.675 239.195 298.005 239.525 ;
        RECT 297.675 237.835 298.005 238.165 ;
        RECT 297.68 237.16 298 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 297.675 -1.525 298.005 -1.195 ;
        RECT 297.675 -2.885 298.005 -2.555 ;
        RECT 297.68 -3.56 298 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 297.675 -91.285 298.005 -90.955 ;
        RECT 297.675 -92.645 298.005 -92.315 ;
        RECT 297.675 -94.005 298.005 -93.675 ;
        RECT 297.675 -95.365 298.005 -95.035 ;
        RECT 297.675 -96.725 298.005 -96.395 ;
        RECT 297.675 -98.085 298.005 -97.755 ;
        RECT 297.675 -99.445 298.005 -99.115 ;
        RECT 297.675 -100.805 298.005 -100.475 ;
        RECT 297.675 -102.165 298.005 -101.835 ;
        RECT 297.675 -103.525 298.005 -103.195 ;
        RECT 297.675 -104.885 298.005 -104.555 ;
        RECT 297.675 -106.245 298.005 -105.915 ;
        RECT 297.675 -107.605 298.005 -107.275 ;
        RECT 297.675 -108.965 298.005 -108.635 ;
        RECT 297.675 -110.325 298.005 -109.995 ;
        RECT 297.675 -111.685 298.005 -111.355 ;
        RECT 297.675 -113.045 298.005 -112.715 ;
        RECT 297.675 -114.405 298.005 -114.075 ;
        RECT 297.675 -115.765 298.005 -115.435 ;
        RECT 297.675 -117.125 298.005 -116.795 ;
        RECT 297.675 -118.485 298.005 -118.155 ;
        RECT 297.675 -119.845 298.005 -119.515 ;
        RECT 297.675 -121.205 298.005 -120.875 ;
        RECT 297.675 -122.565 298.005 -122.235 ;
        RECT 297.675 -123.925 298.005 -123.595 ;
        RECT 297.675 -125.285 298.005 -124.955 ;
        RECT 297.675 -126.645 298.005 -126.315 ;
        RECT 297.675 -128.005 298.005 -127.675 ;
        RECT 297.675 -129.365 298.005 -129.035 ;
        RECT 297.675 -130.725 298.005 -130.395 ;
        RECT 297.675 -132.085 298.005 -131.755 ;
        RECT 297.675 -133.445 298.005 -133.115 ;
        RECT 297.675 -134.805 298.005 -134.475 ;
        RECT 297.675 -136.165 298.005 -135.835 ;
        RECT 297.675 -137.525 298.005 -137.195 ;
        RECT 297.675 -138.885 298.005 -138.555 ;
        RECT 297.675 -140.245 298.005 -139.915 ;
        RECT 297.675 -141.605 298.005 -141.275 ;
        RECT 297.675 -142.965 298.005 -142.635 ;
        RECT 297.675 -144.325 298.005 -143.995 ;
        RECT 297.675 -145.685 298.005 -145.355 ;
        RECT 297.675 -147.045 298.005 -146.715 ;
        RECT 297.675 -148.405 298.005 -148.075 ;
        RECT 297.675 -149.765 298.005 -149.435 ;
        RECT 297.675 -151.125 298.005 -150.795 ;
        RECT 297.675 -152.485 298.005 -152.155 ;
        RECT 297.675 -153.845 298.005 -153.515 ;
        RECT 297.675 -155.205 298.005 -154.875 ;
        RECT 297.675 -156.565 298.005 -156.235 ;
        RECT 297.675 -157.925 298.005 -157.595 ;
        RECT 297.675 -159.285 298.005 -158.955 ;
        RECT 297.675 -160.645 298.005 -160.315 ;
        RECT 297.675 -162.005 298.005 -161.675 ;
        RECT 297.675 -163.365 298.005 -163.035 ;
        RECT 297.675 -164.725 298.005 -164.395 ;
        RECT 297.675 -166.085 298.005 -165.755 ;
        RECT 297.675 -167.445 298.005 -167.115 ;
        RECT 297.675 -168.805 298.005 -168.475 ;
        RECT 297.675 -170.165 298.005 -169.835 ;
        RECT 297.675 -171.525 298.005 -171.195 ;
        RECT 297.675 -172.885 298.005 -172.555 ;
        RECT 297.675 -174.245 298.005 -173.915 ;
        RECT 297.675 -175.605 298.005 -175.275 ;
        RECT 297.675 -176.965 298.005 -176.635 ;
        RECT 297.675 -178.325 298.005 -177.995 ;
        RECT 297.675 -180.57 298.005 -179.44 ;
        RECT 297.68 -180.685 298 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 299.035 241.32 299.365 242.45 ;
        RECT 299.035 239.195 299.365 239.525 ;
        RECT 299.035 237.835 299.365 238.165 ;
        RECT 299.04 237.16 299.36 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 299.035 -1.525 299.365 -1.195 ;
        RECT 299.035 -2.885 299.365 -2.555 ;
        RECT 299.04 -3.56 299.36 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 300.395 241.32 300.725 242.45 ;
        RECT 300.395 239.195 300.725 239.525 ;
        RECT 300.395 237.835 300.725 238.165 ;
        RECT 300.4 237.16 300.72 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 300.395 -1.525 300.725 -1.195 ;
        RECT 300.395 -2.885 300.725 -2.555 ;
        RECT 300.4 -3.56 300.72 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 300.395 -99.445 300.725 -99.115 ;
        RECT 300.395 -100.805 300.725 -100.475 ;
        RECT 300.395 -102.165 300.725 -101.835 ;
        RECT 300.395 -103.525 300.725 -103.195 ;
        RECT 300.395 -104.885 300.725 -104.555 ;
        RECT 300.395 -106.245 300.725 -105.915 ;
        RECT 300.395 -107.605 300.725 -107.275 ;
        RECT 300.395 -108.965 300.725 -108.635 ;
        RECT 300.395 -110.325 300.725 -109.995 ;
        RECT 300.395 -111.685 300.725 -111.355 ;
        RECT 300.395 -113.045 300.725 -112.715 ;
        RECT 300.395 -114.405 300.725 -114.075 ;
        RECT 300.395 -115.765 300.725 -115.435 ;
        RECT 300.395 -117.125 300.725 -116.795 ;
        RECT 300.395 -118.485 300.725 -118.155 ;
        RECT 300.395 -119.845 300.725 -119.515 ;
        RECT 300.395 -121.205 300.725 -120.875 ;
        RECT 300.395 -122.565 300.725 -122.235 ;
        RECT 300.395 -123.925 300.725 -123.595 ;
        RECT 300.395 -125.285 300.725 -124.955 ;
        RECT 300.395 -126.645 300.725 -126.315 ;
        RECT 300.395 -128.005 300.725 -127.675 ;
        RECT 300.395 -129.365 300.725 -129.035 ;
        RECT 300.395 -130.725 300.725 -130.395 ;
        RECT 300.395 -132.085 300.725 -131.755 ;
        RECT 300.395 -133.445 300.725 -133.115 ;
        RECT 300.395 -134.805 300.725 -134.475 ;
        RECT 300.395 -136.165 300.725 -135.835 ;
        RECT 300.395 -137.525 300.725 -137.195 ;
        RECT 300.395 -138.885 300.725 -138.555 ;
        RECT 300.395 -140.245 300.725 -139.915 ;
        RECT 300.395 -141.605 300.725 -141.275 ;
        RECT 300.395 -142.965 300.725 -142.635 ;
        RECT 300.395 -144.325 300.725 -143.995 ;
        RECT 300.395 -145.685 300.725 -145.355 ;
        RECT 300.395 -147.045 300.725 -146.715 ;
        RECT 300.395 -148.405 300.725 -148.075 ;
        RECT 300.395 -149.765 300.725 -149.435 ;
        RECT 300.395 -151.125 300.725 -150.795 ;
        RECT 300.395 -152.485 300.725 -152.155 ;
        RECT 300.395 -153.845 300.725 -153.515 ;
        RECT 300.395 -155.205 300.725 -154.875 ;
        RECT 300.395 -156.565 300.725 -156.235 ;
        RECT 300.395 -157.925 300.725 -157.595 ;
        RECT 300.395 -159.285 300.725 -158.955 ;
        RECT 300.395 -160.645 300.725 -160.315 ;
        RECT 300.395 -162.005 300.725 -161.675 ;
        RECT 300.395 -163.365 300.725 -163.035 ;
        RECT 300.395 -164.725 300.725 -164.395 ;
        RECT 300.395 -166.085 300.725 -165.755 ;
        RECT 300.395 -167.445 300.725 -167.115 ;
        RECT 300.395 -168.805 300.725 -168.475 ;
        RECT 300.395 -170.165 300.725 -169.835 ;
        RECT 300.395 -171.525 300.725 -171.195 ;
        RECT 300.395 -172.885 300.725 -172.555 ;
        RECT 300.395 -174.245 300.725 -173.915 ;
        RECT 300.395 -175.605 300.725 -175.275 ;
        RECT 300.395 -176.965 300.725 -176.635 ;
        RECT 300.395 -178.325 300.725 -177.995 ;
        RECT 300.395 -180.57 300.725 -179.44 ;
        RECT 300.4 -180.685 300.72 -90.955 ;
        RECT 300.395 -91.285 300.725 -90.955 ;
        RECT 300.395 -92.645 300.725 -92.315 ;
        RECT 300.395 -94.005 300.725 -93.675 ;
        RECT 300.395 -95.365 300.725 -95.035 ;
        RECT 300.395 -96.725 300.725 -96.395 ;
        RECT 300.395 -98.085 300.725 -97.755 ;
    END
    PORT
      LAYER met3 ;
        RECT 236.475 241.32 236.805 242.45 ;
        RECT 236.475 239.195 236.805 239.525 ;
        RECT 236.475 237.835 236.805 238.165 ;
        RECT 236.48 237.16 236.8 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 236.475 -1.525 236.805 -1.195 ;
        RECT 236.475 -2.885 236.805 -2.555 ;
        RECT 236.48 -3.56 236.8 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 237.835 241.32 238.165 242.45 ;
        RECT 237.835 239.195 238.165 239.525 ;
        RECT 237.835 237.835 238.165 238.165 ;
        RECT 237.84 237.16 238.16 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 237.835 -1.525 238.165 -1.195 ;
        RECT 237.835 -2.885 238.165 -2.555 ;
        RECT 237.84 -3.56 238.16 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 239.195 241.32 239.525 242.45 ;
        RECT 239.195 239.195 239.525 239.525 ;
        RECT 239.195 237.835 239.525 238.165 ;
        RECT 239.2 237.16 239.52 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 239.195 -1.525 239.525 -1.195 ;
        RECT 239.195 -2.885 239.525 -2.555 ;
        RECT 239.2 -3.56 239.52 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 239.195 -91.285 239.525 -90.955 ;
        RECT 239.195 -92.645 239.525 -92.315 ;
        RECT 239.195 -94.005 239.525 -93.675 ;
        RECT 239.195 -95.365 239.525 -95.035 ;
        RECT 239.195 -96.725 239.525 -96.395 ;
        RECT 239.195 -98.085 239.525 -97.755 ;
        RECT 239.195 -99.445 239.525 -99.115 ;
        RECT 239.195 -100.805 239.525 -100.475 ;
        RECT 239.195 -102.165 239.525 -101.835 ;
        RECT 239.195 -103.525 239.525 -103.195 ;
        RECT 239.195 -104.885 239.525 -104.555 ;
        RECT 239.195 -106.245 239.525 -105.915 ;
        RECT 239.195 -107.605 239.525 -107.275 ;
        RECT 239.195 -108.965 239.525 -108.635 ;
        RECT 239.195 -110.325 239.525 -109.995 ;
        RECT 239.195 -111.685 239.525 -111.355 ;
        RECT 239.195 -113.045 239.525 -112.715 ;
        RECT 239.195 -114.405 239.525 -114.075 ;
        RECT 239.195 -115.765 239.525 -115.435 ;
        RECT 239.195 -117.125 239.525 -116.795 ;
        RECT 239.195 -118.485 239.525 -118.155 ;
        RECT 239.195 -119.845 239.525 -119.515 ;
        RECT 239.195 -121.205 239.525 -120.875 ;
        RECT 239.195 -122.565 239.525 -122.235 ;
        RECT 239.195 -123.925 239.525 -123.595 ;
        RECT 239.195 -125.285 239.525 -124.955 ;
        RECT 239.195 -126.645 239.525 -126.315 ;
        RECT 239.195 -128.005 239.525 -127.675 ;
        RECT 239.195 -129.365 239.525 -129.035 ;
        RECT 239.195 -130.725 239.525 -130.395 ;
        RECT 239.195 -132.085 239.525 -131.755 ;
        RECT 239.195 -133.445 239.525 -133.115 ;
        RECT 239.195 -134.805 239.525 -134.475 ;
        RECT 239.195 -136.165 239.525 -135.835 ;
        RECT 239.195 -137.525 239.525 -137.195 ;
        RECT 239.195 -138.885 239.525 -138.555 ;
        RECT 239.195 -140.245 239.525 -139.915 ;
        RECT 239.195 -141.605 239.525 -141.275 ;
        RECT 239.195 -142.965 239.525 -142.635 ;
        RECT 239.195 -144.325 239.525 -143.995 ;
        RECT 239.195 -145.685 239.525 -145.355 ;
        RECT 239.195 -147.045 239.525 -146.715 ;
        RECT 239.195 -148.405 239.525 -148.075 ;
        RECT 239.195 -149.765 239.525 -149.435 ;
        RECT 239.195 -151.125 239.525 -150.795 ;
        RECT 239.195 -152.485 239.525 -152.155 ;
        RECT 239.195 -153.845 239.525 -153.515 ;
        RECT 239.195 -155.205 239.525 -154.875 ;
        RECT 239.195 -156.565 239.525 -156.235 ;
        RECT 239.195 -157.925 239.525 -157.595 ;
        RECT 239.195 -159.285 239.525 -158.955 ;
        RECT 239.195 -160.645 239.525 -160.315 ;
        RECT 239.195 -162.005 239.525 -161.675 ;
        RECT 239.195 -163.365 239.525 -163.035 ;
        RECT 239.195 -164.725 239.525 -164.395 ;
        RECT 239.195 -166.085 239.525 -165.755 ;
        RECT 239.195 -167.445 239.525 -167.115 ;
        RECT 239.195 -168.805 239.525 -168.475 ;
        RECT 239.195 -170.165 239.525 -169.835 ;
        RECT 239.195 -171.525 239.525 -171.195 ;
        RECT 239.195 -172.885 239.525 -172.555 ;
        RECT 239.195 -174.245 239.525 -173.915 ;
        RECT 239.195 -175.605 239.525 -175.275 ;
        RECT 239.195 -176.965 239.525 -176.635 ;
        RECT 239.195 -178.325 239.525 -177.995 ;
        RECT 239.195 -180.57 239.525 -179.44 ;
        RECT 239.2 -180.685 239.52 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 240.555 241.32 240.885 242.45 ;
        RECT 240.555 239.195 240.885 239.525 ;
        RECT 240.555 237.835 240.885 238.165 ;
        RECT 240.56 237.16 240.88 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 240.555 -95.365 240.885 -95.035 ;
        RECT 240.555 -96.725 240.885 -96.395 ;
        RECT 240.555 -98.085 240.885 -97.755 ;
        RECT 240.555 -99.445 240.885 -99.115 ;
        RECT 240.555 -100.805 240.885 -100.475 ;
        RECT 240.555 -102.165 240.885 -101.835 ;
        RECT 240.555 -103.525 240.885 -103.195 ;
        RECT 240.555 -104.885 240.885 -104.555 ;
        RECT 240.555 -106.245 240.885 -105.915 ;
        RECT 240.555 -107.605 240.885 -107.275 ;
        RECT 240.555 -108.965 240.885 -108.635 ;
        RECT 240.555 -110.325 240.885 -109.995 ;
        RECT 240.555 -111.685 240.885 -111.355 ;
        RECT 240.555 -113.045 240.885 -112.715 ;
        RECT 240.555 -114.405 240.885 -114.075 ;
        RECT 240.555 -115.765 240.885 -115.435 ;
        RECT 240.555 -117.125 240.885 -116.795 ;
        RECT 240.555 -118.485 240.885 -118.155 ;
        RECT 240.555 -119.845 240.885 -119.515 ;
        RECT 240.555 -121.205 240.885 -120.875 ;
        RECT 240.555 -122.565 240.885 -122.235 ;
        RECT 240.555 -123.925 240.885 -123.595 ;
        RECT 240.555 -125.285 240.885 -124.955 ;
        RECT 240.555 -126.645 240.885 -126.315 ;
        RECT 240.555 -128.005 240.885 -127.675 ;
        RECT 240.555 -129.365 240.885 -129.035 ;
        RECT 240.555 -130.725 240.885 -130.395 ;
        RECT 240.555 -132.085 240.885 -131.755 ;
        RECT 240.555 -133.445 240.885 -133.115 ;
        RECT 240.555 -134.805 240.885 -134.475 ;
        RECT 240.555 -136.165 240.885 -135.835 ;
        RECT 240.555 -137.525 240.885 -137.195 ;
        RECT 240.555 -138.885 240.885 -138.555 ;
        RECT 240.555 -140.245 240.885 -139.915 ;
        RECT 240.555 -141.605 240.885 -141.275 ;
        RECT 240.555 -142.965 240.885 -142.635 ;
        RECT 240.555 -144.325 240.885 -143.995 ;
        RECT 240.555 -145.685 240.885 -145.355 ;
        RECT 240.555 -147.045 240.885 -146.715 ;
        RECT 240.555 -148.405 240.885 -148.075 ;
        RECT 240.555 -149.765 240.885 -149.435 ;
        RECT 240.555 -151.125 240.885 -150.795 ;
        RECT 240.555 -152.485 240.885 -152.155 ;
        RECT 240.555 -153.845 240.885 -153.515 ;
        RECT 240.555 -155.205 240.885 -154.875 ;
        RECT 240.555 -156.565 240.885 -156.235 ;
        RECT 240.555 -157.925 240.885 -157.595 ;
        RECT 240.555 -159.285 240.885 -158.955 ;
        RECT 240.555 -160.645 240.885 -160.315 ;
        RECT 240.555 -162.005 240.885 -161.675 ;
        RECT 240.555 -163.365 240.885 -163.035 ;
        RECT 240.555 -164.725 240.885 -164.395 ;
        RECT 240.555 -166.085 240.885 -165.755 ;
        RECT 240.555 -167.445 240.885 -167.115 ;
        RECT 240.555 -168.805 240.885 -168.475 ;
        RECT 240.555 -170.165 240.885 -169.835 ;
        RECT 240.555 -171.525 240.885 -171.195 ;
        RECT 240.555 -172.885 240.885 -172.555 ;
        RECT 240.555 -174.245 240.885 -173.915 ;
        RECT 240.555 -175.605 240.885 -175.275 ;
        RECT 240.555 -176.965 240.885 -176.635 ;
        RECT 240.555 -178.325 240.885 -177.995 ;
        RECT 240.555 -180.57 240.885 -179.44 ;
        RECT 240.56 -180.685 240.88 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 241.21 -94.075 241.54 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 241.915 241.32 242.245 242.45 ;
        RECT 241.915 239.195 242.245 239.525 ;
        RECT 241.915 237.835 242.245 238.165 ;
        RECT 241.92 237.16 242.24 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 241.915 -1.525 242.245 -1.195 ;
        RECT 241.915 -2.885 242.245 -2.555 ;
        RECT 241.92 -3.56 242.24 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 243.275 241.32 243.605 242.45 ;
        RECT 243.275 239.195 243.605 239.525 ;
        RECT 243.275 237.835 243.605 238.165 ;
        RECT 243.28 237.16 243.6 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 243.275 -1.525 243.605 -1.195 ;
        RECT 243.275 -2.885 243.605 -2.555 ;
        RECT 243.28 -3.56 243.6 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 244.635 241.32 244.965 242.45 ;
        RECT 244.635 239.195 244.965 239.525 ;
        RECT 244.635 237.835 244.965 238.165 ;
        RECT 244.64 237.16 244.96 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 244.635 -1.525 244.965 -1.195 ;
        RECT 244.635 -2.885 244.965 -2.555 ;
        RECT 244.64 -3.56 244.96 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 244.635 -91.285 244.965 -90.955 ;
        RECT 244.635 -92.645 244.965 -92.315 ;
        RECT 244.635 -94.005 244.965 -93.675 ;
        RECT 244.635 -95.365 244.965 -95.035 ;
        RECT 244.635 -96.725 244.965 -96.395 ;
        RECT 244.635 -98.085 244.965 -97.755 ;
        RECT 244.635 -99.445 244.965 -99.115 ;
        RECT 244.635 -100.805 244.965 -100.475 ;
        RECT 244.635 -102.165 244.965 -101.835 ;
        RECT 244.635 -103.525 244.965 -103.195 ;
        RECT 244.635 -104.885 244.965 -104.555 ;
        RECT 244.635 -106.245 244.965 -105.915 ;
        RECT 244.635 -107.605 244.965 -107.275 ;
        RECT 244.635 -108.965 244.965 -108.635 ;
        RECT 244.635 -110.325 244.965 -109.995 ;
        RECT 244.635 -111.685 244.965 -111.355 ;
        RECT 244.635 -113.045 244.965 -112.715 ;
        RECT 244.635 -114.405 244.965 -114.075 ;
        RECT 244.635 -115.765 244.965 -115.435 ;
        RECT 244.635 -117.125 244.965 -116.795 ;
        RECT 244.635 -118.485 244.965 -118.155 ;
        RECT 244.635 -119.845 244.965 -119.515 ;
        RECT 244.635 -121.205 244.965 -120.875 ;
        RECT 244.635 -122.565 244.965 -122.235 ;
        RECT 244.635 -123.925 244.965 -123.595 ;
        RECT 244.635 -125.285 244.965 -124.955 ;
        RECT 244.635 -126.645 244.965 -126.315 ;
        RECT 244.635 -128.005 244.965 -127.675 ;
        RECT 244.635 -129.365 244.965 -129.035 ;
        RECT 244.635 -130.725 244.965 -130.395 ;
        RECT 244.635 -132.085 244.965 -131.755 ;
        RECT 244.635 -133.445 244.965 -133.115 ;
        RECT 244.635 -134.805 244.965 -134.475 ;
        RECT 244.635 -136.165 244.965 -135.835 ;
        RECT 244.635 -137.525 244.965 -137.195 ;
        RECT 244.635 -138.885 244.965 -138.555 ;
        RECT 244.635 -140.245 244.965 -139.915 ;
        RECT 244.635 -141.605 244.965 -141.275 ;
        RECT 244.635 -142.965 244.965 -142.635 ;
        RECT 244.635 -144.325 244.965 -143.995 ;
        RECT 244.635 -145.685 244.965 -145.355 ;
        RECT 244.635 -147.045 244.965 -146.715 ;
        RECT 244.635 -148.405 244.965 -148.075 ;
        RECT 244.635 -149.765 244.965 -149.435 ;
        RECT 244.635 -151.125 244.965 -150.795 ;
        RECT 244.635 -152.485 244.965 -152.155 ;
        RECT 244.635 -153.845 244.965 -153.515 ;
        RECT 244.635 -155.205 244.965 -154.875 ;
        RECT 244.635 -156.565 244.965 -156.235 ;
        RECT 244.635 -157.925 244.965 -157.595 ;
        RECT 244.635 -159.285 244.965 -158.955 ;
        RECT 244.635 -160.645 244.965 -160.315 ;
        RECT 244.635 -162.005 244.965 -161.675 ;
        RECT 244.635 -163.365 244.965 -163.035 ;
        RECT 244.635 -164.725 244.965 -164.395 ;
        RECT 244.635 -166.085 244.965 -165.755 ;
        RECT 244.635 -167.445 244.965 -167.115 ;
        RECT 244.635 -168.805 244.965 -168.475 ;
        RECT 244.635 -170.165 244.965 -169.835 ;
        RECT 244.635 -171.525 244.965 -171.195 ;
        RECT 244.635 -172.885 244.965 -172.555 ;
        RECT 244.635 -174.245 244.965 -173.915 ;
        RECT 244.635 -175.605 244.965 -175.275 ;
        RECT 244.635 -176.965 244.965 -176.635 ;
        RECT 244.635 -178.325 244.965 -177.995 ;
        RECT 244.635 -180.57 244.965 -179.44 ;
        RECT 244.64 -180.685 244.96 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 245.995 241.32 246.325 242.45 ;
        RECT 245.995 239.195 246.325 239.525 ;
        RECT 245.995 237.835 246.325 238.165 ;
        RECT 246 237.16 246.32 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 245.995 -95.365 246.325 -95.035 ;
        RECT 245.995 -96.725 246.325 -96.395 ;
        RECT 245.995 -98.085 246.325 -97.755 ;
        RECT 245.995 -99.445 246.325 -99.115 ;
        RECT 245.995 -100.805 246.325 -100.475 ;
        RECT 245.995 -102.165 246.325 -101.835 ;
        RECT 245.995 -103.525 246.325 -103.195 ;
        RECT 245.995 -104.885 246.325 -104.555 ;
        RECT 245.995 -106.245 246.325 -105.915 ;
        RECT 245.995 -107.605 246.325 -107.275 ;
        RECT 245.995 -108.965 246.325 -108.635 ;
        RECT 245.995 -110.325 246.325 -109.995 ;
        RECT 245.995 -111.685 246.325 -111.355 ;
        RECT 245.995 -113.045 246.325 -112.715 ;
        RECT 245.995 -114.405 246.325 -114.075 ;
        RECT 245.995 -115.765 246.325 -115.435 ;
        RECT 245.995 -117.125 246.325 -116.795 ;
        RECT 245.995 -118.485 246.325 -118.155 ;
        RECT 245.995 -119.845 246.325 -119.515 ;
        RECT 245.995 -121.205 246.325 -120.875 ;
        RECT 245.995 -122.565 246.325 -122.235 ;
        RECT 245.995 -123.925 246.325 -123.595 ;
        RECT 245.995 -125.285 246.325 -124.955 ;
        RECT 245.995 -126.645 246.325 -126.315 ;
        RECT 245.995 -128.005 246.325 -127.675 ;
        RECT 245.995 -129.365 246.325 -129.035 ;
        RECT 245.995 -130.725 246.325 -130.395 ;
        RECT 245.995 -132.085 246.325 -131.755 ;
        RECT 245.995 -133.445 246.325 -133.115 ;
        RECT 245.995 -134.805 246.325 -134.475 ;
        RECT 245.995 -136.165 246.325 -135.835 ;
        RECT 245.995 -137.525 246.325 -137.195 ;
        RECT 245.995 -138.885 246.325 -138.555 ;
        RECT 245.995 -140.245 246.325 -139.915 ;
        RECT 245.995 -141.605 246.325 -141.275 ;
        RECT 245.995 -142.965 246.325 -142.635 ;
        RECT 245.995 -144.325 246.325 -143.995 ;
        RECT 245.995 -145.685 246.325 -145.355 ;
        RECT 245.995 -147.045 246.325 -146.715 ;
        RECT 245.995 -148.405 246.325 -148.075 ;
        RECT 245.995 -149.765 246.325 -149.435 ;
        RECT 245.995 -151.125 246.325 -150.795 ;
        RECT 245.995 -152.485 246.325 -152.155 ;
        RECT 245.995 -153.845 246.325 -153.515 ;
        RECT 245.995 -155.205 246.325 -154.875 ;
        RECT 245.995 -156.565 246.325 -156.235 ;
        RECT 245.995 -157.925 246.325 -157.595 ;
        RECT 245.995 -159.285 246.325 -158.955 ;
        RECT 245.995 -160.645 246.325 -160.315 ;
        RECT 245.995 -162.005 246.325 -161.675 ;
        RECT 245.995 -163.365 246.325 -163.035 ;
        RECT 245.995 -164.725 246.325 -164.395 ;
        RECT 245.995 -166.085 246.325 -165.755 ;
        RECT 245.995 -167.445 246.325 -167.115 ;
        RECT 245.995 -168.805 246.325 -168.475 ;
        RECT 245.995 -170.165 246.325 -169.835 ;
        RECT 245.995 -171.525 246.325 -171.195 ;
        RECT 245.995 -172.885 246.325 -172.555 ;
        RECT 245.995 -174.245 246.325 -173.915 ;
        RECT 245.995 -175.605 246.325 -175.275 ;
        RECT 245.995 -176.965 246.325 -176.635 ;
        RECT 245.995 -178.325 246.325 -177.995 ;
        RECT 245.995 -180.57 246.325 -179.44 ;
        RECT 246 -180.685 246.32 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 247.31 -94.075 247.64 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 247.355 241.32 247.685 242.45 ;
        RECT 247.355 239.195 247.685 239.525 ;
        RECT 247.355 237.835 247.685 238.165 ;
        RECT 247.36 237.16 247.68 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 248.715 241.32 249.045 242.45 ;
        RECT 248.715 239.195 249.045 239.525 ;
        RECT 248.715 237.835 249.045 238.165 ;
        RECT 248.72 237.16 249.04 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 248.715 -1.525 249.045 -1.195 ;
        RECT 248.715 -2.885 249.045 -2.555 ;
        RECT 248.72 -3.56 249.04 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 250.075 241.32 250.405 242.45 ;
        RECT 250.075 239.195 250.405 239.525 ;
        RECT 250.075 237.835 250.405 238.165 ;
        RECT 250.08 237.16 250.4 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 250.075 -1.525 250.405 -1.195 ;
        RECT 250.075 -2.885 250.405 -2.555 ;
        RECT 250.08 -3.56 250.4 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 251.435 241.32 251.765 242.45 ;
        RECT 251.435 239.195 251.765 239.525 ;
        RECT 251.435 237.835 251.765 238.165 ;
        RECT 251.44 237.16 251.76 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 251.435 -1.525 251.765 -1.195 ;
        RECT 251.435 -2.885 251.765 -2.555 ;
        RECT 251.44 -3.56 251.76 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 251.435 -91.285 251.765 -90.955 ;
        RECT 251.435 -92.645 251.765 -92.315 ;
        RECT 251.435 -94.005 251.765 -93.675 ;
        RECT 251.435 -95.365 251.765 -95.035 ;
        RECT 251.435 -96.725 251.765 -96.395 ;
        RECT 251.435 -98.085 251.765 -97.755 ;
        RECT 251.435 -99.445 251.765 -99.115 ;
        RECT 251.435 -100.805 251.765 -100.475 ;
        RECT 251.435 -102.165 251.765 -101.835 ;
        RECT 251.435 -103.525 251.765 -103.195 ;
        RECT 251.435 -104.885 251.765 -104.555 ;
        RECT 251.435 -106.245 251.765 -105.915 ;
        RECT 251.435 -107.605 251.765 -107.275 ;
        RECT 251.435 -108.965 251.765 -108.635 ;
        RECT 251.435 -110.325 251.765 -109.995 ;
        RECT 251.435 -111.685 251.765 -111.355 ;
        RECT 251.435 -113.045 251.765 -112.715 ;
        RECT 251.435 -114.405 251.765 -114.075 ;
        RECT 251.435 -115.765 251.765 -115.435 ;
        RECT 251.435 -117.125 251.765 -116.795 ;
        RECT 251.435 -118.485 251.765 -118.155 ;
        RECT 251.435 -119.845 251.765 -119.515 ;
        RECT 251.435 -121.205 251.765 -120.875 ;
        RECT 251.435 -122.565 251.765 -122.235 ;
        RECT 251.435 -123.925 251.765 -123.595 ;
        RECT 251.435 -125.285 251.765 -124.955 ;
        RECT 251.435 -126.645 251.765 -126.315 ;
        RECT 251.435 -128.005 251.765 -127.675 ;
        RECT 251.435 -129.365 251.765 -129.035 ;
        RECT 251.435 -130.725 251.765 -130.395 ;
        RECT 251.435 -132.085 251.765 -131.755 ;
        RECT 251.435 -133.445 251.765 -133.115 ;
        RECT 251.435 -134.805 251.765 -134.475 ;
        RECT 251.435 -136.165 251.765 -135.835 ;
        RECT 251.435 -137.525 251.765 -137.195 ;
        RECT 251.435 -138.885 251.765 -138.555 ;
        RECT 251.435 -140.245 251.765 -139.915 ;
        RECT 251.435 -141.605 251.765 -141.275 ;
        RECT 251.435 -142.965 251.765 -142.635 ;
        RECT 251.435 -144.325 251.765 -143.995 ;
        RECT 251.435 -145.685 251.765 -145.355 ;
        RECT 251.435 -147.045 251.765 -146.715 ;
        RECT 251.435 -148.405 251.765 -148.075 ;
        RECT 251.435 -149.765 251.765 -149.435 ;
        RECT 251.435 -151.125 251.765 -150.795 ;
        RECT 251.435 -152.485 251.765 -152.155 ;
        RECT 251.435 -153.845 251.765 -153.515 ;
        RECT 251.435 -155.205 251.765 -154.875 ;
        RECT 251.435 -156.565 251.765 -156.235 ;
        RECT 251.435 -157.925 251.765 -157.595 ;
        RECT 251.435 -159.285 251.765 -158.955 ;
        RECT 251.435 -160.645 251.765 -160.315 ;
        RECT 251.435 -162.005 251.765 -161.675 ;
        RECT 251.435 -163.365 251.765 -163.035 ;
        RECT 251.435 -164.725 251.765 -164.395 ;
        RECT 251.435 -166.085 251.765 -165.755 ;
        RECT 251.435 -167.445 251.765 -167.115 ;
        RECT 251.435 -168.805 251.765 -168.475 ;
        RECT 251.435 -170.165 251.765 -169.835 ;
        RECT 251.435 -171.525 251.765 -171.195 ;
        RECT 251.435 -172.885 251.765 -172.555 ;
        RECT 251.435 -174.245 251.765 -173.915 ;
        RECT 251.435 -175.605 251.765 -175.275 ;
        RECT 251.435 -176.965 251.765 -176.635 ;
        RECT 251.435 -178.325 251.765 -177.995 ;
        RECT 251.435 -180.57 251.765 -179.44 ;
        RECT 251.44 -180.685 251.76 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 252.795 241.32 253.125 242.45 ;
        RECT 252.795 239.195 253.125 239.525 ;
        RECT 252.795 237.835 253.125 238.165 ;
        RECT 252.8 237.16 253.12 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 252.795 -95.365 253.125 -95.035 ;
        RECT 252.795 -96.725 253.125 -96.395 ;
        RECT 252.795 -98.085 253.125 -97.755 ;
        RECT 252.795 -99.445 253.125 -99.115 ;
        RECT 252.795 -100.805 253.125 -100.475 ;
        RECT 252.795 -102.165 253.125 -101.835 ;
        RECT 252.795 -103.525 253.125 -103.195 ;
        RECT 252.795 -104.885 253.125 -104.555 ;
        RECT 252.795 -106.245 253.125 -105.915 ;
        RECT 252.795 -107.605 253.125 -107.275 ;
        RECT 252.795 -108.965 253.125 -108.635 ;
        RECT 252.795 -110.325 253.125 -109.995 ;
        RECT 252.795 -111.685 253.125 -111.355 ;
        RECT 252.795 -113.045 253.125 -112.715 ;
        RECT 252.795 -114.405 253.125 -114.075 ;
        RECT 252.795 -115.765 253.125 -115.435 ;
        RECT 252.795 -117.125 253.125 -116.795 ;
        RECT 252.795 -118.485 253.125 -118.155 ;
        RECT 252.795 -119.845 253.125 -119.515 ;
        RECT 252.795 -121.205 253.125 -120.875 ;
        RECT 252.795 -122.565 253.125 -122.235 ;
        RECT 252.795 -123.925 253.125 -123.595 ;
        RECT 252.795 -125.285 253.125 -124.955 ;
        RECT 252.795 -126.645 253.125 -126.315 ;
        RECT 252.795 -128.005 253.125 -127.675 ;
        RECT 252.795 -129.365 253.125 -129.035 ;
        RECT 252.795 -130.725 253.125 -130.395 ;
        RECT 252.795 -132.085 253.125 -131.755 ;
        RECT 252.795 -133.445 253.125 -133.115 ;
        RECT 252.795 -134.805 253.125 -134.475 ;
        RECT 252.795 -136.165 253.125 -135.835 ;
        RECT 252.795 -137.525 253.125 -137.195 ;
        RECT 252.795 -138.885 253.125 -138.555 ;
        RECT 252.795 -140.245 253.125 -139.915 ;
        RECT 252.795 -141.605 253.125 -141.275 ;
        RECT 252.795 -142.965 253.125 -142.635 ;
        RECT 252.795 -144.325 253.125 -143.995 ;
        RECT 252.795 -145.685 253.125 -145.355 ;
        RECT 252.795 -147.045 253.125 -146.715 ;
        RECT 252.795 -148.405 253.125 -148.075 ;
        RECT 252.795 -149.765 253.125 -149.435 ;
        RECT 252.795 -151.125 253.125 -150.795 ;
        RECT 252.795 -152.485 253.125 -152.155 ;
        RECT 252.795 -153.845 253.125 -153.515 ;
        RECT 252.795 -155.205 253.125 -154.875 ;
        RECT 252.795 -156.565 253.125 -156.235 ;
        RECT 252.795 -157.925 253.125 -157.595 ;
        RECT 252.795 -159.285 253.125 -158.955 ;
        RECT 252.795 -160.645 253.125 -160.315 ;
        RECT 252.795 -162.005 253.125 -161.675 ;
        RECT 252.795 -163.365 253.125 -163.035 ;
        RECT 252.795 -164.725 253.125 -164.395 ;
        RECT 252.795 -166.085 253.125 -165.755 ;
        RECT 252.795 -167.445 253.125 -167.115 ;
        RECT 252.795 -168.805 253.125 -168.475 ;
        RECT 252.795 -170.165 253.125 -169.835 ;
        RECT 252.795 -171.525 253.125 -171.195 ;
        RECT 252.795 -172.885 253.125 -172.555 ;
        RECT 252.795 -174.245 253.125 -173.915 ;
        RECT 252.795 -175.605 253.125 -175.275 ;
        RECT 252.795 -176.965 253.125 -176.635 ;
        RECT 252.795 -178.325 253.125 -177.995 ;
        RECT 252.795 -180.57 253.125 -179.44 ;
        RECT 252.8 -180.685 253.12 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 253.41 -94.075 253.74 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 254.155 241.32 254.485 242.45 ;
        RECT 254.155 239.195 254.485 239.525 ;
        RECT 254.155 237.835 254.485 238.165 ;
        RECT 254.16 237.16 254.48 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 254.155 -1.525 254.485 -1.195 ;
        RECT 254.155 -2.885 254.485 -2.555 ;
        RECT 254.16 -3.56 254.48 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 255.515 241.32 255.845 242.45 ;
        RECT 255.515 239.195 255.845 239.525 ;
        RECT 255.515 237.835 255.845 238.165 ;
        RECT 255.52 237.16 255.84 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 255.515 -1.525 255.845 -1.195 ;
        RECT 255.515 -2.885 255.845 -2.555 ;
        RECT 255.52 -3.56 255.84 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 256.875 241.32 257.205 242.45 ;
        RECT 256.875 239.195 257.205 239.525 ;
        RECT 256.875 237.835 257.205 238.165 ;
        RECT 256.88 237.16 257.2 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 256.875 -1.525 257.205 -1.195 ;
        RECT 256.875 -2.885 257.205 -2.555 ;
        RECT 256.88 -3.56 257.2 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 256.875 -91.285 257.205 -90.955 ;
        RECT 256.875 -92.645 257.205 -92.315 ;
        RECT 256.875 -94.005 257.205 -93.675 ;
        RECT 256.875 -95.365 257.205 -95.035 ;
        RECT 256.875 -96.725 257.205 -96.395 ;
        RECT 256.875 -98.085 257.205 -97.755 ;
        RECT 256.875 -99.445 257.205 -99.115 ;
        RECT 256.875 -100.805 257.205 -100.475 ;
        RECT 256.875 -102.165 257.205 -101.835 ;
        RECT 256.875 -103.525 257.205 -103.195 ;
        RECT 256.875 -104.885 257.205 -104.555 ;
        RECT 256.875 -106.245 257.205 -105.915 ;
        RECT 256.875 -107.605 257.205 -107.275 ;
        RECT 256.875 -108.965 257.205 -108.635 ;
        RECT 256.875 -110.325 257.205 -109.995 ;
        RECT 256.875 -111.685 257.205 -111.355 ;
        RECT 256.875 -113.045 257.205 -112.715 ;
        RECT 256.875 -114.405 257.205 -114.075 ;
        RECT 256.875 -115.765 257.205 -115.435 ;
        RECT 256.875 -117.125 257.205 -116.795 ;
        RECT 256.875 -118.485 257.205 -118.155 ;
        RECT 256.875 -119.845 257.205 -119.515 ;
        RECT 256.875 -121.205 257.205 -120.875 ;
        RECT 256.875 -122.565 257.205 -122.235 ;
        RECT 256.875 -123.925 257.205 -123.595 ;
        RECT 256.875 -125.285 257.205 -124.955 ;
        RECT 256.875 -126.645 257.205 -126.315 ;
        RECT 256.875 -128.005 257.205 -127.675 ;
        RECT 256.875 -129.365 257.205 -129.035 ;
        RECT 256.875 -130.725 257.205 -130.395 ;
        RECT 256.875 -132.085 257.205 -131.755 ;
        RECT 256.875 -133.445 257.205 -133.115 ;
        RECT 256.875 -134.805 257.205 -134.475 ;
        RECT 256.875 -136.165 257.205 -135.835 ;
        RECT 256.875 -137.525 257.205 -137.195 ;
        RECT 256.875 -138.885 257.205 -138.555 ;
        RECT 256.875 -140.245 257.205 -139.915 ;
        RECT 256.875 -141.605 257.205 -141.275 ;
        RECT 256.875 -142.965 257.205 -142.635 ;
        RECT 256.875 -144.325 257.205 -143.995 ;
        RECT 256.875 -145.685 257.205 -145.355 ;
        RECT 256.875 -147.045 257.205 -146.715 ;
        RECT 256.875 -148.405 257.205 -148.075 ;
        RECT 256.875 -149.765 257.205 -149.435 ;
        RECT 256.875 -151.125 257.205 -150.795 ;
        RECT 256.875 -152.485 257.205 -152.155 ;
        RECT 256.875 -153.845 257.205 -153.515 ;
        RECT 256.875 -155.205 257.205 -154.875 ;
        RECT 256.875 -156.565 257.205 -156.235 ;
        RECT 256.875 -157.925 257.205 -157.595 ;
        RECT 256.875 -159.285 257.205 -158.955 ;
        RECT 256.875 -160.645 257.205 -160.315 ;
        RECT 256.875 -162.005 257.205 -161.675 ;
        RECT 256.875 -163.365 257.205 -163.035 ;
        RECT 256.875 -164.725 257.205 -164.395 ;
        RECT 256.875 -166.085 257.205 -165.755 ;
        RECT 256.875 -167.445 257.205 -167.115 ;
        RECT 256.875 -168.805 257.205 -168.475 ;
        RECT 256.875 -170.165 257.205 -169.835 ;
        RECT 256.875 -171.525 257.205 -171.195 ;
        RECT 256.875 -172.885 257.205 -172.555 ;
        RECT 256.875 -174.245 257.205 -173.915 ;
        RECT 256.875 -175.605 257.205 -175.275 ;
        RECT 256.875 -176.965 257.205 -176.635 ;
        RECT 256.875 -178.325 257.205 -177.995 ;
        RECT 256.875 -180.57 257.205 -179.44 ;
        RECT 256.88 -180.685 257.2 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 258.235 241.32 258.565 242.45 ;
        RECT 258.235 239.195 258.565 239.525 ;
        RECT 258.235 237.835 258.565 238.165 ;
        RECT 258.24 237.16 258.56 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 258.235 -95.365 258.565 -95.035 ;
        RECT 258.235 -96.725 258.565 -96.395 ;
        RECT 258.235 -98.085 258.565 -97.755 ;
        RECT 258.235 -99.445 258.565 -99.115 ;
        RECT 258.235 -100.805 258.565 -100.475 ;
        RECT 258.235 -102.165 258.565 -101.835 ;
        RECT 258.235 -103.525 258.565 -103.195 ;
        RECT 258.235 -104.885 258.565 -104.555 ;
        RECT 258.235 -106.245 258.565 -105.915 ;
        RECT 258.235 -107.605 258.565 -107.275 ;
        RECT 258.235 -108.965 258.565 -108.635 ;
        RECT 258.235 -110.325 258.565 -109.995 ;
        RECT 258.235 -111.685 258.565 -111.355 ;
        RECT 258.235 -113.045 258.565 -112.715 ;
        RECT 258.235 -114.405 258.565 -114.075 ;
        RECT 258.235 -115.765 258.565 -115.435 ;
        RECT 258.235 -117.125 258.565 -116.795 ;
        RECT 258.235 -118.485 258.565 -118.155 ;
        RECT 258.235 -119.845 258.565 -119.515 ;
        RECT 258.235 -121.205 258.565 -120.875 ;
        RECT 258.235 -122.565 258.565 -122.235 ;
        RECT 258.235 -123.925 258.565 -123.595 ;
        RECT 258.235 -125.285 258.565 -124.955 ;
        RECT 258.235 -126.645 258.565 -126.315 ;
        RECT 258.235 -128.005 258.565 -127.675 ;
        RECT 258.235 -129.365 258.565 -129.035 ;
        RECT 258.235 -130.725 258.565 -130.395 ;
        RECT 258.235 -132.085 258.565 -131.755 ;
        RECT 258.235 -133.445 258.565 -133.115 ;
        RECT 258.235 -134.805 258.565 -134.475 ;
        RECT 258.235 -136.165 258.565 -135.835 ;
        RECT 258.235 -137.525 258.565 -137.195 ;
        RECT 258.235 -138.885 258.565 -138.555 ;
        RECT 258.235 -140.245 258.565 -139.915 ;
        RECT 258.235 -141.605 258.565 -141.275 ;
        RECT 258.235 -142.965 258.565 -142.635 ;
        RECT 258.235 -144.325 258.565 -143.995 ;
        RECT 258.235 -145.685 258.565 -145.355 ;
        RECT 258.235 -147.045 258.565 -146.715 ;
        RECT 258.235 -148.405 258.565 -148.075 ;
        RECT 258.235 -149.765 258.565 -149.435 ;
        RECT 258.235 -151.125 258.565 -150.795 ;
        RECT 258.235 -152.485 258.565 -152.155 ;
        RECT 258.235 -153.845 258.565 -153.515 ;
        RECT 258.235 -155.205 258.565 -154.875 ;
        RECT 258.235 -156.565 258.565 -156.235 ;
        RECT 258.235 -157.925 258.565 -157.595 ;
        RECT 258.235 -159.285 258.565 -158.955 ;
        RECT 258.235 -160.645 258.565 -160.315 ;
        RECT 258.235 -162.005 258.565 -161.675 ;
        RECT 258.235 -163.365 258.565 -163.035 ;
        RECT 258.235 -164.725 258.565 -164.395 ;
        RECT 258.235 -166.085 258.565 -165.755 ;
        RECT 258.235 -167.445 258.565 -167.115 ;
        RECT 258.235 -168.805 258.565 -168.475 ;
        RECT 258.235 -170.165 258.565 -169.835 ;
        RECT 258.235 -171.525 258.565 -171.195 ;
        RECT 258.235 -172.885 258.565 -172.555 ;
        RECT 258.235 -174.245 258.565 -173.915 ;
        RECT 258.235 -175.605 258.565 -175.275 ;
        RECT 258.235 -176.965 258.565 -176.635 ;
        RECT 258.235 -178.325 258.565 -177.995 ;
        RECT 258.235 -180.57 258.565 -179.44 ;
        RECT 258.24 -180.685 258.56 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 259.51 -94.075 259.84 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 259.595 241.32 259.925 242.45 ;
        RECT 259.595 239.195 259.925 239.525 ;
        RECT 259.595 237.835 259.925 238.165 ;
        RECT 259.6 237.16 259.92 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 260.955 241.32 261.285 242.45 ;
        RECT 260.955 239.195 261.285 239.525 ;
        RECT 260.955 237.835 261.285 238.165 ;
        RECT 260.96 237.16 261.28 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 260.955 -1.525 261.285 -1.195 ;
        RECT 260.955 -2.885 261.285 -2.555 ;
        RECT 260.96 -3.56 261.28 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 260.955 -91.285 261.285 -90.955 ;
        RECT 260.955 -92.645 261.285 -92.315 ;
        RECT 260.955 -94.005 261.285 -93.675 ;
        RECT 260.955 -95.365 261.285 -95.035 ;
        RECT 260.955 -96.725 261.285 -96.395 ;
        RECT 260.955 -98.085 261.285 -97.755 ;
        RECT 260.955 -99.445 261.285 -99.115 ;
        RECT 260.955 -100.805 261.285 -100.475 ;
        RECT 260.955 -102.165 261.285 -101.835 ;
        RECT 260.955 -103.525 261.285 -103.195 ;
        RECT 260.955 -104.885 261.285 -104.555 ;
        RECT 260.955 -106.245 261.285 -105.915 ;
        RECT 260.955 -107.605 261.285 -107.275 ;
        RECT 260.955 -108.965 261.285 -108.635 ;
        RECT 260.955 -110.325 261.285 -109.995 ;
        RECT 260.955 -111.685 261.285 -111.355 ;
        RECT 260.955 -113.045 261.285 -112.715 ;
        RECT 260.955 -114.405 261.285 -114.075 ;
        RECT 260.955 -115.765 261.285 -115.435 ;
        RECT 260.955 -117.125 261.285 -116.795 ;
        RECT 260.955 -118.485 261.285 -118.155 ;
        RECT 260.955 -119.845 261.285 -119.515 ;
        RECT 260.955 -121.205 261.285 -120.875 ;
        RECT 260.955 -122.565 261.285 -122.235 ;
        RECT 260.955 -123.925 261.285 -123.595 ;
        RECT 260.955 -125.285 261.285 -124.955 ;
        RECT 260.955 -126.645 261.285 -126.315 ;
        RECT 260.955 -128.005 261.285 -127.675 ;
        RECT 260.955 -129.365 261.285 -129.035 ;
        RECT 260.955 -130.725 261.285 -130.395 ;
        RECT 260.955 -132.085 261.285 -131.755 ;
        RECT 260.955 -133.445 261.285 -133.115 ;
        RECT 260.955 -134.805 261.285 -134.475 ;
        RECT 260.955 -136.165 261.285 -135.835 ;
        RECT 260.955 -137.525 261.285 -137.195 ;
        RECT 260.955 -138.885 261.285 -138.555 ;
        RECT 260.955 -140.245 261.285 -139.915 ;
        RECT 260.955 -141.605 261.285 -141.275 ;
        RECT 260.955 -142.965 261.285 -142.635 ;
        RECT 260.955 -144.325 261.285 -143.995 ;
        RECT 260.955 -145.685 261.285 -145.355 ;
        RECT 260.955 -147.045 261.285 -146.715 ;
        RECT 260.955 -148.405 261.285 -148.075 ;
        RECT 260.955 -149.765 261.285 -149.435 ;
        RECT 260.955 -151.125 261.285 -150.795 ;
        RECT 260.955 -152.485 261.285 -152.155 ;
        RECT 260.955 -153.845 261.285 -153.515 ;
        RECT 260.955 -155.205 261.285 -154.875 ;
        RECT 260.955 -156.565 261.285 -156.235 ;
        RECT 260.955 -157.925 261.285 -157.595 ;
        RECT 260.955 -159.285 261.285 -158.955 ;
        RECT 260.955 -160.645 261.285 -160.315 ;
        RECT 260.955 -162.005 261.285 -161.675 ;
        RECT 260.955 -163.365 261.285 -163.035 ;
        RECT 260.955 -164.725 261.285 -164.395 ;
        RECT 260.955 -166.085 261.285 -165.755 ;
        RECT 260.955 -167.445 261.285 -167.115 ;
        RECT 260.955 -168.805 261.285 -168.475 ;
        RECT 260.955 -170.165 261.285 -169.835 ;
        RECT 260.955 -171.525 261.285 -171.195 ;
        RECT 260.955 -172.885 261.285 -172.555 ;
        RECT 260.955 -174.245 261.285 -173.915 ;
        RECT 260.955 -175.605 261.285 -175.275 ;
        RECT 260.955 -176.965 261.285 -176.635 ;
        RECT 260.955 -178.325 261.285 -177.995 ;
        RECT 260.955 -180.57 261.285 -179.44 ;
        RECT 260.96 -180.685 261.28 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 262.315 241.32 262.645 242.45 ;
        RECT 262.315 239.195 262.645 239.525 ;
        RECT 262.315 237.835 262.645 238.165 ;
        RECT 262.32 237.16 262.64 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 262.315 -1.525 262.645 -1.195 ;
        RECT 262.315 -2.885 262.645 -2.555 ;
        RECT 262.32 -3.56 262.64 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 263.675 241.32 264.005 242.45 ;
        RECT 263.675 239.195 264.005 239.525 ;
        RECT 263.675 237.835 264.005 238.165 ;
        RECT 263.68 237.16 264 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 263.675 -1.525 264.005 -1.195 ;
        RECT 263.675 -2.885 264.005 -2.555 ;
        RECT 263.68 -3.56 264 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 263.675 -91.285 264.005 -90.955 ;
        RECT 263.675 -92.645 264.005 -92.315 ;
        RECT 263.675 -94.005 264.005 -93.675 ;
        RECT 263.675 -95.365 264.005 -95.035 ;
        RECT 263.675 -96.725 264.005 -96.395 ;
        RECT 263.675 -98.085 264.005 -97.755 ;
        RECT 263.675 -99.445 264.005 -99.115 ;
        RECT 263.675 -100.805 264.005 -100.475 ;
        RECT 263.675 -102.165 264.005 -101.835 ;
        RECT 263.675 -103.525 264.005 -103.195 ;
        RECT 263.675 -104.885 264.005 -104.555 ;
        RECT 263.675 -106.245 264.005 -105.915 ;
        RECT 263.675 -107.605 264.005 -107.275 ;
        RECT 263.675 -108.965 264.005 -108.635 ;
        RECT 263.675 -110.325 264.005 -109.995 ;
        RECT 263.675 -111.685 264.005 -111.355 ;
        RECT 263.675 -113.045 264.005 -112.715 ;
        RECT 263.675 -114.405 264.005 -114.075 ;
        RECT 263.675 -115.765 264.005 -115.435 ;
        RECT 263.675 -117.125 264.005 -116.795 ;
        RECT 263.675 -118.485 264.005 -118.155 ;
        RECT 263.675 -119.845 264.005 -119.515 ;
        RECT 263.675 -121.205 264.005 -120.875 ;
        RECT 263.675 -122.565 264.005 -122.235 ;
        RECT 263.675 -123.925 264.005 -123.595 ;
        RECT 263.675 -125.285 264.005 -124.955 ;
        RECT 263.675 -126.645 264.005 -126.315 ;
        RECT 263.675 -128.005 264.005 -127.675 ;
        RECT 263.675 -129.365 264.005 -129.035 ;
        RECT 263.675 -130.725 264.005 -130.395 ;
        RECT 263.675 -132.085 264.005 -131.755 ;
        RECT 263.675 -133.445 264.005 -133.115 ;
        RECT 263.675 -134.805 264.005 -134.475 ;
        RECT 263.675 -136.165 264.005 -135.835 ;
        RECT 263.675 -137.525 264.005 -137.195 ;
        RECT 263.675 -138.885 264.005 -138.555 ;
        RECT 263.675 -140.245 264.005 -139.915 ;
        RECT 263.675 -141.605 264.005 -141.275 ;
        RECT 263.675 -142.965 264.005 -142.635 ;
        RECT 263.675 -144.325 264.005 -143.995 ;
        RECT 263.675 -145.685 264.005 -145.355 ;
        RECT 263.675 -147.045 264.005 -146.715 ;
        RECT 263.675 -148.405 264.005 -148.075 ;
        RECT 263.675 -149.765 264.005 -149.435 ;
        RECT 263.675 -151.125 264.005 -150.795 ;
        RECT 263.675 -152.485 264.005 -152.155 ;
        RECT 263.675 -153.845 264.005 -153.515 ;
        RECT 263.675 -155.205 264.005 -154.875 ;
        RECT 263.675 -156.565 264.005 -156.235 ;
        RECT 263.675 -157.925 264.005 -157.595 ;
        RECT 263.675 -159.285 264.005 -158.955 ;
        RECT 263.675 -160.645 264.005 -160.315 ;
        RECT 263.675 -162.005 264.005 -161.675 ;
        RECT 263.675 -163.365 264.005 -163.035 ;
        RECT 263.675 -164.725 264.005 -164.395 ;
        RECT 263.675 -166.085 264.005 -165.755 ;
        RECT 263.675 -167.445 264.005 -167.115 ;
        RECT 263.675 -168.805 264.005 -168.475 ;
        RECT 263.675 -170.165 264.005 -169.835 ;
        RECT 263.675 -171.525 264.005 -171.195 ;
        RECT 263.675 -172.885 264.005 -172.555 ;
        RECT 263.675 -174.245 264.005 -173.915 ;
        RECT 263.675 -175.605 264.005 -175.275 ;
        RECT 263.675 -176.965 264.005 -176.635 ;
        RECT 263.675 -178.325 264.005 -177.995 ;
        RECT 263.675 -180.57 264.005 -179.44 ;
        RECT 263.68 -180.685 264 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 265.035 241.32 265.365 242.45 ;
        RECT 265.035 239.195 265.365 239.525 ;
        RECT 265.035 237.835 265.365 238.165 ;
        RECT 265.04 237.16 265.36 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 265.035 -95.365 265.365 -95.035 ;
        RECT 265.035 -96.725 265.365 -96.395 ;
        RECT 265.035 -98.085 265.365 -97.755 ;
        RECT 265.035 -99.445 265.365 -99.115 ;
        RECT 265.035 -100.805 265.365 -100.475 ;
        RECT 265.035 -102.165 265.365 -101.835 ;
        RECT 265.035 -103.525 265.365 -103.195 ;
        RECT 265.035 -104.885 265.365 -104.555 ;
        RECT 265.035 -106.245 265.365 -105.915 ;
        RECT 265.035 -107.605 265.365 -107.275 ;
        RECT 265.035 -108.965 265.365 -108.635 ;
        RECT 265.035 -110.325 265.365 -109.995 ;
        RECT 265.035 -111.685 265.365 -111.355 ;
        RECT 265.035 -113.045 265.365 -112.715 ;
        RECT 265.035 -114.405 265.365 -114.075 ;
        RECT 265.035 -115.765 265.365 -115.435 ;
        RECT 265.035 -117.125 265.365 -116.795 ;
        RECT 265.035 -118.485 265.365 -118.155 ;
        RECT 265.035 -119.845 265.365 -119.515 ;
        RECT 265.035 -121.205 265.365 -120.875 ;
        RECT 265.035 -122.565 265.365 -122.235 ;
        RECT 265.035 -123.925 265.365 -123.595 ;
        RECT 265.035 -125.285 265.365 -124.955 ;
        RECT 265.035 -126.645 265.365 -126.315 ;
        RECT 265.035 -128.005 265.365 -127.675 ;
        RECT 265.035 -129.365 265.365 -129.035 ;
        RECT 265.035 -130.725 265.365 -130.395 ;
        RECT 265.035 -132.085 265.365 -131.755 ;
        RECT 265.035 -133.445 265.365 -133.115 ;
        RECT 265.035 -134.805 265.365 -134.475 ;
        RECT 265.035 -136.165 265.365 -135.835 ;
        RECT 265.035 -137.525 265.365 -137.195 ;
        RECT 265.035 -138.885 265.365 -138.555 ;
        RECT 265.035 -140.245 265.365 -139.915 ;
        RECT 265.035 -141.605 265.365 -141.275 ;
        RECT 265.035 -142.965 265.365 -142.635 ;
        RECT 265.035 -144.325 265.365 -143.995 ;
        RECT 265.035 -145.685 265.365 -145.355 ;
        RECT 265.035 -147.045 265.365 -146.715 ;
        RECT 265.035 -148.405 265.365 -148.075 ;
        RECT 265.035 -149.765 265.365 -149.435 ;
        RECT 265.035 -151.125 265.365 -150.795 ;
        RECT 265.035 -152.485 265.365 -152.155 ;
        RECT 265.035 -153.845 265.365 -153.515 ;
        RECT 265.035 -155.205 265.365 -154.875 ;
        RECT 265.035 -156.565 265.365 -156.235 ;
        RECT 265.035 -157.925 265.365 -157.595 ;
        RECT 265.035 -159.285 265.365 -158.955 ;
        RECT 265.035 -160.645 265.365 -160.315 ;
        RECT 265.035 -162.005 265.365 -161.675 ;
        RECT 265.035 -163.365 265.365 -163.035 ;
        RECT 265.035 -164.725 265.365 -164.395 ;
        RECT 265.035 -166.085 265.365 -165.755 ;
        RECT 265.035 -167.445 265.365 -167.115 ;
        RECT 265.035 -168.805 265.365 -168.475 ;
        RECT 265.035 -170.165 265.365 -169.835 ;
        RECT 265.035 -171.525 265.365 -171.195 ;
        RECT 265.035 -172.885 265.365 -172.555 ;
        RECT 265.035 -174.245 265.365 -173.915 ;
        RECT 265.035 -175.605 265.365 -175.275 ;
        RECT 265.035 -176.965 265.365 -176.635 ;
        RECT 265.035 -178.325 265.365 -177.995 ;
        RECT 265.035 -180.57 265.365 -179.44 ;
        RECT 265.04 -180.685 265.36 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 265.61 -94.075 265.94 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 266.395 241.32 266.725 242.45 ;
        RECT 266.395 239.195 266.725 239.525 ;
        RECT 266.395 237.835 266.725 238.165 ;
        RECT 266.4 237.16 266.72 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 266.395 -1.525 266.725 -1.195 ;
        RECT 266.395 -2.885 266.725 -2.555 ;
        RECT 266.4 -3.56 266.72 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 267.755 241.32 268.085 242.45 ;
        RECT 267.755 239.195 268.085 239.525 ;
        RECT 267.755 237.835 268.085 238.165 ;
        RECT 267.76 237.16 268.08 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 267.755 -1.525 268.085 -1.195 ;
        RECT 267.755 -2.885 268.085 -2.555 ;
        RECT 267.76 -3.56 268.08 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 269.115 241.32 269.445 242.45 ;
        RECT 269.115 239.195 269.445 239.525 ;
        RECT 269.115 237.835 269.445 238.165 ;
        RECT 269.12 237.16 269.44 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 269.115 -1.525 269.445 -1.195 ;
        RECT 269.115 -2.885 269.445 -2.555 ;
        RECT 269.12 -3.56 269.44 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 269.115 -102.165 269.445 -101.835 ;
        RECT 269.115 -103.525 269.445 -103.195 ;
        RECT 269.115 -104.885 269.445 -104.555 ;
        RECT 269.115 -106.245 269.445 -105.915 ;
        RECT 269.115 -107.605 269.445 -107.275 ;
        RECT 269.115 -108.965 269.445 -108.635 ;
        RECT 269.115 -110.325 269.445 -109.995 ;
        RECT 269.115 -111.685 269.445 -111.355 ;
        RECT 269.115 -113.045 269.445 -112.715 ;
        RECT 269.115 -114.405 269.445 -114.075 ;
        RECT 269.115 -115.765 269.445 -115.435 ;
        RECT 269.115 -117.125 269.445 -116.795 ;
        RECT 269.115 -118.485 269.445 -118.155 ;
        RECT 269.115 -119.845 269.445 -119.515 ;
        RECT 269.115 -121.205 269.445 -120.875 ;
        RECT 269.115 -122.565 269.445 -122.235 ;
        RECT 269.115 -123.925 269.445 -123.595 ;
        RECT 269.115 -125.285 269.445 -124.955 ;
        RECT 269.115 -126.645 269.445 -126.315 ;
        RECT 269.115 -128.005 269.445 -127.675 ;
        RECT 269.115 -129.365 269.445 -129.035 ;
        RECT 269.115 -130.725 269.445 -130.395 ;
        RECT 269.115 -132.085 269.445 -131.755 ;
        RECT 269.115 -133.445 269.445 -133.115 ;
        RECT 269.115 -134.805 269.445 -134.475 ;
        RECT 269.115 -136.165 269.445 -135.835 ;
        RECT 269.115 -137.525 269.445 -137.195 ;
        RECT 269.115 -138.885 269.445 -138.555 ;
        RECT 269.115 -140.245 269.445 -139.915 ;
        RECT 269.115 -141.605 269.445 -141.275 ;
        RECT 269.115 -142.965 269.445 -142.635 ;
        RECT 269.115 -144.325 269.445 -143.995 ;
        RECT 269.115 -145.685 269.445 -145.355 ;
        RECT 269.115 -147.045 269.445 -146.715 ;
        RECT 269.115 -148.405 269.445 -148.075 ;
        RECT 269.115 -149.765 269.445 -149.435 ;
        RECT 269.115 -151.125 269.445 -150.795 ;
        RECT 269.115 -152.485 269.445 -152.155 ;
        RECT 269.115 -153.845 269.445 -153.515 ;
        RECT 269.115 -155.205 269.445 -154.875 ;
        RECT 269.115 -156.565 269.445 -156.235 ;
        RECT 269.115 -157.925 269.445 -157.595 ;
        RECT 269.115 -159.285 269.445 -158.955 ;
        RECT 269.115 -160.645 269.445 -160.315 ;
        RECT 269.115 -162.005 269.445 -161.675 ;
        RECT 269.115 -163.365 269.445 -163.035 ;
        RECT 269.115 -164.725 269.445 -164.395 ;
        RECT 269.115 -166.085 269.445 -165.755 ;
        RECT 269.115 -167.445 269.445 -167.115 ;
        RECT 269.115 -168.805 269.445 -168.475 ;
        RECT 269.115 -170.165 269.445 -169.835 ;
        RECT 269.115 -171.525 269.445 -171.195 ;
        RECT 269.115 -172.885 269.445 -172.555 ;
        RECT 269.115 -174.245 269.445 -173.915 ;
        RECT 269.115 -175.605 269.445 -175.275 ;
        RECT 269.115 -176.965 269.445 -176.635 ;
        RECT 269.115 -178.325 269.445 -177.995 ;
        RECT 269.115 -180.57 269.445 -179.44 ;
        RECT 269.12 -180.685 269.44 -90.955 ;
        RECT 269.115 -91.285 269.445 -90.955 ;
        RECT 269.115 -92.645 269.445 -92.315 ;
        RECT 269.115 -94.005 269.445 -93.675 ;
        RECT 269.115 -95.365 269.445 -95.035 ;
        RECT 269.115 -96.725 269.445 -96.395 ;
        RECT 269.115 -98.085 269.445 -97.755 ;
        RECT 269.115 -99.445 269.445 -99.115 ;
        RECT 269.115 -100.805 269.445 -100.475 ;
    END
    PORT
      LAYER met3 ;
        RECT 204.61 -94.075 204.94 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 205.195 241.32 205.525 242.45 ;
        RECT 205.195 239.195 205.525 239.525 ;
        RECT 205.195 237.835 205.525 238.165 ;
        RECT 205.2 237.16 205.52 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 206.555 241.32 206.885 242.45 ;
        RECT 206.555 239.195 206.885 239.525 ;
        RECT 206.555 237.835 206.885 238.165 ;
        RECT 206.56 237.16 206.88 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 206.555 -1.525 206.885 -1.195 ;
        RECT 206.555 -2.885 206.885 -2.555 ;
        RECT 206.56 -3.56 206.88 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 207.915 241.32 208.245 242.45 ;
        RECT 207.915 239.195 208.245 239.525 ;
        RECT 207.915 237.835 208.245 238.165 ;
        RECT 207.92 237.16 208.24 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 207.915 -1.525 208.245 -1.195 ;
        RECT 207.915 -2.885 208.245 -2.555 ;
        RECT 207.92 -3.56 208.24 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 207.915 -91.285 208.245 -90.955 ;
        RECT 207.915 -92.645 208.245 -92.315 ;
        RECT 207.915 -94.005 208.245 -93.675 ;
        RECT 207.915 -95.365 208.245 -95.035 ;
        RECT 207.915 -96.725 208.245 -96.395 ;
        RECT 207.915 -98.085 208.245 -97.755 ;
        RECT 207.915 -99.445 208.245 -99.115 ;
        RECT 207.915 -100.805 208.245 -100.475 ;
        RECT 207.915 -102.165 208.245 -101.835 ;
        RECT 207.915 -103.525 208.245 -103.195 ;
        RECT 207.915 -104.885 208.245 -104.555 ;
        RECT 207.915 -106.245 208.245 -105.915 ;
        RECT 207.915 -107.605 208.245 -107.275 ;
        RECT 207.915 -108.965 208.245 -108.635 ;
        RECT 207.915 -110.325 208.245 -109.995 ;
        RECT 207.915 -111.685 208.245 -111.355 ;
        RECT 207.915 -113.045 208.245 -112.715 ;
        RECT 207.915 -114.405 208.245 -114.075 ;
        RECT 207.915 -115.765 208.245 -115.435 ;
        RECT 207.915 -117.125 208.245 -116.795 ;
        RECT 207.915 -118.485 208.245 -118.155 ;
        RECT 207.915 -119.845 208.245 -119.515 ;
        RECT 207.915 -121.205 208.245 -120.875 ;
        RECT 207.915 -122.565 208.245 -122.235 ;
        RECT 207.915 -123.925 208.245 -123.595 ;
        RECT 207.915 -125.285 208.245 -124.955 ;
        RECT 207.915 -126.645 208.245 -126.315 ;
        RECT 207.915 -128.005 208.245 -127.675 ;
        RECT 207.915 -129.365 208.245 -129.035 ;
        RECT 207.915 -130.725 208.245 -130.395 ;
        RECT 207.915 -132.085 208.245 -131.755 ;
        RECT 207.915 -133.445 208.245 -133.115 ;
        RECT 207.915 -134.805 208.245 -134.475 ;
        RECT 207.915 -136.165 208.245 -135.835 ;
        RECT 207.915 -137.525 208.245 -137.195 ;
        RECT 207.915 -138.885 208.245 -138.555 ;
        RECT 207.915 -140.245 208.245 -139.915 ;
        RECT 207.915 -141.605 208.245 -141.275 ;
        RECT 207.915 -142.965 208.245 -142.635 ;
        RECT 207.915 -144.325 208.245 -143.995 ;
        RECT 207.915 -145.685 208.245 -145.355 ;
        RECT 207.915 -147.045 208.245 -146.715 ;
        RECT 207.915 -148.405 208.245 -148.075 ;
        RECT 207.915 -149.765 208.245 -149.435 ;
        RECT 207.915 -151.125 208.245 -150.795 ;
        RECT 207.915 -152.485 208.245 -152.155 ;
        RECT 207.915 -153.845 208.245 -153.515 ;
        RECT 207.915 -155.205 208.245 -154.875 ;
        RECT 207.915 -156.565 208.245 -156.235 ;
        RECT 207.915 -157.925 208.245 -157.595 ;
        RECT 207.915 -159.285 208.245 -158.955 ;
        RECT 207.915 -160.645 208.245 -160.315 ;
        RECT 207.915 -162.005 208.245 -161.675 ;
        RECT 207.915 -163.365 208.245 -163.035 ;
        RECT 207.915 -164.725 208.245 -164.395 ;
        RECT 207.915 -166.085 208.245 -165.755 ;
        RECT 207.915 -167.445 208.245 -167.115 ;
        RECT 207.915 -168.805 208.245 -168.475 ;
        RECT 207.915 -170.165 208.245 -169.835 ;
        RECT 207.915 -171.525 208.245 -171.195 ;
        RECT 207.915 -172.885 208.245 -172.555 ;
        RECT 207.915 -174.245 208.245 -173.915 ;
        RECT 207.915 -175.605 208.245 -175.275 ;
        RECT 207.915 -176.965 208.245 -176.635 ;
        RECT 207.915 -178.325 208.245 -177.995 ;
        RECT 207.915 -180.57 208.245 -179.44 ;
        RECT 207.92 -180.685 208.24 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 209.275 241.32 209.605 242.45 ;
        RECT 209.275 239.195 209.605 239.525 ;
        RECT 209.275 237.835 209.605 238.165 ;
        RECT 209.28 237.16 209.6 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 209.275 -1.525 209.605 -1.195 ;
        RECT 209.275 -2.885 209.605 -2.555 ;
        RECT 209.28 -3.56 209.6 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 209.275 -91.285 209.605 -90.955 ;
        RECT 209.275 -92.645 209.605 -92.315 ;
        RECT 209.275 -94.005 209.605 -93.675 ;
        RECT 209.275 -95.365 209.605 -95.035 ;
        RECT 209.275 -96.725 209.605 -96.395 ;
        RECT 209.275 -98.085 209.605 -97.755 ;
        RECT 209.275 -99.445 209.605 -99.115 ;
        RECT 209.275 -100.805 209.605 -100.475 ;
        RECT 209.275 -102.165 209.605 -101.835 ;
        RECT 209.275 -103.525 209.605 -103.195 ;
        RECT 209.275 -104.885 209.605 -104.555 ;
        RECT 209.275 -106.245 209.605 -105.915 ;
        RECT 209.275 -107.605 209.605 -107.275 ;
        RECT 209.275 -108.965 209.605 -108.635 ;
        RECT 209.275 -110.325 209.605 -109.995 ;
        RECT 209.275 -111.685 209.605 -111.355 ;
        RECT 209.275 -113.045 209.605 -112.715 ;
        RECT 209.275 -114.405 209.605 -114.075 ;
        RECT 209.275 -115.765 209.605 -115.435 ;
        RECT 209.275 -117.125 209.605 -116.795 ;
        RECT 209.275 -118.485 209.605 -118.155 ;
        RECT 209.275 -119.845 209.605 -119.515 ;
        RECT 209.275 -121.205 209.605 -120.875 ;
        RECT 209.275 -122.565 209.605 -122.235 ;
        RECT 209.275 -123.925 209.605 -123.595 ;
        RECT 209.275 -125.285 209.605 -124.955 ;
        RECT 209.275 -126.645 209.605 -126.315 ;
        RECT 209.275 -128.005 209.605 -127.675 ;
        RECT 209.275 -129.365 209.605 -129.035 ;
        RECT 209.275 -130.725 209.605 -130.395 ;
        RECT 209.275 -132.085 209.605 -131.755 ;
        RECT 209.275 -133.445 209.605 -133.115 ;
        RECT 209.275 -134.805 209.605 -134.475 ;
        RECT 209.275 -136.165 209.605 -135.835 ;
        RECT 209.275 -137.525 209.605 -137.195 ;
        RECT 209.275 -138.885 209.605 -138.555 ;
        RECT 209.275 -140.245 209.605 -139.915 ;
        RECT 209.275 -141.605 209.605 -141.275 ;
        RECT 209.275 -142.965 209.605 -142.635 ;
        RECT 209.275 -144.325 209.605 -143.995 ;
        RECT 209.275 -145.685 209.605 -145.355 ;
        RECT 209.275 -147.045 209.605 -146.715 ;
        RECT 209.275 -148.405 209.605 -148.075 ;
        RECT 209.275 -149.765 209.605 -149.435 ;
        RECT 209.275 -151.125 209.605 -150.795 ;
        RECT 209.275 -152.485 209.605 -152.155 ;
        RECT 209.275 -153.845 209.605 -153.515 ;
        RECT 209.275 -155.205 209.605 -154.875 ;
        RECT 209.275 -156.565 209.605 -156.235 ;
        RECT 209.275 -157.925 209.605 -157.595 ;
        RECT 209.275 -159.285 209.605 -158.955 ;
        RECT 209.275 -160.645 209.605 -160.315 ;
        RECT 209.275 -162.005 209.605 -161.675 ;
        RECT 209.275 -163.365 209.605 -163.035 ;
        RECT 209.275 -164.725 209.605 -164.395 ;
        RECT 209.275 -166.085 209.605 -165.755 ;
        RECT 209.275 -167.445 209.605 -167.115 ;
        RECT 209.275 -168.805 209.605 -168.475 ;
        RECT 209.275 -170.165 209.605 -169.835 ;
        RECT 209.275 -171.525 209.605 -171.195 ;
        RECT 209.275 -172.885 209.605 -172.555 ;
        RECT 209.275 -174.245 209.605 -173.915 ;
        RECT 209.275 -175.605 209.605 -175.275 ;
        RECT 209.275 -176.965 209.605 -176.635 ;
        RECT 209.275 -178.325 209.605 -177.995 ;
        RECT 209.275 -180.57 209.605 -179.44 ;
        RECT 209.28 -180.685 209.6 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 210.635 241.32 210.965 242.45 ;
        RECT 210.635 239.195 210.965 239.525 ;
        RECT 210.635 237.835 210.965 238.165 ;
        RECT 210.64 237.16 210.96 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 210.635 -95.365 210.965 -95.035 ;
        RECT 210.635 -96.725 210.965 -96.395 ;
        RECT 210.635 -98.085 210.965 -97.755 ;
        RECT 210.635 -99.445 210.965 -99.115 ;
        RECT 210.635 -100.805 210.965 -100.475 ;
        RECT 210.635 -102.165 210.965 -101.835 ;
        RECT 210.635 -103.525 210.965 -103.195 ;
        RECT 210.635 -104.885 210.965 -104.555 ;
        RECT 210.635 -106.245 210.965 -105.915 ;
        RECT 210.635 -107.605 210.965 -107.275 ;
        RECT 210.635 -108.965 210.965 -108.635 ;
        RECT 210.635 -110.325 210.965 -109.995 ;
        RECT 210.635 -111.685 210.965 -111.355 ;
        RECT 210.635 -113.045 210.965 -112.715 ;
        RECT 210.635 -114.405 210.965 -114.075 ;
        RECT 210.635 -115.765 210.965 -115.435 ;
        RECT 210.635 -117.125 210.965 -116.795 ;
        RECT 210.635 -118.485 210.965 -118.155 ;
        RECT 210.635 -119.845 210.965 -119.515 ;
        RECT 210.635 -121.205 210.965 -120.875 ;
        RECT 210.635 -122.565 210.965 -122.235 ;
        RECT 210.635 -123.925 210.965 -123.595 ;
        RECT 210.635 -125.285 210.965 -124.955 ;
        RECT 210.635 -126.645 210.965 -126.315 ;
        RECT 210.635 -128.005 210.965 -127.675 ;
        RECT 210.635 -129.365 210.965 -129.035 ;
        RECT 210.635 -130.725 210.965 -130.395 ;
        RECT 210.635 -132.085 210.965 -131.755 ;
        RECT 210.635 -133.445 210.965 -133.115 ;
        RECT 210.635 -134.805 210.965 -134.475 ;
        RECT 210.635 -136.165 210.965 -135.835 ;
        RECT 210.635 -137.525 210.965 -137.195 ;
        RECT 210.635 -138.885 210.965 -138.555 ;
        RECT 210.635 -140.245 210.965 -139.915 ;
        RECT 210.635 -141.605 210.965 -141.275 ;
        RECT 210.635 -142.965 210.965 -142.635 ;
        RECT 210.635 -144.325 210.965 -143.995 ;
        RECT 210.635 -145.685 210.965 -145.355 ;
        RECT 210.635 -147.045 210.965 -146.715 ;
        RECT 210.635 -148.405 210.965 -148.075 ;
        RECT 210.635 -149.765 210.965 -149.435 ;
        RECT 210.635 -151.125 210.965 -150.795 ;
        RECT 210.635 -152.485 210.965 -152.155 ;
        RECT 210.635 -153.845 210.965 -153.515 ;
        RECT 210.635 -155.205 210.965 -154.875 ;
        RECT 210.635 -156.565 210.965 -156.235 ;
        RECT 210.635 -157.925 210.965 -157.595 ;
        RECT 210.635 -159.285 210.965 -158.955 ;
        RECT 210.635 -160.645 210.965 -160.315 ;
        RECT 210.635 -162.005 210.965 -161.675 ;
        RECT 210.635 -163.365 210.965 -163.035 ;
        RECT 210.635 -164.725 210.965 -164.395 ;
        RECT 210.635 -166.085 210.965 -165.755 ;
        RECT 210.635 -167.445 210.965 -167.115 ;
        RECT 210.635 -168.805 210.965 -168.475 ;
        RECT 210.635 -170.165 210.965 -169.835 ;
        RECT 210.635 -171.525 210.965 -171.195 ;
        RECT 210.635 -172.885 210.965 -172.555 ;
        RECT 210.635 -174.245 210.965 -173.915 ;
        RECT 210.635 -175.605 210.965 -175.275 ;
        RECT 210.635 -176.965 210.965 -176.635 ;
        RECT 210.635 -178.325 210.965 -177.995 ;
        RECT 210.635 -180.57 210.965 -179.44 ;
        RECT 210.64 -180.685 210.96 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 210.71 -94.075 211.04 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 211.995 241.32 212.325 242.45 ;
        RECT 211.995 239.195 212.325 239.525 ;
        RECT 211.995 237.835 212.325 238.165 ;
        RECT 212 237.16 212.32 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 211.995 -1.525 212.325 -1.195 ;
        RECT 211.995 -2.885 212.325 -2.555 ;
        RECT 212 -3.56 212.32 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 213.355 241.32 213.685 242.45 ;
        RECT 213.355 239.195 213.685 239.525 ;
        RECT 213.355 237.835 213.685 238.165 ;
        RECT 213.36 237.16 213.68 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 213.355 -1.525 213.685 -1.195 ;
        RECT 213.355 -2.885 213.685 -2.555 ;
        RECT 213.36 -3.56 213.68 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 214.715 241.32 215.045 242.45 ;
        RECT 214.715 239.195 215.045 239.525 ;
        RECT 214.715 237.835 215.045 238.165 ;
        RECT 214.72 237.16 215.04 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 214.715 -1.525 215.045 -1.195 ;
        RECT 214.715 -2.885 215.045 -2.555 ;
        RECT 214.72 -3.56 215.04 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 214.715 -91.285 215.045 -90.955 ;
        RECT 214.715 -92.645 215.045 -92.315 ;
        RECT 214.715 -94.005 215.045 -93.675 ;
        RECT 214.715 -95.365 215.045 -95.035 ;
        RECT 214.715 -96.725 215.045 -96.395 ;
        RECT 214.715 -98.085 215.045 -97.755 ;
        RECT 214.715 -99.445 215.045 -99.115 ;
        RECT 214.715 -100.805 215.045 -100.475 ;
        RECT 214.715 -102.165 215.045 -101.835 ;
        RECT 214.715 -103.525 215.045 -103.195 ;
        RECT 214.715 -104.885 215.045 -104.555 ;
        RECT 214.715 -106.245 215.045 -105.915 ;
        RECT 214.715 -107.605 215.045 -107.275 ;
        RECT 214.715 -108.965 215.045 -108.635 ;
        RECT 214.715 -110.325 215.045 -109.995 ;
        RECT 214.715 -111.685 215.045 -111.355 ;
        RECT 214.715 -113.045 215.045 -112.715 ;
        RECT 214.715 -114.405 215.045 -114.075 ;
        RECT 214.715 -115.765 215.045 -115.435 ;
        RECT 214.715 -117.125 215.045 -116.795 ;
        RECT 214.715 -118.485 215.045 -118.155 ;
        RECT 214.715 -119.845 215.045 -119.515 ;
        RECT 214.715 -121.205 215.045 -120.875 ;
        RECT 214.715 -122.565 215.045 -122.235 ;
        RECT 214.715 -123.925 215.045 -123.595 ;
        RECT 214.715 -125.285 215.045 -124.955 ;
        RECT 214.715 -126.645 215.045 -126.315 ;
        RECT 214.715 -128.005 215.045 -127.675 ;
        RECT 214.715 -129.365 215.045 -129.035 ;
        RECT 214.715 -130.725 215.045 -130.395 ;
        RECT 214.715 -132.085 215.045 -131.755 ;
        RECT 214.715 -133.445 215.045 -133.115 ;
        RECT 214.715 -134.805 215.045 -134.475 ;
        RECT 214.715 -136.165 215.045 -135.835 ;
        RECT 214.715 -137.525 215.045 -137.195 ;
        RECT 214.715 -138.885 215.045 -138.555 ;
        RECT 214.715 -140.245 215.045 -139.915 ;
        RECT 214.715 -141.605 215.045 -141.275 ;
        RECT 214.715 -142.965 215.045 -142.635 ;
        RECT 214.715 -144.325 215.045 -143.995 ;
        RECT 214.715 -145.685 215.045 -145.355 ;
        RECT 214.715 -147.045 215.045 -146.715 ;
        RECT 214.715 -148.405 215.045 -148.075 ;
        RECT 214.715 -149.765 215.045 -149.435 ;
        RECT 214.715 -151.125 215.045 -150.795 ;
        RECT 214.715 -152.485 215.045 -152.155 ;
        RECT 214.715 -153.845 215.045 -153.515 ;
        RECT 214.715 -155.205 215.045 -154.875 ;
        RECT 214.715 -156.565 215.045 -156.235 ;
        RECT 214.715 -157.925 215.045 -157.595 ;
        RECT 214.715 -159.285 215.045 -158.955 ;
        RECT 214.715 -160.645 215.045 -160.315 ;
        RECT 214.715 -162.005 215.045 -161.675 ;
        RECT 214.715 -163.365 215.045 -163.035 ;
        RECT 214.715 -164.725 215.045 -164.395 ;
        RECT 214.715 -166.085 215.045 -165.755 ;
        RECT 214.715 -167.445 215.045 -167.115 ;
        RECT 214.715 -168.805 215.045 -168.475 ;
        RECT 214.715 -170.165 215.045 -169.835 ;
        RECT 214.715 -171.525 215.045 -171.195 ;
        RECT 214.715 -172.885 215.045 -172.555 ;
        RECT 214.715 -174.245 215.045 -173.915 ;
        RECT 214.715 -175.605 215.045 -175.275 ;
        RECT 214.715 -176.965 215.045 -176.635 ;
        RECT 214.715 -178.325 215.045 -177.995 ;
        RECT 214.715 -180.57 215.045 -179.44 ;
        RECT 214.72 -180.685 215.04 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 216.075 241.32 216.405 242.45 ;
        RECT 216.075 239.195 216.405 239.525 ;
        RECT 216.075 237.835 216.405 238.165 ;
        RECT 216.08 237.16 216.4 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 216.075 -95.365 216.405 -95.035 ;
        RECT 216.075 -96.725 216.405 -96.395 ;
        RECT 216.075 -98.085 216.405 -97.755 ;
        RECT 216.075 -99.445 216.405 -99.115 ;
        RECT 216.075 -100.805 216.405 -100.475 ;
        RECT 216.075 -102.165 216.405 -101.835 ;
        RECT 216.075 -103.525 216.405 -103.195 ;
        RECT 216.075 -104.885 216.405 -104.555 ;
        RECT 216.075 -106.245 216.405 -105.915 ;
        RECT 216.075 -107.605 216.405 -107.275 ;
        RECT 216.075 -108.965 216.405 -108.635 ;
        RECT 216.075 -110.325 216.405 -109.995 ;
        RECT 216.075 -111.685 216.405 -111.355 ;
        RECT 216.075 -113.045 216.405 -112.715 ;
        RECT 216.075 -114.405 216.405 -114.075 ;
        RECT 216.075 -115.765 216.405 -115.435 ;
        RECT 216.075 -117.125 216.405 -116.795 ;
        RECT 216.075 -118.485 216.405 -118.155 ;
        RECT 216.075 -119.845 216.405 -119.515 ;
        RECT 216.075 -121.205 216.405 -120.875 ;
        RECT 216.075 -122.565 216.405 -122.235 ;
        RECT 216.075 -123.925 216.405 -123.595 ;
        RECT 216.075 -125.285 216.405 -124.955 ;
        RECT 216.075 -126.645 216.405 -126.315 ;
        RECT 216.075 -128.005 216.405 -127.675 ;
        RECT 216.075 -129.365 216.405 -129.035 ;
        RECT 216.075 -130.725 216.405 -130.395 ;
        RECT 216.075 -132.085 216.405 -131.755 ;
        RECT 216.075 -133.445 216.405 -133.115 ;
        RECT 216.075 -134.805 216.405 -134.475 ;
        RECT 216.075 -136.165 216.405 -135.835 ;
        RECT 216.075 -137.525 216.405 -137.195 ;
        RECT 216.075 -138.885 216.405 -138.555 ;
        RECT 216.075 -140.245 216.405 -139.915 ;
        RECT 216.075 -141.605 216.405 -141.275 ;
        RECT 216.075 -142.965 216.405 -142.635 ;
        RECT 216.075 -144.325 216.405 -143.995 ;
        RECT 216.075 -145.685 216.405 -145.355 ;
        RECT 216.075 -147.045 216.405 -146.715 ;
        RECT 216.075 -148.405 216.405 -148.075 ;
        RECT 216.075 -149.765 216.405 -149.435 ;
        RECT 216.075 -151.125 216.405 -150.795 ;
        RECT 216.075 -152.485 216.405 -152.155 ;
        RECT 216.075 -153.845 216.405 -153.515 ;
        RECT 216.075 -155.205 216.405 -154.875 ;
        RECT 216.075 -156.565 216.405 -156.235 ;
        RECT 216.075 -157.925 216.405 -157.595 ;
        RECT 216.075 -159.285 216.405 -158.955 ;
        RECT 216.075 -160.645 216.405 -160.315 ;
        RECT 216.075 -162.005 216.405 -161.675 ;
        RECT 216.075 -163.365 216.405 -163.035 ;
        RECT 216.075 -164.725 216.405 -164.395 ;
        RECT 216.075 -166.085 216.405 -165.755 ;
        RECT 216.075 -167.445 216.405 -167.115 ;
        RECT 216.075 -168.805 216.405 -168.475 ;
        RECT 216.075 -170.165 216.405 -169.835 ;
        RECT 216.075 -171.525 216.405 -171.195 ;
        RECT 216.075 -172.885 216.405 -172.555 ;
        RECT 216.075 -174.245 216.405 -173.915 ;
        RECT 216.075 -175.605 216.405 -175.275 ;
        RECT 216.075 -176.965 216.405 -176.635 ;
        RECT 216.075 -178.325 216.405 -177.995 ;
        RECT 216.075 -180.57 216.405 -179.44 ;
        RECT 216.08 -180.685 216.4 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 216.81 -94.075 217.14 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 217.435 241.32 217.765 242.45 ;
        RECT 217.435 239.195 217.765 239.525 ;
        RECT 217.435 237.835 217.765 238.165 ;
        RECT 217.44 237.16 217.76 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 218.795 241.32 219.125 242.45 ;
        RECT 218.795 239.195 219.125 239.525 ;
        RECT 218.795 237.835 219.125 238.165 ;
        RECT 218.8 237.16 219.12 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 218.795 -1.525 219.125 -1.195 ;
        RECT 218.795 -2.885 219.125 -2.555 ;
        RECT 218.8 -3.56 219.12 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 220.155 241.32 220.485 242.45 ;
        RECT 220.155 239.195 220.485 239.525 ;
        RECT 220.155 237.835 220.485 238.165 ;
        RECT 220.16 237.16 220.48 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 220.155 -1.525 220.485 -1.195 ;
        RECT 220.155 -2.885 220.485 -2.555 ;
        RECT 220.16 -3.56 220.48 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 220.155 -91.285 220.485 -90.955 ;
        RECT 220.155 -92.645 220.485 -92.315 ;
        RECT 220.155 -94.005 220.485 -93.675 ;
        RECT 220.155 -95.365 220.485 -95.035 ;
        RECT 220.155 -96.725 220.485 -96.395 ;
        RECT 220.155 -98.085 220.485 -97.755 ;
        RECT 220.155 -99.445 220.485 -99.115 ;
        RECT 220.155 -100.805 220.485 -100.475 ;
        RECT 220.155 -102.165 220.485 -101.835 ;
        RECT 220.155 -103.525 220.485 -103.195 ;
        RECT 220.155 -104.885 220.485 -104.555 ;
        RECT 220.155 -106.245 220.485 -105.915 ;
        RECT 220.155 -107.605 220.485 -107.275 ;
        RECT 220.155 -108.965 220.485 -108.635 ;
        RECT 220.155 -110.325 220.485 -109.995 ;
        RECT 220.155 -111.685 220.485 -111.355 ;
        RECT 220.155 -113.045 220.485 -112.715 ;
        RECT 220.155 -114.405 220.485 -114.075 ;
        RECT 220.155 -115.765 220.485 -115.435 ;
        RECT 220.155 -117.125 220.485 -116.795 ;
        RECT 220.155 -118.485 220.485 -118.155 ;
        RECT 220.155 -119.845 220.485 -119.515 ;
        RECT 220.155 -121.205 220.485 -120.875 ;
        RECT 220.155 -122.565 220.485 -122.235 ;
        RECT 220.155 -123.925 220.485 -123.595 ;
        RECT 220.155 -125.285 220.485 -124.955 ;
        RECT 220.155 -126.645 220.485 -126.315 ;
        RECT 220.155 -128.005 220.485 -127.675 ;
        RECT 220.155 -129.365 220.485 -129.035 ;
        RECT 220.155 -130.725 220.485 -130.395 ;
        RECT 220.155 -132.085 220.485 -131.755 ;
        RECT 220.155 -133.445 220.485 -133.115 ;
        RECT 220.155 -134.805 220.485 -134.475 ;
        RECT 220.155 -136.165 220.485 -135.835 ;
        RECT 220.155 -137.525 220.485 -137.195 ;
        RECT 220.155 -138.885 220.485 -138.555 ;
        RECT 220.155 -140.245 220.485 -139.915 ;
        RECT 220.155 -141.605 220.485 -141.275 ;
        RECT 220.155 -142.965 220.485 -142.635 ;
        RECT 220.155 -144.325 220.485 -143.995 ;
        RECT 220.155 -145.685 220.485 -145.355 ;
        RECT 220.155 -147.045 220.485 -146.715 ;
        RECT 220.155 -148.405 220.485 -148.075 ;
        RECT 220.155 -149.765 220.485 -149.435 ;
        RECT 220.155 -151.125 220.485 -150.795 ;
        RECT 220.155 -152.485 220.485 -152.155 ;
        RECT 220.155 -153.845 220.485 -153.515 ;
        RECT 220.155 -155.205 220.485 -154.875 ;
        RECT 220.155 -156.565 220.485 -156.235 ;
        RECT 220.155 -157.925 220.485 -157.595 ;
        RECT 220.155 -159.285 220.485 -158.955 ;
        RECT 220.155 -160.645 220.485 -160.315 ;
        RECT 220.155 -162.005 220.485 -161.675 ;
        RECT 220.155 -163.365 220.485 -163.035 ;
        RECT 220.155 -164.725 220.485 -164.395 ;
        RECT 220.155 -166.085 220.485 -165.755 ;
        RECT 220.155 -167.445 220.485 -167.115 ;
        RECT 220.155 -168.805 220.485 -168.475 ;
        RECT 220.155 -170.165 220.485 -169.835 ;
        RECT 220.155 -171.525 220.485 -171.195 ;
        RECT 220.155 -172.885 220.485 -172.555 ;
        RECT 220.155 -174.245 220.485 -173.915 ;
        RECT 220.155 -175.605 220.485 -175.275 ;
        RECT 220.155 -176.965 220.485 -176.635 ;
        RECT 220.155 -178.325 220.485 -177.995 ;
        RECT 220.155 -180.57 220.485 -179.44 ;
        RECT 220.16 -180.685 220.48 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 221.515 241.32 221.845 242.45 ;
        RECT 221.515 239.195 221.845 239.525 ;
        RECT 221.515 237.835 221.845 238.165 ;
        RECT 221.52 237.16 221.84 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 221.515 -1.525 221.845 -1.195 ;
        RECT 221.515 -2.885 221.845 -2.555 ;
        RECT 221.52 -3.56 221.84 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 221.515 -91.285 221.845 -90.955 ;
        RECT 221.515 -92.645 221.845 -92.315 ;
        RECT 221.515 -94.005 221.845 -93.675 ;
        RECT 221.515 -95.365 221.845 -95.035 ;
        RECT 221.515 -96.725 221.845 -96.395 ;
        RECT 221.515 -98.085 221.845 -97.755 ;
        RECT 221.515 -99.445 221.845 -99.115 ;
        RECT 221.515 -100.805 221.845 -100.475 ;
        RECT 221.515 -102.165 221.845 -101.835 ;
        RECT 221.515 -103.525 221.845 -103.195 ;
        RECT 221.515 -104.885 221.845 -104.555 ;
        RECT 221.515 -106.245 221.845 -105.915 ;
        RECT 221.515 -107.605 221.845 -107.275 ;
        RECT 221.515 -108.965 221.845 -108.635 ;
        RECT 221.515 -110.325 221.845 -109.995 ;
        RECT 221.515 -111.685 221.845 -111.355 ;
        RECT 221.515 -113.045 221.845 -112.715 ;
        RECT 221.515 -114.405 221.845 -114.075 ;
        RECT 221.515 -115.765 221.845 -115.435 ;
        RECT 221.515 -117.125 221.845 -116.795 ;
        RECT 221.515 -118.485 221.845 -118.155 ;
        RECT 221.515 -119.845 221.845 -119.515 ;
        RECT 221.515 -121.205 221.845 -120.875 ;
        RECT 221.515 -122.565 221.845 -122.235 ;
        RECT 221.515 -123.925 221.845 -123.595 ;
        RECT 221.515 -125.285 221.845 -124.955 ;
        RECT 221.515 -126.645 221.845 -126.315 ;
        RECT 221.515 -128.005 221.845 -127.675 ;
        RECT 221.515 -129.365 221.845 -129.035 ;
        RECT 221.515 -130.725 221.845 -130.395 ;
        RECT 221.515 -132.085 221.845 -131.755 ;
        RECT 221.515 -133.445 221.845 -133.115 ;
        RECT 221.515 -134.805 221.845 -134.475 ;
        RECT 221.515 -136.165 221.845 -135.835 ;
        RECT 221.515 -137.525 221.845 -137.195 ;
        RECT 221.515 -138.885 221.845 -138.555 ;
        RECT 221.515 -140.245 221.845 -139.915 ;
        RECT 221.515 -141.605 221.845 -141.275 ;
        RECT 221.515 -142.965 221.845 -142.635 ;
        RECT 221.515 -144.325 221.845 -143.995 ;
        RECT 221.515 -145.685 221.845 -145.355 ;
        RECT 221.515 -147.045 221.845 -146.715 ;
        RECT 221.515 -148.405 221.845 -148.075 ;
        RECT 221.515 -149.765 221.845 -149.435 ;
        RECT 221.515 -151.125 221.845 -150.795 ;
        RECT 221.515 -152.485 221.845 -152.155 ;
        RECT 221.515 -153.845 221.845 -153.515 ;
        RECT 221.515 -155.205 221.845 -154.875 ;
        RECT 221.515 -156.565 221.845 -156.235 ;
        RECT 221.515 -157.925 221.845 -157.595 ;
        RECT 221.515 -159.285 221.845 -158.955 ;
        RECT 221.515 -160.645 221.845 -160.315 ;
        RECT 221.515 -162.005 221.845 -161.675 ;
        RECT 221.515 -163.365 221.845 -163.035 ;
        RECT 221.515 -164.725 221.845 -164.395 ;
        RECT 221.515 -166.085 221.845 -165.755 ;
        RECT 221.515 -167.445 221.845 -167.115 ;
        RECT 221.515 -168.805 221.845 -168.475 ;
        RECT 221.515 -170.165 221.845 -169.835 ;
        RECT 221.515 -171.525 221.845 -171.195 ;
        RECT 221.515 -172.885 221.845 -172.555 ;
        RECT 221.515 -174.245 221.845 -173.915 ;
        RECT 221.515 -175.605 221.845 -175.275 ;
        RECT 221.515 -176.965 221.845 -176.635 ;
        RECT 221.515 -178.325 221.845 -177.995 ;
        RECT 221.515 -180.57 221.845 -179.44 ;
        RECT 221.52 -180.685 221.84 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 222.875 241.32 223.205 242.45 ;
        RECT 222.875 239.195 223.205 239.525 ;
        RECT 222.875 237.835 223.205 238.165 ;
        RECT 222.88 237.16 223.2 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 222.875 -95.365 223.205 -95.035 ;
        RECT 222.875 -96.725 223.205 -96.395 ;
        RECT 222.875 -98.085 223.205 -97.755 ;
        RECT 222.875 -99.445 223.205 -99.115 ;
        RECT 222.875 -100.805 223.205 -100.475 ;
        RECT 222.875 -102.165 223.205 -101.835 ;
        RECT 222.875 -103.525 223.205 -103.195 ;
        RECT 222.875 -104.885 223.205 -104.555 ;
        RECT 222.875 -106.245 223.205 -105.915 ;
        RECT 222.875 -107.605 223.205 -107.275 ;
        RECT 222.875 -108.965 223.205 -108.635 ;
        RECT 222.875 -110.325 223.205 -109.995 ;
        RECT 222.875 -111.685 223.205 -111.355 ;
        RECT 222.875 -113.045 223.205 -112.715 ;
        RECT 222.875 -114.405 223.205 -114.075 ;
        RECT 222.875 -115.765 223.205 -115.435 ;
        RECT 222.875 -117.125 223.205 -116.795 ;
        RECT 222.875 -118.485 223.205 -118.155 ;
        RECT 222.875 -119.845 223.205 -119.515 ;
        RECT 222.875 -121.205 223.205 -120.875 ;
        RECT 222.875 -122.565 223.205 -122.235 ;
        RECT 222.875 -123.925 223.205 -123.595 ;
        RECT 222.875 -125.285 223.205 -124.955 ;
        RECT 222.875 -126.645 223.205 -126.315 ;
        RECT 222.875 -128.005 223.205 -127.675 ;
        RECT 222.875 -129.365 223.205 -129.035 ;
        RECT 222.875 -130.725 223.205 -130.395 ;
        RECT 222.875 -132.085 223.205 -131.755 ;
        RECT 222.875 -133.445 223.205 -133.115 ;
        RECT 222.875 -134.805 223.205 -134.475 ;
        RECT 222.875 -136.165 223.205 -135.835 ;
        RECT 222.875 -137.525 223.205 -137.195 ;
        RECT 222.875 -138.885 223.205 -138.555 ;
        RECT 222.875 -140.245 223.205 -139.915 ;
        RECT 222.875 -141.605 223.205 -141.275 ;
        RECT 222.875 -142.965 223.205 -142.635 ;
        RECT 222.875 -144.325 223.205 -143.995 ;
        RECT 222.875 -145.685 223.205 -145.355 ;
        RECT 222.875 -147.045 223.205 -146.715 ;
        RECT 222.875 -148.405 223.205 -148.075 ;
        RECT 222.875 -149.765 223.205 -149.435 ;
        RECT 222.875 -151.125 223.205 -150.795 ;
        RECT 222.875 -152.485 223.205 -152.155 ;
        RECT 222.875 -153.845 223.205 -153.515 ;
        RECT 222.875 -155.205 223.205 -154.875 ;
        RECT 222.875 -156.565 223.205 -156.235 ;
        RECT 222.875 -157.925 223.205 -157.595 ;
        RECT 222.875 -159.285 223.205 -158.955 ;
        RECT 222.875 -160.645 223.205 -160.315 ;
        RECT 222.875 -162.005 223.205 -161.675 ;
        RECT 222.875 -163.365 223.205 -163.035 ;
        RECT 222.875 -164.725 223.205 -164.395 ;
        RECT 222.875 -166.085 223.205 -165.755 ;
        RECT 222.875 -167.445 223.205 -167.115 ;
        RECT 222.875 -168.805 223.205 -168.475 ;
        RECT 222.875 -170.165 223.205 -169.835 ;
        RECT 222.875 -171.525 223.205 -171.195 ;
        RECT 222.875 -172.885 223.205 -172.555 ;
        RECT 222.875 -174.245 223.205 -173.915 ;
        RECT 222.875 -175.605 223.205 -175.275 ;
        RECT 222.875 -176.965 223.205 -176.635 ;
        RECT 222.875 -178.325 223.205 -177.995 ;
        RECT 222.875 -180.57 223.205 -179.44 ;
        RECT 222.88 -180.685 223.2 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 222.91 -94.075 223.24 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 224.235 241.32 224.565 242.45 ;
        RECT 224.235 239.195 224.565 239.525 ;
        RECT 224.235 237.835 224.565 238.165 ;
        RECT 224.24 237.16 224.56 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 224.235 -1.525 224.565 -1.195 ;
        RECT 224.235 -2.885 224.565 -2.555 ;
        RECT 224.24 -3.56 224.56 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 225.595 241.32 225.925 242.45 ;
        RECT 225.595 239.195 225.925 239.525 ;
        RECT 225.595 237.835 225.925 238.165 ;
        RECT 225.6 237.16 225.92 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 225.595 -1.525 225.925 -1.195 ;
        RECT 225.595 -2.885 225.925 -2.555 ;
        RECT 225.6 -3.56 225.92 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 226.955 241.32 227.285 242.45 ;
        RECT 226.955 239.195 227.285 239.525 ;
        RECT 226.955 237.835 227.285 238.165 ;
        RECT 226.96 237.16 227.28 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 226.955 -1.525 227.285 -1.195 ;
        RECT 226.955 -2.885 227.285 -2.555 ;
        RECT 226.96 -3.56 227.28 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 226.955 -91.285 227.285 -90.955 ;
        RECT 226.955 -92.645 227.285 -92.315 ;
        RECT 226.955 -94.005 227.285 -93.675 ;
        RECT 226.955 -95.365 227.285 -95.035 ;
        RECT 226.955 -96.725 227.285 -96.395 ;
        RECT 226.955 -98.085 227.285 -97.755 ;
        RECT 226.955 -99.445 227.285 -99.115 ;
        RECT 226.955 -100.805 227.285 -100.475 ;
        RECT 226.955 -102.165 227.285 -101.835 ;
        RECT 226.955 -103.525 227.285 -103.195 ;
        RECT 226.955 -104.885 227.285 -104.555 ;
        RECT 226.955 -106.245 227.285 -105.915 ;
        RECT 226.955 -107.605 227.285 -107.275 ;
        RECT 226.955 -108.965 227.285 -108.635 ;
        RECT 226.955 -110.325 227.285 -109.995 ;
        RECT 226.955 -111.685 227.285 -111.355 ;
        RECT 226.955 -113.045 227.285 -112.715 ;
        RECT 226.955 -114.405 227.285 -114.075 ;
        RECT 226.955 -115.765 227.285 -115.435 ;
        RECT 226.955 -117.125 227.285 -116.795 ;
        RECT 226.955 -118.485 227.285 -118.155 ;
        RECT 226.955 -119.845 227.285 -119.515 ;
        RECT 226.955 -121.205 227.285 -120.875 ;
        RECT 226.955 -122.565 227.285 -122.235 ;
        RECT 226.955 -123.925 227.285 -123.595 ;
        RECT 226.955 -125.285 227.285 -124.955 ;
        RECT 226.955 -126.645 227.285 -126.315 ;
        RECT 226.955 -128.005 227.285 -127.675 ;
        RECT 226.955 -129.365 227.285 -129.035 ;
        RECT 226.955 -130.725 227.285 -130.395 ;
        RECT 226.955 -132.085 227.285 -131.755 ;
        RECT 226.955 -133.445 227.285 -133.115 ;
        RECT 226.955 -134.805 227.285 -134.475 ;
        RECT 226.955 -136.165 227.285 -135.835 ;
        RECT 226.955 -137.525 227.285 -137.195 ;
        RECT 226.955 -138.885 227.285 -138.555 ;
        RECT 226.955 -140.245 227.285 -139.915 ;
        RECT 226.955 -141.605 227.285 -141.275 ;
        RECT 226.955 -142.965 227.285 -142.635 ;
        RECT 226.955 -144.325 227.285 -143.995 ;
        RECT 226.955 -145.685 227.285 -145.355 ;
        RECT 226.955 -147.045 227.285 -146.715 ;
        RECT 226.955 -148.405 227.285 -148.075 ;
        RECT 226.955 -149.765 227.285 -149.435 ;
        RECT 226.955 -151.125 227.285 -150.795 ;
        RECT 226.955 -152.485 227.285 -152.155 ;
        RECT 226.955 -153.845 227.285 -153.515 ;
        RECT 226.955 -155.205 227.285 -154.875 ;
        RECT 226.955 -156.565 227.285 -156.235 ;
        RECT 226.955 -157.925 227.285 -157.595 ;
        RECT 226.955 -159.285 227.285 -158.955 ;
        RECT 226.955 -160.645 227.285 -160.315 ;
        RECT 226.955 -162.005 227.285 -161.675 ;
        RECT 226.955 -163.365 227.285 -163.035 ;
        RECT 226.955 -164.725 227.285 -164.395 ;
        RECT 226.955 -166.085 227.285 -165.755 ;
        RECT 226.955 -167.445 227.285 -167.115 ;
        RECT 226.955 -168.805 227.285 -168.475 ;
        RECT 226.955 -170.165 227.285 -169.835 ;
        RECT 226.955 -171.525 227.285 -171.195 ;
        RECT 226.955 -172.885 227.285 -172.555 ;
        RECT 226.955 -174.245 227.285 -173.915 ;
        RECT 226.955 -175.605 227.285 -175.275 ;
        RECT 226.955 -176.965 227.285 -176.635 ;
        RECT 226.955 -178.325 227.285 -177.995 ;
        RECT 226.955 -180.57 227.285 -179.44 ;
        RECT 226.96 -180.685 227.28 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 228.315 241.32 228.645 242.45 ;
        RECT 228.315 239.195 228.645 239.525 ;
        RECT 228.315 237.835 228.645 238.165 ;
        RECT 228.32 237.16 228.64 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 228.315 -95.365 228.645 -95.035 ;
        RECT 228.315 -96.725 228.645 -96.395 ;
        RECT 228.315 -98.085 228.645 -97.755 ;
        RECT 228.315 -99.445 228.645 -99.115 ;
        RECT 228.315 -100.805 228.645 -100.475 ;
        RECT 228.315 -102.165 228.645 -101.835 ;
        RECT 228.315 -103.525 228.645 -103.195 ;
        RECT 228.315 -104.885 228.645 -104.555 ;
        RECT 228.315 -106.245 228.645 -105.915 ;
        RECT 228.315 -107.605 228.645 -107.275 ;
        RECT 228.315 -108.965 228.645 -108.635 ;
        RECT 228.315 -110.325 228.645 -109.995 ;
        RECT 228.315 -111.685 228.645 -111.355 ;
        RECT 228.315 -113.045 228.645 -112.715 ;
        RECT 228.315 -114.405 228.645 -114.075 ;
        RECT 228.315 -115.765 228.645 -115.435 ;
        RECT 228.315 -117.125 228.645 -116.795 ;
        RECT 228.315 -118.485 228.645 -118.155 ;
        RECT 228.315 -119.845 228.645 -119.515 ;
        RECT 228.315 -121.205 228.645 -120.875 ;
        RECT 228.315 -122.565 228.645 -122.235 ;
        RECT 228.315 -123.925 228.645 -123.595 ;
        RECT 228.315 -125.285 228.645 -124.955 ;
        RECT 228.315 -126.645 228.645 -126.315 ;
        RECT 228.315 -128.005 228.645 -127.675 ;
        RECT 228.315 -129.365 228.645 -129.035 ;
        RECT 228.315 -130.725 228.645 -130.395 ;
        RECT 228.315 -132.085 228.645 -131.755 ;
        RECT 228.315 -133.445 228.645 -133.115 ;
        RECT 228.315 -134.805 228.645 -134.475 ;
        RECT 228.315 -136.165 228.645 -135.835 ;
        RECT 228.315 -137.525 228.645 -137.195 ;
        RECT 228.315 -138.885 228.645 -138.555 ;
        RECT 228.315 -140.245 228.645 -139.915 ;
        RECT 228.315 -141.605 228.645 -141.275 ;
        RECT 228.315 -142.965 228.645 -142.635 ;
        RECT 228.315 -144.325 228.645 -143.995 ;
        RECT 228.315 -145.685 228.645 -145.355 ;
        RECT 228.315 -147.045 228.645 -146.715 ;
        RECT 228.315 -148.405 228.645 -148.075 ;
        RECT 228.315 -149.765 228.645 -149.435 ;
        RECT 228.315 -151.125 228.645 -150.795 ;
        RECT 228.315 -152.485 228.645 -152.155 ;
        RECT 228.315 -153.845 228.645 -153.515 ;
        RECT 228.315 -155.205 228.645 -154.875 ;
        RECT 228.315 -156.565 228.645 -156.235 ;
        RECT 228.315 -157.925 228.645 -157.595 ;
        RECT 228.315 -159.285 228.645 -158.955 ;
        RECT 228.315 -160.645 228.645 -160.315 ;
        RECT 228.315 -162.005 228.645 -161.675 ;
        RECT 228.315 -163.365 228.645 -163.035 ;
        RECT 228.315 -164.725 228.645 -164.395 ;
        RECT 228.315 -166.085 228.645 -165.755 ;
        RECT 228.315 -167.445 228.645 -167.115 ;
        RECT 228.315 -168.805 228.645 -168.475 ;
        RECT 228.315 -170.165 228.645 -169.835 ;
        RECT 228.315 -171.525 228.645 -171.195 ;
        RECT 228.315 -172.885 228.645 -172.555 ;
        RECT 228.315 -174.245 228.645 -173.915 ;
        RECT 228.315 -175.605 228.645 -175.275 ;
        RECT 228.315 -176.965 228.645 -176.635 ;
        RECT 228.315 -178.325 228.645 -177.995 ;
        RECT 228.315 -180.57 228.645 -179.44 ;
        RECT 228.32 -180.685 228.64 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 229.01 -94.075 229.34 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 229.675 241.32 230.005 242.45 ;
        RECT 229.675 239.195 230.005 239.525 ;
        RECT 229.675 237.835 230.005 238.165 ;
        RECT 229.68 237.16 230 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 231.035 241.32 231.365 242.45 ;
        RECT 231.035 239.195 231.365 239.525 ;
        RECT 231.035 237.835 231.365 238.165 ;
        RECT 231.04 237.16 231.36 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 231.035 -1.525 231.365 -1.195 ;
        RECT 231.035 -2.885 231.365 -2.555 ;
        RECT 231.04 -3.56 231.36 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 232.395 241.32 232.725 242.45 ;
        RECT 232.395 239.195 232.725 239.525 ;
        RECT 232.395 237.835 232.725 238.165 ;
        RECT 232.4 237.16 232.72 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 232.395 -1.525 232.725 -1.195 ;
        RECT 232.395 -2.885 232.725 -2.555 ;
        RECT 232.4 -3.56 232.72 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 232.395 -91.285 232.725 -90.955 ;
        RECT 232.395 -92.645 232.725 -92.315 ;
        RECT 232.395 -94.005 232.725 -93.675 ;
        RECT 232.395 -95.365 232.725 -95.035 ;
        RECT 232.395 -96.725 232.725 -96.395 ;
        RECT 232.395 -98.085 232.725 -97.755 ;
        RECT 232.395 -99.445 232.725 -99.115 ;
        RECT 232.395 -100.805 232.725 -100.475 ;
        RECT 232.395 -102.165 232.725 -101.835 ;
        RECT 232.395 -103.525 232.725 -103.195 ;
        RECT 232.395 -104.885 232.725 -104.555 ;
        RECT 232.395 -106.245 232.725 -105.915 ;
        RECT 232.395 -107.605 232.725 -107.275 ;
        RECT 232.395 -108.965 232.725 -108.635 ;
        RECT 232.395 -110.325 232.725 -109.995 ;
        RECT 232.395 -111.685 232.725 -111.355 ;
        RECT 232.395 -113.045 232.725 -112.715 ;
        RECT 232.395 -114.405 232.725 -114.075 ;
        RECT 232.395 -115.765 232.725 -115.435 ;
        RECT 232.395 -117.125 232.725 -116.795 ;
        RECT 232.395 -118.485 232.725 -118.155 ;
        RECT 232.395 -119.845 232.725 -119.515 ;
        RECT 232.395 -121.205 232.725 -120.875 ;
        RECT 232.395 -122.565 232.725 -122.235 ;
        RECT 232.395 -123.925 232.725 -123.595 ;
        RECT 232.395 -125.285 232.725 -124.955 ;
        RECT 232.395 -126.645 232.725 -126.315 ;
        RECT 232.395 -128.005 232.725 -127.675 ;
        RECT 232.395 -129.365 232.725 -129.035 ;
        RECT 232.395 -130.725 232.725 -130.395 ;
        RECT 232.395 -132.085 232.725 -131.755 ;
        RECT 232.395 -133.445 232.725 -133.115 ;
        RECT 232.395 -134.805 232.725 -134.475 ;
        RECT 232.395 -136.165 232.725 -135.835 ;
        RECT 232.395 -137.525 232.725 -137.195 ;
        RECT 232.395 -138.885 232.725 -138.555 ;
        RECT 232.395 -140.245 232.725 -139.915 ;
        RECT 232.395 -141.605 232.725 -141.275 ;
        RECT 232.395 -142.965 232.725 -142.635 ;
        RECT 232.395 -144.325 232.725 -143.995 ;
        RECT 232.395 -145.685 232.725 -145.355 ;
        RECT 232.395 -147.045 232.725 -146.715 ;
        RECT 232.395 -148.405 232.725 -148.075 ;
        RECT 232.395 -149.765 232.725 -149.435 ;
        RECT 232.395 -151.125 232.725 -150.795 ;
        RECT 232.395 -152.485 232.725 -152.155 ;
        RECT 232.395 -153.845 232.725 -153.515 ;
        RECT 232.395 -155.205 232.725 -154.875 ;
        RECT 232.395 -156.565 232.725 -156.235 ;
        RECT 232.395 -157.925 232.725 -157.595 ;
        RECT 232.395 -159.285 232.725 -158.955 ;
        RECT 232.395 -160.645 232.725 -160.315 ;
        RECT 232.395 -162.005 232.725 -161.675 ;
        RECT 232.395 -163.365 232.725 -163.035 ;
        RECT 232.395 -164.725 232.725 -164.395 ;
        RECT 232.395 -166.085 232.725 -165.755 ;
        RECT 232.395 -167.445 232.725 -167.115 ;
        RECT 232.395 -168.805 232.725 -168.475 ;
        RECT 232.395 -170.165 232.725 -169.835 ;
        RECT 232.395 -171.525 232.725 -171.195 ;
        RECT 232.395 -172.885 232.725 -172.555 ;
        RECT 232.395 -174.245 232.725 -173.915 ;
        RECT 232.395 -175.605 232.725 -175.275 ;
        RECT 232.395 -176.965 232.725 -176.635 ;
        RECT 232.395 -178.325 232.725 -177.995 ;
        RECT 232.395 -180.57 232.725 -179.44 ;
        RECT 232.4 -180.685 232.72 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 233.755 241.32 234.085 242.45 ;
        RECT 233.755 239.195 234.085 239.525 ;
        RECT 233.755 237.835 234.085 238.165 ;
        RECT 233.76 237.16 234.08 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 233.755 -1.525 234.085 -1.195 ;
        RECT 233.755 -2.885 234.085 -2.555 ;
        RECT 233.76 -3.56 234.08 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 233.755 -91.285 234.085 -90.955 ;
        RECT 233.755 -92.645 234.085 -92.315 ;
        RECT 233.755 -94.005 234.085 -93.675 ;
        RECT 233.755 -95.365 234.085 -95.035 ;
        RECT 233.755 -96.725 234.085 -96.395 ;
        RECT 233.755 -98.085 234.085 -97.755 ;
        RECT 233.755 -99.445 234.085 -99.115 ;
        RECT 233.755 -100.805 234.085 -100.475 ;
        RECT 233.755 -102.165 234.085 -101.835 ;
        RECT 233.755 -103.525 234.085 -103.195 ;
        RECT 233.755 -104.885 234.085 -104.555 ;
        RECT 233.755 -106.245 234.085 -105.915 ;
        RECT 233.755 -107.605 234.085 -107.275 ;
        RECT 233.755 -108.965 234.085 -108.635 ;
        RECT 233.755 -110.325 234.085 -109.995 ;
        RECT 233.755 -111.685 234.085 -111.355 ;
        RECT 233.755 -113.045 234.085 -112.715 ;
        RECT 233.755 -114.405 234.085 -114.075 ;
        RECT 233.755 -115.765 234.085 -115.435 ;
        RECT 233.755 -117.125 234.085 -116.795 ;
        RECT 233.755 -118.485 234.085 -118.155 ;
        RECT 233.755 -119.845 234.085 -119.515 ;
        RECT 233.755 -121.205 234.085 -120.875 ;
        RECT 233.755 -122.565 234.085 -122.235 ;
        RECT 233.755 -123.925 234.085 -123.595 ;
        RECT 233.755 -125.285 234.085 -124.955 ;
        RECT 233.755 -126.645 234.085 -126.315 ;
        RECT 233.755 -128.005 234.085 -127.675 ;
        RECT 233.755 -129.365 234.085 -129.035 ;
        RECT 233.755 -130.725 234.085 -130.395 ;
        RECT 233.755 -132.085 234.085 -131.755 ;
        RECT 233.755 -133.445 234.085 -133.115 ;
        RECT 233.755 -134.805 234.085 -134.475 ;
        RECT 233.755 -136.165 234.085 -135.835 ;
        RECT 233.755 -137.525 234.085 -137.195 ;
        RECT 233.755 -138.885 234.085 -138.555 ;
        RECT 233.755 -140.245 234.085 -139.915 ;
        RECT 233.755 -141.605 234.085 -141.275 ;
        RECT 233.755 -142.965 234.085 -142.635 ;
        RECT 233.755 -144.325 234.085 -143.995 ;
        RECT 233.755 -145.685 234.085 -145.355 ;
        RECT 233.755 -147.045 234.085 -146.715 ;
        RECT 233.755 -148.405 234.085 -148.075 ;
        RECT 233.755 -149.765 234.085 -149.435 ;
        RECT 233.755 -151.125 234.085 -150.795 ;
        RECT 233.755 -152.485 234.085 -152.155 ;
        RECT 233.755 -153.845 234.085 -153.515 ;
        RECT 233.755 -155.205 234.085 -154.875 ;
        RECT 233.755 -156.565 234.085 -156.235 ;
        RECT 233.755 -157.925 234.085 -157.595 ;
        RECT 233.755 -159.285 234.085 -158.955 ;
        RECT 233.755 -160.645 234.085 -160.315 ;
        RECT 233.755 -162.005 234.085 -161.675 ;
        RECT 233.755 -163.365 234.085 -163.035 ;
        RECT 233.755 -164.725 234.085 -164.395 ;
        RECT 233.755 -166.085 234.085 -165.755 ;
        RECT 233.755 -167.445 234.085 -167.115 ;
        RECT 233.755 -168.805 234.085 -168.475 ;
        RECT 233.755 -170.165 234.085 -169.835 ;
        RECT 233.755 -171.525 234.085 -171.195 ;
        RECT 233.755 -172.885 234.085 -172.555 ;
        RECT 233.755 -174.245 234.085 -173.915 ;
        RECT 233.755 -175.605 234.085 -175.275 ;
        RECT 233.755 -176.965 234.085 -176.635 ;
        RECT 233.755 -178.325 234.085 -177.995 ;
        RECT 233.755 -180.57 234.085 -179.44 ;
        RECT 233.76 -180.685 234.08 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 235.11 -94.075 235.44 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 235.115 241.32 235.445 242.45 ;
        RECT 235.115 239.195 235.445 239.525 ;
        RECT 235.115 237.835 235.445 238.165 ;
        RECT 235.12 237.16 235.44 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 235.115 -176.965 235.445 -176.635 ;
        RECT 235.115 -178.325 235.445 -177.995 ;
        RECT 235.115 -180.57 235.445 -179.44 ;
        RECT 235.12 -180.685 235.44 -95.035 ;
        RECT 235.115 -95.365 235.445 -95.035 ;
        RECT 235.115 -96.725 235.445 -96.395 ;
        RECT 235.115 -98.085 235.445 -97.755 ;
        RECT 235.115 -99.445 235.445 -99.115 ;
        RECT 235.115 -100.805 235.445 -100.475 ;
        RECT 235.115 -102.165 235.445 -101.835 ;
        RECT 235.115 -103.525 235.445 -103.195 ;
        RECT 235.115 -104.885 235.445 -104.555 ;
        RECT 235.115 -106.245 235.445 -105.915 ;
        RECT 235.115 -107.605 235.445 -107.275 ;
        RECT 235.115 -108.965 235.445 -108.635 ;
        RECT 235.115 -110.325 235.445 -109.995 ;
        RECT 235.115 -111.685 235.445 -111.355 ;
        RECT 235.115 -113.045 235.445 -112.715 ;
        RECT 235.115 -114.405 235.445 -114.075 ;
        RECT 235.115 -115.765 235.445 -115.435 ;
        RECT 235.115 -117.125 235.445 -116.795 ;
        RECT 235.115 -118.485 235.445 -118.155 ;
        RECT 235.115 -119.845 235.445 -119.515 ;
        RECT 235.115 -121.205 235.445 -120.875 ;
        RECT 235.115 -122.565 235.445 -122.235 ;
        RECT 235.115 -123.925 235.445 -123.595 ;
        RECT 235.115 -125.285 235.445 -124.955 ;
        RECT 235.115 -126.645 235.445 -126.315 ;
        RECT 235.115 -128.005 235.445 -127.675 ;
        RECT 235.115 -129.365 235.445 -129.035 ;
        RECT 235.115 -130.725 235.445 -130.395 ;
        RECT 235.115 -132.085 235.445 -131.755 ;
        RECT 235.115 -133.445 235.445 -133.115 ;
        RECT 235.115 -134.805 235.445 -134.475 ;
        RECT 235.115 -136.165 235.445 -135.835 ;
        RECT 235.115 -137.525 235.445 -137.195 ;
        RECT 235.115 -138.885 235.445 -138.555 ;
        RECT 235.115 -140.245 235.445 -139.915 ;
        RECT 235.115 -141.605 235.445 -141.275 ;
        RECT 235.115 -142.965 235.445 -142.635 ;
        RECT 235.115 -144.325 235.445 -143.995 ;
        RECT 235.115 -145.685 235.445 -145.355 ;
        RECT 235.115 -147.045 235.445 -146.715 ;
        RECT 235.115 -148.405 235.445 -148.075 ;
        RECT 235.115 -149.765 235.445 -149.435 ;
        RECT 235.115 -151.125 235.445 -150.795 ;
        RECT 235.115 -152.485 235.445 -152.155 ;
        RECT 235.115 -153.845 235.445 -153.515 ;
        RECT 235.115 -155.205 235.445 -154.875 ;
        RECT 235.115 -156.565 235.445 -156.235 ;
        RECT 235.115 -157.925 235.445 -157.595 ;
        RECT 235.115 -159.285 235.445 -158.955 ;
        RECT 235.115 -160.645 235.445 -160.315 ;
        RECT 235.115 -162.005 235.445 -161.675 ;
        RECT 235.115 -163.365 235.445 -163.035 ;
        RECT 235.115 -164.725 235.445 -164.395 ;
        RECT 235.115 -166.085 235.445 -165.755 ;
        RECT 235.115 -167.445 235.445 -167.115 ;
        RECT 235.115 -168.805 235.445 -168.475 ;
        RECT 235.115 -170.165 235.445 -169.835 ;
        RECT 235.115 -171.525 235.445 -171.195 ;
        RECT 235.115 -172.885 235.445 -172.555 ;
        RECT 235.115 -174.245 235.445 -173.915 ;
        RECT 235.115 -175.605 235.445 -175.275 ;
    END
    PORT
      LAYER met3 ;
        RECT 173.915 241.32 174.245 242.45 ;
        RECT 173.915 239.195 174.245 239.525 ;
        RECT 173.915 237.835 174.245 238.165 ;
        RECT 173.92 237.16 174.24 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 173.915 -95.365 174.245 -95.035 ;
        RECT 173.915 -96.725 174.245 -96.395 ;
        RECT 173.915 -98.085 174.245 -97.755 ;
        RECT 173.915 -99.445 174.245 -99.115 ;
        RECT 173.915 -100.805 174.245 -100.475 ;
        RECT 173.915 -102.165 174.245 -101.835 ;
        RECT 173.915 -103.525 174.245 -103.195 ;
        RECT 173.915 -104.885 174.245 -104.555 ;
        RECT 173.915 -106.245 174.245 -105.915 ;
        RECT 173.915 -107.605 174.245 -107.275 ;
        RECT 173.915 -108.965 174.245 -108.635 ;
        RECT 173.915 -110.325 174.245 -109.995 ;
        RECT 173.915 -111.685 174.245 -111.355 ;
        RECT 173.915 -113.045 174.245 -112.715 ;
        RECT 173.915 -114.405 174.245 -114.075 ;
        RECT 173.915 -115.765 174.245 -115.435 ;
        RECT 173.915 -117.125 174.245 -116.795 ;
        RECT 173.915 -118.485 174.245 -118.155 ;
        RECT 173.915 -119.845 174.245 -119.515 ;
        RECT 173.915 -121.205 174.245 -120.875 ;
        RECT 173.915 -122.565 174.245 -122.235 ;
        RECT 173.915 -123.925 174.245 -123.595 ;
        RECT 173.915 -125.285 174.245 -124.955 ;
        RECT 173.915 -126.645 174.245 -126.315 ;
        RECT 173.915 -128.005 174.245 -127.675 ;
        RECT 173.915 -129.365 174.245 -129.035 ;
        RECT 173.915 -130.725 174.245 -130.395 ;
        RECT 173.915 -132.085 174.245 -131.755 ;
        RECT 173.915 -133.445 174.245 -133.115 ;
        RECT 173.915 -134.805 174.245 -134.475 ;
        RECT 173.915 -136.165 174.245 -135.835 ;
        RECT 173.915 -137.525 174.245 -137.195 ;
        RECT 173.915 -138.885 174.245 -138.555 ;
        RECT 173.915 -140.245 174.245 -139.915 ;
        RECT 173.915 -141.605 174.245 -141.275 ;
        RECT 173.915 -142.965 174.245 -142.635 ;
        RECT 173.915 -144.325 174.245 -143.995 ;
        RECT 173.915 -145.685 174.245 -145.355 ;
        RECT 173.915 -147.045 174.245 -146.715 ;
        RECT 173.915 -148.405 174.245 -148.075 ;
        RECT 173.915 -149.765 174.245 -149.435 ;
        RECT 173.915 -151.125 174.245 -150.795 ;
        RECT 173.915 -152.485 174.245 -152.155 ;
        RECT 173.915 -153.845 174.245 -153.515 ;
        RECT 173.915 -155.205 174.245 -154.875 ;
        RECT 173.915 -156.565 174.245 -156.235 ;
        RECT 173.915 -157.925 174.245 -157.595 ;
        RECT 173.915 -159.285 174.245 -158.955 ;
        RECT 173.915 -160.645 174.245 -160.315 ;
        RECT 173.915 -162.005 174.245 -161.675 ;
        RECT 173.915 -163.365 174.245 -163.035 ;
        RECT 173.915 -164.725 174.245 -164.395 ;
        RECT 173.915 -166.085 174.245 -165.755 ;
        RECT 173.915 -167.445 174.245 -167.115 ;
        RECT 173.915 -168.805 174.245 -168.475 ;
        RECT 173.915 -170.165 174.245 -169.835 ;
        RECT 173.915 -171.525 174.245 -171.195 ;
        RECT 173.915 -172.885 174.245 -172.555 ;
        RECT 173.915 -174.245 174.245 -173.915 ;
        RECT 173.915 -175.605 174.245 -175.275 ;
        RECT 173.915 -176.965 174.245 -176.635 ;
        RECT 173.915 -178.325 174.245 -177.995 ;
        RECT 173.915 -180.57 174.245 -179.44 ;
        RECT 173.92 -180.685 174.24 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 174.11 -94.075 174.44 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 175.275 241.32 175.605 242.45 ;
        RECT 175.275 239.195 175.605 239.525 ;
        RECT 175.275 237.835 175.605 238.165 ;
        RECT 175.28 237.16 175.6 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 175.275 -1.525 175.605 -1.195 ;
        RECT 175.275 -2.885 175.605 -2.555 ;
        RECT 175.28 -3.56 175.6 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 176.635 241.32 176.965 242.45 ;
        RECT 176.635 239.195 176.965 239.525 ;
        RECT 176.635 237.835 176.965 238.165 ;
        RECT 176.64 237.16 176.96 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 176.635 -1.525 176.965 -1.195 ;
        RECT 176.635 -2.885 176.965 -2.555 ;
        RECT 176.64 -3.56 176.96 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 177.995 241.32 178.325 242.45 ;
        RECT 177.995 239.195 178.325 239.525 ;
        RECT 177.995 237.835 178.325 238.165 ;
        RECT 178 237.16 178.32 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 177.995 -1.525 178.325 -1.195 ;
        RECT 177.995 -2.885 178.325 -2.555 ;
        RECT 178 -3.56 178.32 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 177.995 -91.285 178.325 -90.955 ;
        RECT 177.995 -92.645 178.325 -92.315 ;
        RECT 177.995 -94.005 178.325 -93.675 ;
        RECT 177.995 -95.365 178.325 -95.035 ;
        RECT 177.995 -96.725 178.325 -96.395 ;
        RECT 177.995 -98.085 178.325 -97.755 ;
        RECT 177.995 -99.445 178.325 -99.115 ;
        RECT 177.995 -100.805 178.325 -100.475 ;
        RECT 177.995 -102.165 178.325 -101.835 ;
        RECT 177.995 -103.525 178.325 -103.195 ;
        RECT 177.995 -104.885 178.325 -104.555 ;
        RECT 177.995 -106.245 178.325 -105.915 ;
        RECT 177.995 -107.605 178.325 -107.275 ;
        RECT 177.995 -108.965 178.325 -108.635 ;
        RECT 177.995 -110.325 178.325 -109.995 ;
        RECT 177.995 -111.685 178.325 -111.355 ;
        RECT 177.995 -113.045 178.325 -112.715 ;
        RECT 177.995 -114.405 178.325 -114.075 ;
        RECT 177.995 -115.765 178.325 -115.435 ;
        RECT 177.995 -117.125 178.325 -116.795 ;
        RECT 177.995 -118.485 178.325 -118.155 ;
        RECT 177.995 -119.845 178.325 -119.515 ;
        RECT 177.995 -121.205 178.325 -120.875 ;
        RECT 177.995 -122.565 178.325 -122.235 ;
        RECT 177.995 -123.925 178.325 -123.595 ;
        RECT 177.995 -125.285 178.325 -124.955 ;
        RECT 177.995 -126.645 178.325 -126.315 ;
        RECT 177.995 -128.005 178.325 -127.675 ;
        RECT 177.995 -129.365 178.325 -129.035 ;
        RECT 177.995 -130.725 178.325 -130.395 ;
        RECT 177.995 -132.085 178.325 -131.755 ;
        RECT 177.995 -133.445 178.325 -133.115 ;
        RECT 177.995 -134.805 178.325 -134.475 ;
        RECT 177.995 -136.165 178.325 -135.835 ;
        RECT 177.995 -137.525 178.325 -137.195 ;
        RECT 177.995 -138.885 178.325 -138.555 ;
        RECT 177.995 -140.245 178.325 -139.915 ;
        RECT 177.995 -141.605 178.325 -141.275 ;
        RECT 177.995 -142.965 178.325 -142.635 ;
        RECT 177.995 -144.325 178.325 -143.995 ;
        RECT 177.995 -145.685 178.325 -145.355 ;
        RECT 177.995 -147.045 178.325 -146.715 ;
        RECT 177.995 -148.405 178.325 -148.075 ;
        RECT 177.995 -149.765 178.325 -149.435 ;
        RECT 177.995 -151.125 178.325 -150.795 ;
        RECT 177.995 -152.485 178.325 -152.155 ;
        RECT 177.995 -153.845 178.325 -153.515 ;
        RECT 177.995 -155.205 178.325 -154.875 ;
        RECT 177.995 -156.565 178.325 -156.235 ;
        RECT 177.995 -157.925 178.325 -157.595 ;
        RECT 177.995 -159.285 178.325 -158.955 ;
        RECT 177.995 -160.645 178.325 -160.315 ;
        RECT 177.995 -162.005 178.325 -161.675 ;
        RECT 177.995 -163.365 178.325 -163.035 ;
        RECT 177.995 -164.725 178.325 -164.395 ;
        RECT 177.995 -166.085 178.325 -165.755 ;
        RECT 177.995 -167.445 178.325 -167.115 ;
        RECT 177.995 -168.805 178.325 -168.475 ;
        RECT 177.995 -170.165 178.325 -169.835 ;
        RECT 177.995 -171.525 178.325 -171.195 ;
        RECT 177.995 -172.885 178.325 -172.555 ;
        RECT 177.995 -174.245 178.325 -173.915 ;
        RECT 177.995 -175.605 178.325 -175.275 ;
        RECT 177.995 -176.965 178.325 -176.635 ;
        RECT 177.995 -178.325 178.325 -177.995 ;
        RECT 177.995 -180.57 178.325 -179.44 ;
        RECT 178 -180.685 178.32 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 179.355 241.32 179.685 242.45 ;
        RECT 179.355 239.195 179.685 239.525 ;
        RECT 179.355 237.835 179.685 238.165 ;
        RECT 179.36 237.16 179.68 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 179.355 -95.365 179.685 -95.035 ;
        RECT 179.355 -96.725 179.685 -96.395 ;
        RECT 179.355 -98.085 179.685 -97.755 ;
        RECT 179.355 -99.445 179.685 -99.115 ;
        RECT 179.355 -100.805 179.685 -100.475 ;
        RECT 179.355 -102.165 179.685 -101.835 ;
        RECT 179.355 -103.525 179.685 -103.195 ;
        RECT 179.355 -104.885 179.685 -104.555 ;
        RECT 179.355 -106.245 179.685 -105.915 ;
        RECT 179.355 -107.605 179.685 -107.275 ;
        RECT 179.355 -108.965 179.685 -108.635 ;
        RECT 179.355 -110.325 179.685 -109.995 ;
        RECT 179.355 -111.685 179.685 -111.355 ;
        RECT 179.355 -113.045 179.685 -112.715 ;
        RECT 179.355 -114.405 179.685 -114.075 ;
        RECT 179.355 -115.765 179.685 -115.435 ;
        RECT 179.355 -117.125 179.685 -116.795 ;
        RECT 179.355 -118.485 179.685 -118.155 ;
        RECT 179.355 -119.845 179.685 -119.515 ;
        RECT 179.355 -121.205 179.685 -120.875 ;
        RECT 179.355 -122.565 179.685 -122.235 ;
        RECT 179.355 -123.925 179.685 -123.595 ;
        RECT 179.355 -125.285 179.685 -124.955 ;
        RECT 179.355 -126.645 179.685 -126.315 ;
        RECT 179.355 -128.005 179.685 -127.675 ;
        RECT 179.355 -129.365 179.685 -129.035 ;
        RECT 179.355 -130.725 179.685 -130.395 ;
        RECT 179.355 -132.085 179.685 -131.755 ;
        RECT 179.355 -133.445 179.685 -133.115 ;
        RECT 179.355 -134.805 179.685 -134.475 ;
        RECT 179.355 -136.165 179.685 -135.835 ;
        RECT 179.355 -137.525 179.685 -137.195 ;
        RECT 179.355 -138.885 179.685 -138.555 ;
        RECT 179.355 -140.245 179.685 -139.915 ;
        RECT 179.355 -141.605 179.685 -141.275 ;
        RECT 179.355 -142.965 179.685 -142.635 ;
        RECT 179.355 -144.325 179.685 -143.995 ;
        RECT 179.355 -145.685 179.685 -145.355 ;
        RECT 179.355 -147.045 179.685 -146.715 ;
        RECT 179.355 -148.405 179.685 -148.075 ;
        RECT 179.355 -149.765 179.685 -149.435 ;
        RECT 179.355 -151.125 179.685 -150.795 ;
        RECT 179.355 -152.485 179.685 -152.155 ;
        RECT 179.355 -153.845 179.685 -153.515 ;
        RECT 179.355 -155.205 179.685 -154.875 ;
        RECT 179.355 -156.565 179.685 -156.235 ;
        RECT 179.355 -157.925 179.685 -157.595 ;
        RECT 179.355 -159.285 179.685 -158.955 ;
        RECT 179.355 -160.645 179.685 -160.315 ;
        RECT 179.355 -162.005 179.685 -161.675 ;
        RECT 179.355 -163.365 179.685 -163.035 ;
        RECT 179.355 -164.725 179.685 -164.395 ;
        RECT 179.355 -166.085 179.685 -165.755 ;
        RECT 179.355 -167.445 179.685 -167.115 ;
        RECT 179.355 -168.805 179.685 -168.475 ;
        RECT 179.355 -170.165 179.685 -169.835 ;
        RECT 179.355 -171.525 179.685 -171.195 ;
        RECT 179.355 -172.885 179.685 -172.555 ;
        RECT 179.355 -174.245 179.685 -173.915 ;
        RECT 179.355 -175.605 179.685 -175.275 ;
        RECT 179.355 -176.965 179.685 -176.635 ;
        RECT 179.355 -178.325 179.685 -177.995 ;
        RECT 179.355 -180.57 179.685 -179.44 ;
        RECT 179.36 -180.685 179.68 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 180.21 -94.075 180.54 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 180.715 241.32 181.045 242.45 ;
        RECT 180.715 239.195 181.045 239.525 ;
        RECT 180.715 237.835 181.045 238.165 ;
        RECT 180.72 237.16 181.04 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 182.075 241.32 182.405 242.45 ;
        RECT 182.075 239.195 182.405 239.525 ;
        RECT 182.075 237.835 182.405 238.165 ;
        RECT 182.08 237.16 182.4 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 182.075 -1.525 182.405 -1.195 ;
        RECT 182.075 -2.885 182.405 -2.555 ;
        RECT 182.08 -3.56 182.4 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 183.435 241.32 183.765 242.45 ;
        RECT 183.435 239.195 183.765 239.525 ;
        RECT 183.435 237.835 183.765 238.165 ;
        RECT 183.44 237.16 183.76 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 183.435 -1.525 183.765 -1.195 ;
        RECT 183.435 -2.885 183.765 -2.555 ;
        RECT 183.44 -3.56 183.76 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 183.435 -91.285 183.765 -90.955 ;
        RECT 183.435 -92.645 183.765 -92.315 ;
        RECT 183.435 -94.005 183.765 -93.675 ;
        RECT 183.435 -95.365 183.765 -95.035 ;
        RECT 183.435 -96.725 183.765 -96.395 ;
        RECT 183.435 -98.085 183.765 -97.755 ;
        RECT 183.435 -99.445 183.765 -99.115 ;
        RECT 183.435 -100.805 183.765 -100.475 ;
        RECT 183.435 -102.165 183.765 -101.835 ;
        RECT 183.435 -103.525 183.765 -103.195 ;
        RECT 183.435 -104.885 183.765 -104.555 ;
        RECT 183.435 -106.245 183.765 -105.915 ;
        RECT 183.435 -107.605 183.765 -107.275 ;
        RECT 183.435 -108.965 183.765 -108.635 ;
        RECT 183.435 -110.325 183.765 -109.995 ;
        RECT 183.435 -111.685 183.765 -111.355 ;
        RECT 183.435 -113.045 183.765 -112.715 ;
        RECT 183.435 -114.405 183.765 -114.075 ;
        RECT 183.435 -115.765 183.765 -115.435 ;
        RECT 183.435 -117.125 183.765 -116.795 ;
        RECT 183.435 -118.485 183.765 -118.155 ;
        RECT 183.435 -119.845 183.765 -119.515 ;
        RECT 183.435 -121.205 183.765 -120.875 ;
        RECT 183.435 -122.565 183.765 -122.235 ;
        RECT 183.435 -123.925 183.765 -123.595 ;
        RECT 183.435 -125.285 183.765 -124.955 ;
        RECT 183.435 -126.645 183.765 -126.315 ;
        RECT 183.435 -128.005 183.765 -127.675 ;
        RECT 183.435 -129.365 183.765 -129.035 ;
        RECT 183.435 -130.725 183.765 -130.395 ;
        RECT 183.435 -132.085 183.765 -131.755 ;
        RECT 183.435 -133.445 183.765 -133.115 ;
        RECT 183.435 -134.805 183.765 -134.475 ;
        RECT 183.435 -136.165 183.765 -135.835 ;
        RECT 183.435 -137.525 183.765 -137.195 ;
        RECT 183.435 -138.885 183.765 -138.555 ;
        RECT 183.435 -140.245 183.765 -139.915 ;
        RECT 183.435 -141.605 183.765 -141.275 ;
        RECT 183.435 -142.965 183.765 -142.635 ;
        RECT 183.435 -144.325 183.765 -143.995 ;
        RECT 183.435 -145.685 183.765 -145.355 ;
        RECT 183.435 -147.045 183.765 -146.715 ;
        RECT 183.435 -148.405 183.765 -148.075 ;
        RECT 183.435 -149.765 183.765 -149.435 ;
        RECT 183.435 -151.125 183.765 -150.795 ;
        RECT 183.435 -152.485 183.765 -152.155 ;
        RECT 183.435 -153.845 183.765 -153.515 ;
        RECT 183.435 -155.205 183.765 -154.875 ;
        RECT 183.435 -156.565 183.765 -156.235 ;
        RECT 183.435 -157.925 183.765 -157.595 ;
        RECT 183.435 -159.285 183.765 -158.955 ;
        RECT 183.435 -160.645 183.765 -160.315 ;
        RECT 183.435 -162.005 183.765 -161.675 ;
        RECT 183.435 -163.365 183.765 -163.035 ;
        RECT 183.435 -164.725 183.765 -164.395 ;
        RECT 183.435 -166.085 183.765 -165.755 ;
        RECT 183.435 -167.445 183.765 -167.115 ;
        RECT 183.435 -168.805 183.765 -168.475 ;
        RECT 183.435 -170.165 183.765 -169.835 ;
        RECT 183.435 -171.525 183.765 -171.195 ;
        RECT 183.435 -172.885 183.765 -172.555 ;
        RECT 183.435 -174.245 183.765 -173.915 ;
        RECT 183.435 -175.605 183.765 -175.275 ;
        RECT 183.435 -176.965 183.765 -176.635 ;
        RECT 183.435 -178.325 183.765 -177.995 ;
        RECT 183.435 -180.57 183.765 -179.44 ;
        RECT 183.44 -180.685 183.76 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 184.795 241.32 185.125 242.45 ;
        RECT 184.795 239.195 185.125 239.525 ;
        RECT 184.795 237.835 185.125 238.165 ;
        RECT 184.8 237.16 185.12 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 184.795 -1.525 185.125 -1.195 ;
        RECT 184.795 -2.885 185.125 -2.555 ;
        RECT 184.8 -3.56 185.12 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 184.795 -91.285 185.125 -90.955 ;
        RECT 184.795 -92.645 185.125 -92.315 ;
        RECT 184.795 -94.005 185.125 -93.675 ;
        RECT 184.795 -95.365 185.125 -95.035 ;
        RECT 184.795 -96.725 185.125 -96.395 ;
        RECT 184.795 -98.085 185.125 -97.755 ;
        RECT 184.795 -99.445 185.125 -99.115 ;
        RECT 184.795 -100.805 185.125 -100.475 ;
        RECT 184.795 -102.165 185.125 -101.835 ;
        RECT 184.795 -103.525 185.125 -103.195 ;
        RECT 184.795 -104.885 185.125 -104.555 ;
        RECT 184.795 -106.245 185.125 -105.915 ;
        RECT 184.795 -107.605 185.125 -107.275 ;
        RECT 184.795 -108.965 185.125 -108.635 ;
        RECT 184.795 -110.325 185.125 -109.995 ;
        RECT 184.795 -111.685 185.125 -111.355 ;
        RECT 184.795 -113.045 185.125 -112.715 ;
        RECT 184.795 -114.405 185.125 -114.075 ;
        RECT 184.795 -115.765 185.125 -115.435 ;
        RECT 184.795 -117.125 185.125 -116.795 ;
        RECT 184.795 -118.485 185.125 -118.155 ;
        RECT 184.795 -119.845 185.125 -119.515 ;
        RECT 184.795 -121.205 185.125 -120.875 ;
        RECT 184.795 -122.565 185.125 -122.235 ;
        RECT 184.795 -123.925 185.125 -123.595 ;
        RECT 184.795 -125.285 185.125 -124.955 ;
        RECT 184.795 -126.645 185.125 -126.315 ;
        RECT 184.795 -128.005 185.125 -127.675 ;
        RECT 184.795 -129.365 185.125 -129.035 ;
        RECT 184.795 -130.725 185.125 -130.395 ;
        RECT 184.795 -132.085 185.125 -131.755 ;
        RECT 184.795 -133.445 185.125 -133.115 ;
        RECT 184.795 -134.805 185.125 -134.475 ;
        RECT 184.795 -136.165 185.125 -135.835 ;
        RECT 184.795 -137.525 185.125 -137.195 ;
        RECT 184.795 -138.885 185.125 -138.555 ;
        RECT 184.795 -140.245 185.125 -139.915 ;
        RECT 184.795 -141.605 185.125 -141.275 ;
        RECT 184.795 -142.965 185.125 -142.635 ;
        RECT 184.795 -144.325 185.125 -143.995 ;
        RECT 184.795 -145.685 185.125 -145.355 ;
        RECT 184.795 -147.045 185.125 -146.715 ;
        RECT 184.795 -148.405 185.125 -148.075 ;
        RECT 184.795 -149.765 185.125 -149.435 ;
        RECT 184.795 -151.125 185.125 -150.795 ;
        RECT 184.795 -152.485 185.125 -152.155 ;
        RECT 184.795 -153.845 185.125 -153.515 ;
        RECT 184.795 -155.205 185.125 -154.875 ;
        RECT 184.795 -156.565 185.125 -156.235 ;
        RECT 184.795 -157.925 185.125 -157.595 ;
        RECT 184.795 -159.285 185.125 -158.955 ;
        RECT 184.795 -160.645 185.125 -160.315 ;
        RECT 184.795 -162.005 185.125 -161.675 ;
        RECT 184.795 -163.365 185.125 -163.035 ;
        RECT 184.795 -164.725 185.125 -164.395 ;
        RECT 184.795 -166.085 185.125 -165.755 ;
        RECT 184.795 -167.445 185.125 -167.115 ;
        RECT 184.795 -168.805 185.125 -168.475 ;
        RECT 184.795 -170.165 185.125 -169.835 ;
        RECT 184.795 -171.525 185.125 -171.195 ;
        RECT 184.795 -172.885 185.125 -172.555 ;
        RECT 184.795 -174.245 185.125 -173.915 ;
        RECT 184.795 -175.605 185.125 -175.275 ;
        RECT 184.795 -176.965 185.125 -176.635 ;
        RECT 184.795 -178.325 185.125 -177.995 ;
        RECT 184.795 -180.57 185.125 -179.44 ;
        RECT 184.8 -180.685 185.12 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 186.155 241.32 186.485 242.45 ;
        RECT 186.155 239.195 186.485 239.525 ;
        RECT 186.155 237.835 186.485 238.165 ;
        RECT 186.16 237.16 186.48 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 186.155 -95.365 186.485 -95.035 ;
        RECT 186.155 -96.725 186.485 -96.395 ;
        RECT 186.155 -98.085 186.485 -97.755 ;
        RECT 186.155 -99.445 186.485 -99.115 ;
        RECT 186.155 -100.805 186.485 -100.475 ;
        RECT 186.155 -102.165 186.485 -101.835 ;
        RECT 186.155 -103.525 186.485 -103.195 ;
        RECT 186.155 -104.885 186.485 -104.555 ;
        RECT 186.155 -106.245 186.485 -105.915 ;
        RECT 186.155 -107.605 186.485 -107.275 ;
        RECT 186.155 -108.965 186.485 -108.635 ;
        RECT 186.155 -110.325 186.485 -109.995 ;
        RECT 186.155 -111.685 186.485 -111.355 ;
        RECT 186.155 -113.045 186.485 -112.715 ;
        RECT 186.155 -114.405 186.485 -114.075 ;
        RECT 186.155 -115.765 186.485 -115.435 ;
        RECT 186.155 -117.125 186.485 -116.795 ;
        RECT 186.155 -118.485 186.485 -118.155 ;
        RECT 186.155 -119.845 186.485 -119.515 ;
        RECT 186.155 -121.205 186.485 -120.875 ;
        RECT 186.155 -122.565 186.485 -122.235 ;
        RECT 186.155 -123.925 186.485 -123.595 ;
        RECT 186.155 -125.285 186.485 -124.955 ;
        RECT 186.155 -126.645 186.485 -126.315 ;
        RECT 186.155 -128.005 186.485 -127.675 ;
        RECT 186.155 -129.365 186.485 -129.035 ;
        RECT 186.155 -130.725 186.485 -130.395 ;
        RECT 186.155 -132.085 186.485 -131.755 ;
        RECT 186.155 -133.445 186.485 -133.115 ;
        RECT 186.155 -134.805 186.485 -134.475 ;
        RECT 186.155 -136.165 186.485 -135.835 ;
        RECT 186.155 -137.525 186.485 -137.195 ;
        RECT 186.155 -138.885 186.485 -138.555 ;
        RECT 186.155 -140.245 186.485 -139.915 ;
        RECT 186.155 -141.605 186.485 -141.275 ;
        RECT 186.155 -142.965 186.485 -142.635 ;
        RECT 186.155 -144.325 186.485 -143.995 ;
        RECT 186.155 -145.685 186.485 -145.355 ;
        RECT 186.155 -147.045 186.485 -146.715 ;
        RECT 186.155 -148.405 186.485 -148.075 ;
        RECT 186.155 -149.765 186.485 -149.435 ;
        RECT 186.155 -151.125 186.485 -150.795 ;
        RECT 186.155 -152.485 186.485 -152.155 ;
        RECT 186.155 -153.845 186.485 -153.515 ;
        RECT 186.155 -155.205 186.485 -154.875 ;
        RECT 186.155 -156.565 186.485 -156.235 ;
        RECT 186.155 -157.925 186.485 -157.595 ;
        RECT 186.155 -159.285 186.485 -158.955 ;
        RECT 186.155 -160.645 186.485 -160.315 ;
        RECT 186.155 -162.005 186.485 -161.675 ;
        RECT 186.155 -163.365 186.485 -163.035 ;
        RECT 186.155 -164.725 186.485 -164.395 ;
        RECT 186.155 -166.085 186.485 -165.755 ;
        RECT 186.155 -167.445 186.485 -167.115 ;
        RECT 186.155 -168.805 186.485 -168.475 ;
        RECT 186.155 -170.165 186.485 -169.835 ;
        RECT 186.155 -171.525 186.485 -171.195 ;
        RECT 186.155 -172.885 186.485 -172.555 ;
        RECT 186.155 -174.245 186.485 -173.915 ;
        RECT 186.155 -175.605 186.485 -175.275 ;
        RECT 186.155 -176.965 186.485 -176.635 ;
        RECT 186.155 -178.325 186.485 -177.995 ;
        RECT 186.155 -180.57 186.485 -179.44 ;
        RECT 186.16 -180.685 186.48 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 186.31 -94.075 186.64 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 187.515 241.32 187.845 242.45 ;
        RECT 187.515 239.195 187.845 239.525 ;
        RECT 187.515 237.835 187.845 238.165 ;
        RECT 187.52 237.16 187.84 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 187.515 -1.525 187.845 -1.195 ;
        RECT 187.515 -2.885 187.845 -2.555 ;
        RECT 187.52 -3.56 187.84 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 188.875 241.32 189.205 242.45 ;
        RECT 188.875 239.195 189.205 239.525 ;
        RECT 188.875 237.835 189.205 238.165 ;
        RECT 188.88 237.16 189.2 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 188.875 -1.525 189.205 -1.195 ;
        RECT 188.875 -2.885 189.205 -2.555 ;
        RECT 188.88 -3.56 189.2 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 190.235 241.32 190.565 242.45 ;
        RECT 190.235 239.195 190.565 239.525 ;
        RECT 190.235 237.835 190.565 238.165 ;
        RECT 190.24 237.16 190.56 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 190.235 -1.525 190.565 -1.195 ;
        RECT 190.235 -2.885 190.565 -2.555 ;
        RECT 190.24 -3.56 190.56 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 190.235 -91.285 190.565 -90.955 ;
        RECT 190.235 -92.645 190.565 -92.315 ;
        RECT 190.235 -94.005 190.565 -93.675 ;
        RECT 190.235 -95.365 190.565 -95.035 ;
        RECT 190.235 -96.725 190.565 -96.395 ;
        RECT 190.235 -98.085 190.565 -97.755 ;
        RECT 190.235 -99.445 190.565 -99.115 ;
        RECT 190.235 -100.805 190.565 -100.475 ;
        RECT 190.235 -102.165 190.565 -101.835 ;
        RECT 190.235 -103.525 190.565 -103.195 ;
        RECT 190.235 -104.885 190.565 -104.555 ;
        RECT 190.235 -106.245 190.565 -105.915 ;
        RECT 190.235 -107.605 190.565 -107.275 ;
        RECT 190.235 -108.965 190.565 -108.635 ;
        RECT 190.235 -110.325 190.565 -109.995 ;
        RECT 190.235 -111.685 190.565 -111.355 ;
        RECT 190.235 -113.045 190.565 -112.715 ;
        RECT 190.235 -114.405 190.565 -114.075 ;
        RECT 190.235 -115.765 190.565 -115.435 ;
        RECT 190.235 -117.125 190.565 -116.795 ;
        RECT 190.235 -118.485 190.565 -118.155 ;
        RECT 190.235 -119.845 190.565 -119.515 ;
        RECT 190.235 -121.205 190.565 -120.875 ;
        RECT 190.235 -122.565 190.565 -122.235 ;
        RECT 190.235 -123.925 190.565 -123.595 ;
        RECT 190.235 -125.285 190.565 -124.955 ;
        RECT 190.235 -126.645 190.565 -126.315 ;
        RECT 190.235 -128.005 190.565 -127.675 ;
        RECT 190.235 -129.365 190.565 -129.035 ;
        RECT 190.235 -130.725 190.565 -130.395 ;
        RECT 190.235 -132.085 190.565 -131.755 ;
        RECT 190.235 -133.445 190.565 -133.115 ;
        RECT 190.235 -134.805 190.565 -134.475 ;
        RECT 190.235 -136.165 190.565 -135.835 ;
        RECT 190.235 -137.525 190.565 -137.195 ;
        RECT 190.235 -138.885 190.565 -138.555 ;
        RECT 190.235 -140.245 190.565 -139.915 ;
        RECT 190.235 -141.605 190.565 -141.275 ;
        RECT 190.235 -142.965 190.565 -142.635 ;
        RECT 190.235 -144.325 190.565 -143.995 ;
        RECT 190.235 -145.685 190.565 -145.355 ;
        RECT 190.235 -147.045 190.565 -146.715 ;
        RECT 190.235 -148.405 190.565 -148.075 ;
        RECT 190.235 -149.765 190.565 -149.435 ;
        RECT 190.235 -151.125 190.565 -150.795 ;
        RECT 190.235 -152.485 190.565 -152.155 ;
        RECT 190.235 -153.845 190.565 -153.515 ;
        RECT 190.235 -155.205 190.565 -154.875 ;
        RECT 190.235 -156.565 190.565 -156.235 ;
        RECT 190.235 -157.925 190.565 -157.595 ;
        RECT 190.235 -159.285 190.565 -158.955 ;
        RECT 190.235 -160.645 190.565 -160.315 ;
        RECT 190.235 -162.005 190.565 -161.675 ;
        RECT 190.235 -163.365 190.565 -163.035 ;
        RECT 190.235 -164.725 190.565 -164.395 ;
        RECT 190.235 -166.085 190.565 -165.755 ;
        RECT 190.235 -167.445 190.565 -167.115 ;
        RECT 190.235 -168.805 190.565 -168.475 ;
        RECT 190.235 -170.165 190.565 -169.835 ;
        RECT 190.235 -171.525 190.565 -171.195 ;
        RECT 190.235 -172.885 190.565 -172.555 ;
        RECT 190.235 -174.245 190.565 -173.915 ;
        RECT 190.235 -175.605 190.565 -175.275 ;
        RECT 190.235 -176.965 190.565 -176.635 ;
        RECT 190.235 -178.325 190.565 -177.995 ;
        RECT 190.235 -180.57 190.565 -179.44 ;
        RECT 190.24 -180.685 190.56 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 191.595 241.32 191.925 242.45 ;
        RECT 191.595 239.195 191.925 239.525 ;
        RECT 191.595 237.835 191.925 238.165 ;
        RECT 191.6 237.16 191.92 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 191.595 -95.365 191.925 -95.035 ;
        RECT 191.595 -96.725 191.925 -96.395 ;
        RECT 191.595 -98.085 191.925 -97.755 ;
        RECT 191.595 -99.445 191.925 -99.115 ;
        RECT 191.595 -100.805 191.925 -100.475 ;
        RECT 191.595 -102.165 191.925 -101.835 ;
        RECT 191.595 -103.525 191.925 -103.195 ;
        RECT 191.595 -104.885 191.925 -104.555 ;
        RECT 191.595 -106.245 191.925 -105.915 ;
        RECT 191.595 -107.605 191.925 -107.275 ;
        RECT 191.595 -108.965 191.925 -108.635 ;
        RECT 191.595 -110.325 191.925 -109.995 ;
        RECT 191.595 -111.685 191.925 -111.355 ;
        RECT 191.595 -113.045 191.925 -112.715 ;
        RECT 191.595 -114.405 191.925 -114.075 ;
        RECT 191.595 -115.765 191.925 -115.435 ;
        RECT 191.595 -117.125 191.925 -116.795 ;
        RECT 191.595 -118.485 191.925 -118.155 ;
        RECT 191.595 -119.845 191.925 -119.515 ;
        RECT 191.595 -121.205 191.925 -120.875 ;
        RECT 191.595 -122.565 191.925 -122.235 ;
        RECT 191.595 -123.925 191.925 -123.595 ;
        RECT 191.595 -125.285 191.925 -124.955 ;
        RECT 191.595 -126.645 191.925 -126.315 ;
        RECT 191.595 -128.005 191.925 -127.675 ;
        RECT 191.595 -129.365 191.925 -129.035 ;
        RECT 191.595 -130.725 191.925 -130.395 ;
        RECT 191.595 -132.085 191.925 -131.755 ;
        RECT 191.595 -133.445 191.925 -133.115 ;
        RECT 191.595 -134.805 191.925 -134.475 ;
        RECT 191.595 -136.165 191.925 -135.835 ;
        RECT 191.595 -137.525 191.925 -137.195 ;
        RECT 191.595 -138.885 191.925 -138.555 ;
        RECT 191.595 -140.245 191.925 -139.915 ;
        RECT 191.595 -141.605 191.925 -141.275 ;
        RECT 191.595 -142.965 191.925 -142.635 ;
        RECT 191.595 -144.325 191.925 -143.995 ;
        RECT 191.595 -145.685 191.925 -145.355 ;
        RECT 191.595 -147.045 191.925 -146.715 ;
        RECT 191.595 -148.405 191.925 -148.075 ;
        RECT 191.595 -149.765 191.925 -149.435 ;
        RECT 191.595 -151.125 191.925 -150.795 ;
        RECT 191.595 -152.485 191.925 -152.155 ;
        RECT 191.595 -153.845 191.925 -153.515 ;
        RECT 191.595 -155.205 191.925 -154.875 ;
        RECT 191.595 -156.565 191.925 -156.235 ;
        RECT 191.595 -157.925 191.925 -157.595 ;
        RECT 191.595 -159.285 191.925 -158.955 ;
        RECT 191.595 -160.645 191.925 -160.315 ;
        RECT 191.595 -162.005 191.925 -161.675 ;
        RECT 191.595 -163.365 191.925 -163.035 ;
        RECT 191.595 -164.725 191.925 -164.395 ;
        RECT 191.595 -166.085 191.925 -165.755 ;
        RECT 191.595 -167.445 191.925 -167.115 ;
        RECT 191.595 -168.805 191.925 -168.475 ;
        RECT 191.595 -170.165 191.925 -169.835 ;
        RECT 191.595 -171.525 191.925 -171.195 ;
        RECT 191.595 -172.885 191.925 -172.555 ;
        RECT 191.595 -174.245 191.925 -173.915 ;
        RECT 191.595 -175.605 191.925 -175.275 ;
        RECT 191.595 -176.965 191.925 -176.635 ;
        RECT 191.595 -178.325 191.925 -177.995 ;
        RECT 191.595 -180.57 191.925 -179.44 ;
        RECT 191.6 -180.685 191.92 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 192.41 -94.075 192.74 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 192.955 241.32 193.285 242.45 ;
        RECT 192.955 239.195 193.285 239.525 ;
        RECT 192.955 237.835 193.285 238.165 ;
        RECT 192.96 237.16 193.28 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 194.315 241.32 194.645 242.45 ;
        RECT 194.315 239.195 194.645 239.525 ;
        RECT 194.315 237.835 194.645 238.165 ;
        RECT 194.32 237.16 194.64 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 194.315 -1.525 194.645 -1.195 ;
        RECT 194.315 -2.885 194.645 -2.555 ;
        RECT 194.32 -3.56 194.64 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 195.675 241.32 196.005 242.45 ;
        RECT 195.675 239.195 196.005 239.525 ;
        RECT 195.675 237.835 196.005 238.165 ;
        RECT 195.68 237.16 196 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 195.675 -1.525 196.005 -1.195 ;
        RECT 195.675 -2.885 196.005 -2.555 ;
        RECT 195.68 -3.56 196 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 195.675 -91.285 196.005 -90.955 ;
        RECT 195.675 -92.645 196.005 -92.315 ;
        RECT 195.675 -94.005 196.005 -93.675 ;
        RECT 195.675 -95.365 196.005 -95.035 ;
        RECT 195.675 -96.725 196.005 -96.395 ;
        RECT 195.675 -98.085 196.005 -97.755 ;
        RECT 195.675 -99.445 196.005 -99.115 ;
        RECT 195.675 -100.805 196.005 -100.475 ;
        RECT 195.675 -102.165 196.005 -101.835 ;
        RECT 195.675 -103.525 196.005 -103.195 ;
        RECT 195.675 -104.885 196.005 -104.555 ;
        RECT 195.675 -106.245 196.005 -105.915 ;
        RECT 195.675 -107.605 196.005 -107.275 ;
        RECT 195.675 -108.965 196.005 -108.635 ;
        RECT 195.675 -110.325 196.005 -109.995 ;
        RECT 195.675 -111.685 196.005 -111.355 ;
        RECT 195.675 -113.045 196.005 -112.715 ;
        RECT 195.675 -114.405 196.005 -114.075 ;
        RECT 195.675 -115.765 196.005 -115.435 ;
        RECT 195.675 -117.125 196.005 -116.795 ;
        RECT 195.675 -118.485 196.005 -118.155 ;
        RECT 195.675 -119.845 196.005 -119.515 ;
        RECT 195.675 -121.205 196.005 -120.875 ;
        RECT 195.675 -122.565 196.005 -122.235 ;
        RECT 195.675 -123.925 196.005 -123.595 ;
        RECT 195.675 -125.285 196.005 -124.955 ;
        RECT 195.675 -126.645 196.005 -126.315 ;
        RECT 195.675 -128.005 196.005 -127.675 ;
        RECT 195.675 -129.365 196.005 -129.035 ;
        RECT 195.675 -130.725 196.005 -130.395 ;
        RECT 195.675 -132.085 196.005 -131.755 ;
        RECT 195.675 -133.445 196.005 -133.115 ;
        RECT 195.675 -134.805 196.005 -134.475 ;
        RECT 195.675 -136.165 196.005 -135.835 ;
        RECT 195.675 -137.525 196.005 -137.195 ;
        RECT 195.675 -138.885 196.005 -138.555 ;
        RECT 195.675 -140.245 196.005 -139.915 ;
        RECT 195.675 -141.605 196.005 -141.275 ;
        RECT 195.675 -142.965 196.005 -142.635 ;
        RECT 195.675 -144.325 196.005 -143.995 ;
        RECT 195.675 -145.685 196.005 -145.355 ;
        RECT 195.675 -147.045 196.005 -146.715 ;
        RECT 195.675 -148.405 196.005 -148.075 ;
        RECT 195.675 -149.765 196.005 -149.435 ;
        RECT 195.675 -151.125 196.005 -150.795 ;
        RECT 195.675 -152.485 196.005 -152.155 ;
        RECT 195.675 -153.845 196.005 -153.515 ;
        RECT 195.675 -155.205 196.005 -154.875 ;
        RECT 195.675 -156.565 196.005 -156.235 ;
        RECT 195.675 -157.925 196.005 -157.595 ;
        RECT 195.675 -159.285 196.005 -158.955 ;
        RECT 195.675 -160.645 196.005 -160.315 ;
        RECT 195.675 -162.005 196.005 -161.675 ;
        RECT 195.675 -163.365 196.005 -163.035 ;
        RECT 195.675 -164.725 196.005 -164.395 ;
        RECT 195.675 -166.085 196.005 -165.755 ;
        RECT 195.675 -167.445 196.005 -167.115 ;
        RECT 195.675 -168.805 196.005 -168.475 ;
        RECT 195.675 -170.165 196.005 -169.835 ;
        RECT 195.675 -171.525 196.005 -171.195 ;
        RECT 195.675 -172.885 196.005 -172.555 ;
        RECT 195.675 -174.245 196.005 -173.915 ;
        RECT 195.675 -175.605 196.005 -175.275 ;
        RECT 195.675 -176.965 196.005 -176.635 ;
        RECT 195.675 -178.325 196.005 -177.995 ;
        RECT 195.675 -180.57 196.005 -179.44 ;
        RECT 195.68 -180.685 196 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 197.035 241.32 197.365 242.45 ;
        RECT 197.035 239.195 197.365 239.525 ;
        RECT 197.035 237.835 197.365 238.165 ;
        RECT 197.04 237.16 197.36 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 197.035 -1.525 197.365 -1.195 ;
        RECT 197.035 -2.885 197.365 -2.555 ;
        RECT 197.04 -3.56 197.36 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 197.035 -91.285 197.365 -90.955 ;
        RECT 197.035 -92.645 197.365 -92.315 ;
        RECT 197.035 -94.005 197.365 -93.675 ;
        RECT 197.035 -95.365 197.365 -95.035 ;
        RECT 197.035 -96.725 197.365 -96.395 ;
        RECT 197.035 -98.085 197.365 -97.755 ;
        RECT 197.035 -99.445 197.365 -99.115 ;
        RECT 197.035 -100.805 197.365 -100.475 ;
        RECT 197.035 -102.165 197.365 -101.835 ;
        RECT 197.035 -103.525 197.365 -103.195 ;
        RECT 197.035 -104.885 197.365 -104.555 ;
        RECT 197.035 -106.245 197.365 -105.915 ;
        RECT 197.035 -107.605 197.365 -107.275 ;
        RECT 197.035 -108.965 197.365 -108.635 ;
        RECT 197.035 -110.325 197.365 -109.995 ;
        RECT 197.035 -111.685 197.365 -111.355 ;
        RECT 197.035 -113.045 197.365 -112.715 ;
        RECT 197.035 -114.405 197.365 -114.075 ;
        RECT 197.035 -115.765 197.365 -115.435 ;
        RECT 197.035 -117.125 197.365 -116.795 ;
        RECT 197.035 -118.485 197.365 -118.155 ;
        RECT 197.035 -119.845 197.365 -119.515 ;
        RECT 197.035 -121.205 197.365 -120.875 ;
        RECT 197.035 -122.565 197.365 -122.235 ;
        RECT 197.035 -123.925 197.365 -123.595 ;
        RECT 197.035 -125.285 197.365 -124.955 ;
        RECT 197.035 -126.645 197.365 -126.315 ;
        RECT 197.035 -128.005 197.365 -127.675 ;
        RECT 197.035 -129.365 197.365 -129.035 ;
        RECT 197.035 -130.725 197.365 -130.395 ;
        RECT 197.035 -132.085 197.365 -131.755 ;
        RECT 197.035 -133.445 197.365 -133.115 ;
        RECT 197.035 -134.805 197.365 -134.475 ;
        RECT 197.035 -136.165 197.365 -135.835 ;
        RECT 197.035 -137.525 197.365 -137.195 ;
        RECT 197.035 -138.885 197.365 -138.555 ;
        RECT 197.035 -140.245 197.365 -139.915 ;
        RECT 197.035 -141.605 197.365 -141.275 ;
        RECT 197.035 -142.965 197.365 -142.635 ;
        RECT 197.035 -144.325 197.365 -143.995 ;
        RECT 197.035 -145.685 197.365 -145.355 ;
        RECT 197.035 -147.045 197.365 -146.715 ;
        RECT 197.035 -148.405 197.365 -148.075 ;
        RECT 197.035 -149.765 197.365 -149.435 ;
        RECT 197.035 -151.125 197.365 -150.795 ;
        RECT 197.035 -152.485 197.365 -152.155 ;
        RECT 197.035 -153.845 197.365 -153.515 ;
        RECT 197.035 -155.205 197.365 -154.875 ;
        RECT 197.035 -156.565 197.365 -156.235 ;
        RECT 197.035 -157.925 197.365 -157.595 ;
        RECT 197.035 -159.285 197.365 -158.955 ;
        RECT 197.035 -160.645 197.365 -160.315 ;
        RECT 197.035 -162.005 197.365 -161.675 ;
        RECT 197.035 -163.365 197.365 -163.035 ;
        RECT 197.035 -164.725 197.365 -164.395 ;
        RECT 197.035 -166.085 197.365 -165.755 ;
        RECT 197.035 -167.445 197.365 -167.115 ;
        RECT 197.035 -168.805 197.365 -168.475 ;
        RECT 197.035 -170.165 197.365 -169.835 ;
        RECT 197.035 -171.525 197.365 -171.195 ;
        RECT 197.035 -172.885 197.365 -172.555 ;
        RECT 197.035 -174.245 197.365 -173.915 ;
        RECT 197.035 -175.605 197.365 -175.275 ;
        RECT 197.035 -176.965 197.365 -176.635 ;
        RECT 197.035 -178.325 197.365 -177.995 ;
        RECT 197.035 -180.57 197.365 -179.44 ;
        RECT 197.04 -180.685 197.36 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 198.395 241.32 198.725 242.45 ;
        RECT 198.395 239.195 198.725 239.525 ;
        RECT 198.395 237.835 198.725 238.165 ;
        RECT 198.4 237.16 198.72 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 198.395 -95.365 198.725 -95.035 ;
        RECT 198.395 -96.725 198.725 -96.395 ;
        RECT 198.395 -98.085 198.725 -97.755 ;
        RECT 198.395 -99.445 198.725 -99.115 ;
        RECT 198.395 -100.805 198.725 -100.475 ;
        RECT 198.395 -102.165 198.725 -101.835 ;
        RECT 198.395 -103.525 198.725 -103.195 ;
        RECT 198.395 -104.885 198.725 -104.555 ;
        RECT 198.395 -106.245 198.725 -105.915 ;
        RECT 198.395 -107.605 198.725 -107.275 ;
        RECT 198.395 -108.965 198.725 -108.635 ;
        RECT 198.395 -110.325 198.725 -109.995 ;
        RECT 198.395 -111.685 198.725 -111.355 ;
        RECT 198.395 -113.045 198.725 -112.715 ;
        RECT 198.395 -114.405 198.725 -114.075 ;
        RECT 198.395 -115.765 198.725 -115.435 ;
        RECT 198.395 -117.125 198.725 -116.795 ;
        RECT 198.395 -118.485 198.725 -118.155 ;
        RECT 198.395 -119.845 198.725 -119.515 ;
        RECT 198.395 -121.205 198.725 -120.875 ;
        RECT 198.395 -122.565 198.725 -122.235 ;
        RECT 198.395 -123.925 198.725 -123.595 ;
        RECT 198.395 -125.285 198.725 -124.955 ;
        RECT 198.395 -126.645 198.725 -126.315 ;
        RECT 198.395 -128.005 198.725 -127.675 ;
        RECT 198.395 -129.365 198.725 -129.035 ;
        RECT 198.395 -130.725 198.725 -130.395 ;
        RECT 198.395 -132.085 198.725 -131.755 ;
        RECT 198.395 -133.445 198.725 -133.115 ;
        RECT 198.395 -134.805 198.725 -134.475 ;
        RECT 198.395 -136.165 198.725 -135.835 ;
        RECT 198.395 -137.525 198.725 -137.195 ;
        RECT 198.395 -138.885 198.725 -138.555 ;
        RECT 198.395 -140.245 198.725 -139.915 ;
        RECT 198.395 -141.605 198.725 -141.275 ;
        RECT 198.395 -142.965 198.725 -142.635 ;
        RECT 198.395 -144.325 198.725 -143.995 ;
        RECT 198.395 -145.685 198.725 -145.355 ;
        RECT 198.395 -147.045 198.725 -146.715 ;
        RECT 198.395 -148.405 198.725 -148.075 ;
        RECT 198.395 -149.765 198.725 -149.435 ;
        RECT 198.395 -151.125 198.725 -150.795 ;
        RECT 198.395 -152.485 198.725 -152.155 ;
        RECT 198.395 -153.845 198.725 -153.515 ;
        RECT 198.395 -155.205 198.725 -154.875 ;
        RECT 198.395 -156.565 198.725 -156.235 ;
        RECT 198.395 -157.925 198.725 -157.595 ;
        RECT 198.395 -159.285 198.725 -158.955 ;
        RECT 198.395 -160.645 198.725 -160.315 ;
        RECT 198.395 -162.005 198.725 -161.675 ;
        RECT 198.395 -163.365 198.725 -163.035 ;
        RECT 198.395 -164.725 198.725 -164.395 ;
        RECT 198.395 -166.085 198.725 -165.755 ;
        RECT 198.395 -167.445 198.725 -167.115 ;
        RECT 198.395 -168.805 198.725 -168.475 ;
        RECT 198.395 -170.165 198.725 -169.835 ;
        RECT 198.395 -171.525 198.725 -171.195 ;
        RECT 198.395 -172.885 198.725 -172.555 ;
        RECT 198.395 -174.245 198.725 -173.915 ;
        RECT 198.395 -175.605 198.725 -175.275 ;
        RECT 198.395 -176.965 198.725 -176.635 ;
        RECT 198.395 -178.325 198.725 -177.995 ;
        RECT 198.395 -180.57 198.725 -179.44 ;
        RECT 198.4 -180.685 198.72 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 198.51 -94.075 198.84 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 199.755 241.32 200.085 242.45 ;
        RECT 199.755 239.195 200.085 239.525 ;
        RECT 199.755 237.835 200.085 238.165 ;
        RECT 199.76 237.16 200.08 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 199.755 -1.525 200.085 -1.195 ;
        RECT 199.755 -2.885 200.085 -2.555 ;
        RECT 199.76 -3.56 200.08 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 201.115 241.32 201.445 242.45 ;
        RECT 201.115 239.195 201.445 239.525 ;
        RECT 201.115 237.835 201.445 238.165 ;
        RECT 201.12 237.16 201.44 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 201.115 -1.525 201.445 -1.195 ;
        RECT 201.115 -2.885 201.445 -2.555 ;
        RECT 201.12 -3.56 201.44 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 202.475 241.32 202.805 242.45 ;
        RECT 202.475 239.195 202.805 239.525 ;
        RECT 202.475 237.835 202.805 238.165 ;
        RECT 202.48 237.16 202.8 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 202.475 -1.525 202.805 -1.195 ;
        RECT 202.475 -2.885 202.805 -2.555 ;
        RECT 202.48 -3.56 202.8 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 202.475 -91.285 202.805 -90.955 ;
        RECT 202.475 -92.645 202.805 -92.315 ;
        RECT 202.475 -94.005 202.805 -93.675 ;
        RECT 202.475 -95.365 202.805 -95.035 ;
        RECT 202.475 -96.725 202.805 -96.395 ;
        RECT 202.475 -98.085 202.805 -97.755 ;
        RECT 202.475 -99.445 202.805 -99.115 ;
        RECT 202.475 -100.805 202.805 -100.475 ;
        RECT 202.475 -102.165 202.805 -101.835 ;
        RECT 202.475 -103.525 202.805 -103.195 ;
        RECT 202.475 -104.885 202.805 -104.555 ;
        RECT 202.475 -106.245 202.805 -105.915 ;
        RECT 202.475 -107.605 202.805 -107.275 ;
        RECT 202.475 -108.965 202.805 -108.635 ;
        RECT 202.475 -110.325 202.805 -109.995 ;
        RECT 202.475 -111.685 202.805 -111.355 ;
        RECT 202.475 -113.045 202.805 -112.715 ;
        RECT 202.475 -114.405 202.805 -114.075 ;
        RECT 202.475 -115.765 202.805 -115.435 ;
        RECT 202.475 -117.125 202.805 -116.795 ;
        RECT 202.475 -118.485 202.805 -118.155 ;
        RECT 202.475 -119.845 202.805 -119.515 ;
        RECT 202.475 -121.205 202.805 -120.875 ;
        RECT 202.475 -122.565 202.805 -122.235 ;
        RECT 202.475 -123.925 202.805 -123.595 ;
        RECT 202.475 -125.285 202.805 -124.955 ;
        RECT 202.475 -126.645 202.805 -126.315 ;
        RECT 202.475 -128.005 202.805 -127.675 ;
        RECT 202.475 -129.365 202.805 -129.035 ;
        RECT 202.475 -130.725 202.805 -130.395 ;
        RECT 202.475 -132.085 202.805 -131.755 ;
        RECT 202.475 -133.445 202.805 -133.115 ;
        RECT 202.475 -134.805 202.805 -134.475 ;
        RECT 202.475 -136.165 202.805 -135.835 ;
        RECT 202.475 -137.525 202.805 -137.195 ;
        RECT 202.475 -138.885 202.805 -138.555 ;
        RECT 202.475 -140.245 202.805 -139.915 ;
        RECT 202.475 -141.605 202.805 -141.275 ;
        RECT 202.475 -142.965 202.805 -142.635 ;
        RECT 202.475 -144.325 202.805 -143.995 ;
        RECT 202.475 -145.685 202.805 -145.355 ;
        RECT 202.475 -147.045 202.805 -146.715 ;
        RECT 202.475 -148.405 202.805 -148.075 ;
        RECT 202.475 -149.765 202.805 -149.435 ;
        RECT 202.475 -151.125 202.805 -150.795 ;
        RECT 202.475 -152.485 202.805 -152.155 ;
        RECT 202.475 -153.845 202.805 -153.515 ;
        RECT 202.475 -155.205 202.805 -154.875 ;
        RECT 202.475 -156.565 202.805 -156.235 ;
        RECT 202.475 -157.925 202.805 -157.595 ;
        RECT 202.475 -159.285 202.805 -158.955 ;
        RECT 202.475 -160.645 202.805 -160.315 ;
        RECT 202.475 -162.005 202.805 -161.675 ;
        RECT 202.475 -163.365 202.805 -163.035 ;
        RECT 202.475 -164.725 202.805 -164.395 ;
        RECT 202.475 -166.085 202.805 -165.755 ;
        RECT 202.475 -167.445 202.805 -167.115 ;
        RECT 202.475 -168.805 202.805 -168.475 ;
        RECT 202.475 -170.165 202.805 -169.835 ;
        RECT 202.475 -171.525 202.805 -171.195 ;
        RECT 202.475 -172.885 202.805 -172.555 ;
        RECT 202.475 -174.245 202.805 -173.915 ;
        RECT 202.475 -175.605 202.805 -175.275 ;
        RECT 202.475 -176.965 202.805 -176.635 ;
        RECT 202.475 -178.325 202.805 -177.995 ;
        RECT 202.475 -180.57 202.805 -179.44 ;
        RECT 202.48 -180.685 202.8 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 203.835 241.32 204.165 242.45 ;
        RECT 203.835 239.195 204.165 239.525 ;
        RECT 203.835 237.835 204.165 238.165 ;
        RECT 203.84 237.16 204.16 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 203.835 -178.325 204.165 -177.995 ;
        RECT 203.835 -180.57 204.165 -179.44 ;
        RECT 203.84 -180.685 204.16 -95.035 ;
        RECT 203.835 -95.365 204.165 -95.035 ;
        RECT 203.835 -96.725 204.165 -96.395 ;
        RECT 203.835 -98.085 204.165 -97.755 ;
        RECT 203.835 -99.445 204.165 -99.115 ;
        RECT 203.835 -100.805 204.165 -100.475 ;
        RECT 203.835 -102.165 204.165 -101.835 ;
        RECT 203.835 -103.525 204.165 -103.195 ;
        RECT 203.835 -104.885 204.165 -104.555 ;
        RECT 203.835 -106.245 204.165 -105.915 ;
        RECT 203.835 -107.605 204.165 -107.275 ;
        RECT 203.835 -108.965 204.165 -108.635 ;
        RECT 203.835 -110.325 204.165 -109.995 ;
        RECT 203.835 -111.685 204.165 -111.355 ;
        RECT 203.835 -113.045 204.165 -112.715 ;
        RECT 203.835 -114.405 204.165 -114.075 ;
        RECT 203.835 -115.765 204.165 -115.435 ;
        RECT 203.835 -117.125 204.165 -116.795 ;
        RECT 203.835 -118.485 204.165 -118.155 ;
        RECT 203.835 -119.845 204.165 -119.515 ;
        RECT 203.835 -121.205 204.165 -120.875 ;
        RECT 203.835 -122.565 204.165 -122.235 ;
        RECT 203.835 -123.925 204.165 -123.595 ;
        RECT 203.835 -125.285 204.165 -124.955 ;
        RECT 203.835 -126.645 204.165 -126.315 ;
        RECT 203.835 -128.005 204.165 -127.675 ;
        RECT 203.835 -129.365 204.165 -129.035 ;
        RECT 203.835 -130.725 204.165 -130.395 ;
        RECT 203.835 -132.085 204.165 -131.755 ;
        RECT 203.835 -133.445 204.165 -133.115 ;
        RECT 203.835 -134.805 204.165 -134.475 ;
        RECT 203.835 -136.165 204.165 -135.835 ;
        RECT 203.835 -137.525 204.165 -137.195 ;
        RECT 203.835 -138.885 204.165 -138.555 ;
        RECT 203.835 -140.245 204.165 -139.915 ;
        RECT 203.835 -141.605 204.165 -141.275 ;
        RECT 203.835 -142.965 204.165 -142.635 ;
        RECT 203.835 -144.325 204.165 -143.995 ;
        RECT 203.835 -145.685 204.165 -145.355 ;
        RECT 203.835 -147.045 204.165 -146.715 ;
        RECT 203.835 -148.405 204.165 -148.075 ;
        RECT 203.835 -149.765 204.165 -149.435 ;
        RECT 203.835 -151.125 204.165 -150.795 ;
        RECT 203.835 -152.485 204.165 -152.155 ;
        RECT 203.835 -153.845 204.165 -153.515 ;
        RECT 203.835 -155.205 204.165 -154.875 ;
        RECT 203.835 -156.565 204.165 -156.235 ;
        RECT 203.835 -157.925 204.165 -157.595 ;
        RECT 203.835 -159.285 204.165 -158.955 ;
        RECT 203.835 -160.645 204.165 -160.315 ;
        RECT 203.835 -162.005 204.165 -161.675 ;
        RECT 203.835 -163.365 204.165 -163.035 ;
        RECT 203.835 -164.725 204.165 -164.395 ;
        RECT 203.835 -166.085 204.165 -165.755 ;
        RECT 203.835 -167.445 204.165 -167.115 ;
        RECT 203.835 -168.805 204.165 -168.475 ;
        RECT 203.835 -170.165 204.165 -169.835 ;
        RECT 203.835 -171.525 204.165 -171.195 ;
        RECT 203.835 -172.885 204.165 -172.555 ;
        RECT 203.835 -174.245 204.165 -173.915 ;
        RECT 203.835 -175.605 204.165 -175.275 ;
        RECT 203.835 -176.965 204.165 -176.635 ;
    END
    PORT
      LAYER met3 ;
        RECT 137.51 -94.075 137.84 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 138.555 241.32 138.885 242.45 ;
        RECT 138.555 239.195 138.885 239.525 ;
        RECT 138.555 237.835 138.885 238.165 ;
        RECT 138.56 237.16 138.88 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 138.555 -1.525 138.885 -1.195 ;
        RECT 138.555 -2.885 138.885 -2.555 ;
        RECT 138.56 -3.56 138.88 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 139.915 241.32 140.245 242.45 ;
        RECT 139.915 239.195 140.245 239.525 ;
        RECT 139.915 237.835 140.245 238.165 ;
        RECT 139.92 237.16 140.24 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 139.915 -1.525 140.245 -1.195 ;
        RECT 139.915 -2.885 140.245 -2.555 ;
        RECT 139.92 -3.56 140.24 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 141.275 241.32 141.605 242.45 ;
        RECT 141.275 239.195 141.605 239.525 ;
        RECT 141.275 237.835 141.605 238.165 ;
        RECT 141.28 237.16 141.6 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 141.275 -1.525 141.605 -1.195 ;
        RECT 141.275 -2.885 141.605 -2.555 ;
        RECT 141.28 -3.56 141.6 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 141.275 -91.285 141.605 -90.955 ;
        RECT 141.275 -92.645 141.605 -92.315 ;
        RECT 141.275 -94.005 141.605 -93.675 ;
        RECT 141.275 -95.365 141.605 -95.035 ;
        RECT 141.275 -96.725 141.605 -96.395 ;
        RECT 141.275 -98.085 141.605 -97.755 ;
        RECT 141.275 -99.445 141.605 -99.115 ;
        RECT 141.275 -100.805 141.605 -100.475 ;
        RECT 141.275 -102.165 141.605 -101.835 ;
        RECT 141.275 -103.525 141.605 -103.195 ;
        RECT 141.275 -104.885 141.605 -104.555 ;
        RECT 141.275 -106.245 141.605 -105.915 ;
        RECT 141.275 -107.605 141.605 -107.275 ;
        RECT 141.275 -108.965 141.605 -108.635 ;
        RECT 141.275 -110.325 141.605 -109.995 ;
        RECT 141.275 -111.685 141.605 -111.355 ;
        RECT 141.275 -113.045 141.605 -112.715 ;
        RECT 141.275 -114.405 141.605 -114.075 ;
        RECT 141.275 -115.765 141.605 -115.435 ;
        RECT 141.275 -117.125 141.605 -116.795 ;
        RECT 141.275 -118.485 141.605 -118.155 ;
        RECT 141.275 -119.845 141.605 -119.515 ;
        RECT 141.275 -121.205 141.605 -120.875 ;
        RECT 141.275 -122.565 141.605 -122.235 ;
        RECT 141.275 -123.925 141.605 -123.595 ;
        RECT 141.275 -125.285 141.605 -124.955 ;
        RECT 141.275 -126.645 141.605 -126.315 ;
        RECT 141.275 -128.005 141.605 -127.675 ;
        RECT 141.275 -129.365 141.605 -129.035 ;
        RECT 141.275 -130.725 141.605 -130.395 ;
        RECT 141.275 -132.085 141.605 -131.755 ;
        RECT 141.275 -133.445 141.605 -133.115 ;
        RECT 141.275 -134.805 141.605 -134.475 ;
        RECT 141.275 -136.165 141.605 -135.835 ;
        RECT 141.275 -137.525 141.605 -137.195 ;
        RECT 141.275 -138.885 141.605 -138.555 ;
        RECT 141.275 -140.245 141.605 -139.915 ;
        RECT 141.275 -141.605 141.605 -141.275 ;
        RECT 141.275 -142.965 141.605 -142.635 ;
        RECT 141.275 -144.325 141.605 -143.995 ;
        RECT 141.275 -145.685 141.605 -145.355 ;
        RECT 141.275 -147.045 141.605 -146.715 ;
        RECT 141.275 -148.405 141.605 -148.075 ;
        RECT 141.275 -149.765 141.605 -149.435 ;
        RECT 141.275 -151.125 141.605 -150.795 ;
        RECT 141.275 -152.485 141.605 -152.155 ;
        RECT 141.275 -153.845 141.605 -153.515 ;
        RECT 141.275 -155.205 141.605 -154.875 ;
        RECT 141.275 -156.565 141.605 -156.235 ;
        RECT 141.275 -157.925 141.605 -157.595 ;
        RECT 141.275 -159.285 141.605 -158.955 ;
        RECT 141.275 -160.645 141.605 -160.315 ;
        RECT 141.275 -162.005 141.605 -161.675 ;
        RECT 141.275 -163.365 141.605 -163.035 ;
        RECT 141.275 -164.725 141.605 -164.395 ;
        RECT 141.275 -166.085 141.605 -165.755 ;
        RECT 141.275 -167.445 141.605 -167.115 ;
        RECT 141.275 -168.805 141.605 -168.475 ;
        RECT 141.275 -170.165 141.605 -169.835 ;
        RECT 141.275 -171.525 141.605 -171.195 ;
        RECT 141.275 -172.885 141.605 -172.555 ;
        RECT 141.275 -174.245 141.605 -173.915 ;
        RECT 141.275 -175.605 141.605 -175.275 ;
        RECT 141.275 -176.965 141.605 -176.635 ;
        RECT 141.275 -178.325 141.605 -177.995 ;
        RECT 141.275 -180.57 141.605 -179.44 ;
        RECT 141.28 -180.685 141.6 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 142.635 241.32 142.965 242.45 ;
        RECT 142.635 239.195 142.965 239.525 ;
        RECT 142.635 237.835 142.965 238.165 ;
        RECT 142.64 237.16 142.96 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 142.635 -95.365 142.965 -95.035 ;
        RECT 142.635 -96.725 142.965 -96.395 ;
        RECT 142.635 -98.085 142.965 -97.755 ;
        RECT 142.635 -99.445 142.965 -99.115 ;
        RECT 142.635 -100.805 142.965 -100.475 ;
        RECT 142.635 -102.165 142.965 -101.835 ;
        RECT 142.635 -103.525 142.965 -103.195 ;
        RECT 142.635 -104.885 142.965 -104.555 ;
        RECT 142.635 -106.245 142.965 -105.915 ;
        RECT 142.635 -107.605 142.965 -107.275 ;
        RECT 142.635 -108.965 142.965 -108.635 ;
        RECT 142.635 -110.325 142.965 -109.995 ;
        RECT 142.635 -111.685 142.965 -111.355 ;
        RECT 142.635 -113.045 142.965 -112.715 ;
        RECT 142.635 -114.405 142.965 -114.075 ;
        RECT 142.635 -115.765 142.965 -115.435 ;
        RECT 142.635 -117.125 142.965 -116.795 ;
        RECT 142.635 -118.485 142.965 -118.155 ;
        RECT 142.635 -119.845 142.965 -119.515 ;
        RECT 142.635 -121.205 142.965 -120.875 ;
        RECT 142.635 -122.565 142.965 -122.235 ;
        RECT 142.635 -123.925 142.965 -123.595 ;
        RECT 142.635 -125.285 142.965 -124.955 ;
        RECT 142.635 -126.645 142.965 -126.315 ;
        RECT 142.635 -128.005 142.965 -127.675 ;
        RECT 142.635 -129.365 142.965 -129.035 ;
        RECT 142.635 -130.725 142.965 -130.395 ;
        RECT 142.635 -132.085 142.965 -131.755 ;
        RECT 142.635 -133.445 142.965 -133.115 ;
        RECT 142.635 -134.805 142.965 -134.475 ;
        RECT 142.635 -136.165 142.965 -135.835 ;
        RECT 142.635 -137.525 142.965 -137.195 ;
        RECT 142.635 -138.885 142.965 -138.555 ;
        RECT 142.635 -140.245 142.965 -139.915 ;
        RECT 142.635 -141.605 142.965 -141.275 ;
        RECT 142.635 -142.965 142.965 -142.635 ;
        RECT 142.635 -144.325 142.965 -143.995 ;
        RECT 142.635 -145.685 142.965 -145.355 ;
        RECT 142.635 -147.045 142.965 -146.715 ;
        RECT 142.635 -148.405 142.965 -148.075 ;
        RECT 142.635 -149.765 142.965 -149.435 ;
        RECT 142.635 -151.125 142.965 -150.795 ;
        RECT 142.635 -152.485 142.965 -152.155 ;
        RECT 142.635 -153.845 142.965 -153.515 ;
        RECT 142.635 -155.205 142.965 -154.875 ;
        RECT 142.635 -156.565 142.965 -156.235 ;
        RECT 142.635 -157.925 142.965 -157.595 ;
        RECT 142.635 -159.285 142.965 -158.955 ;
        RECT 142.635 -160.645 142.965 -160.315 ;
        RECT 142.635 -162.005 142.965 -161.675 ;
        RECT 142.635 -163.365 142.965 -163.035 ;
        RECT 142.635 -164.725 142.965 -164.395 ;
        RECT 142.635 -166.085 142.965 -165.755 ;
        RECT 142.635 -167.445 142.965 -167.115 ;
        RECT 142.635 -168.805 142.965 -168.475 ;
        RECT 142.635 -170.165 142.965 -169.835 ;
        RECT 142.635 -171.525 142.965 -171.195 ;
        RECT 142.635 -172.885 142.965 -172.555 ;
        RECT 142.635 -174.245 142.965 -173.915 ;
        RECT 142.635 -175.605 142.965 -175.275 ;
        RECT 142.635 -176.965 142.965 -176.635 ;
        RECT 142.635 -178.325 142.965 -177.995 ;
        RECT 142.635 -180.57 142.965 -179.44 ;
        RECT 142.64 -180.685 142.96 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 143.61 -94.075 143.94 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 143.995 241.32 144.325 242.45 ;
        RECT 143.995 239.195 144.325 239.525 ;
        RECT 143.995 237.835 144.325 238.165 ;
        RECT 144 237.16 144.32 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 145.355 241.32 145.685 242.45 ;
        RECT 145.355 239.195 145.685 239.525 ;
        RECT 145.355 237.835 145.685 238.165 ;
        RECT 145.36 237.16 145.68 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 145.355 -1.525 145.685 -1.195 ;
        RECT 145.355 -2.885 145.685 -2.555 ;
        RECT 145.36 -3.56 145.68 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 146.715 241.32 147.045 242.45 ;
        RECT 146.715 239.195 147.045 239.525 ;
        RECT 146.715 237.835 147.045 238.165 ;
        RECT 146.72 237.16 147.04 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 146.715 -1.525 147.045 -1.195 ;
        RECT 146.715 -2.885 147.045 -2.555 ;
        RECT 146.72 -3.56 147.04 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 146.715 -91.285 147.045 -90.955 ;
        RECT 146.715 -92.645 147.045 -92.315 ;
        RECT 146.715 -94.005 147.045 -93.675 ;
        RECT 146.715 -95.365 147.045 -95.035 ;
        RECT 146.715 -96.725 147.045 -96.395 ;
        RECT 146.715 -98.085 147.045 -97.755 ;
        RECT 146.715 -99.445 147.045 -99.115 ;
        RECT 146.715 -100.805 147.045 -100.475 ;
        RECT 146.715 -102.165 147.045 -101.835 ;
        RECT 146.715 -103.525 147.045 -103.195 ;
        RECT 146.715 -104.885 147.045 -104.555 ;
        RECT 146.715 -106.245 147.045 -105.915 ;
        RECT 146.715 -107.605 147.045 -107.275 ;
        RECT 146.715 -108.965 147.045 -108.635 ;
        RECT 146.715 -110.325 147.045 -109.995 ;
        RECT 146.715 -111.685 147.045 -111.355 ;
        RECT 146.715 -113.045 147.045 -112.715 ;
        RECT 146.715 -114.405 147.045 -114.075 ;
        RECT 146.715 -115.765 147.045 -115.435 ;
        RECT 146.715 -117.125 147.045 -116.795 ;
        RECT 146.715 -118.485 147.045 -118.155 ;
        RECT 146.715 -119.845 147.045 -119.515 ;
        RECT 146.715 -121.205 147.045 -120.875 ;
        RECT 146.715 -122.565 147.045 -122.235 ;
        RECT 146.715 -123.925 147.045 -123.595 ;
        RECT 146.715 -125.285 147.045 -124.955 ;
        RECT 146.715 -126.645 147.045 -126.315 ;
        RECT 146.715 -128.005 147.045 -127.675 ;
        RECT 146.715 -129.365 147.045 -129.035 ;
        RECT 146.715 -130.725 147.045 -130.395 ;
        RECT 146.715 -132.085 147.045 -131.755 ;
        RECT 146.715 -133.445 147.045 -133.115 ;
        RECT 146.715 -134.805 147.045 -134.475 ;
        RECT 146.715 -136.165 147.045 -135.835 ;
        RECT 146.715 -137.525 147.045 -137.195 ;
        RECT 146.715 -138.885 147.045 -138.555 ;
        RECT 146.715 -140.245 147.045 -139.915 ;
        RECT 146.715 -141.605 147.045 -141.275 ;
        RECT 146.715 -142.965 147.045 -142.635 ;
        RECT 146.715 -144.325 147.045 -143.995 ;
        RECT 146.715 -145.685 147.045 -145.355 ;
        RECT 146.715 -147.045 147.045 -146.715 ;
        RECT 146.715 -148.405 147.045 -148.075 ;
        RECT 146.715 -149.765 147.045 -149.435 ;
        RECT 146.715 -151.125 147.045 -150.795 ;
        RECT 146.715 -152.485 147.045 -152.155 ;
        RECT 146.715 -153.845 147.045 -153.515 ;
        RECT 146.715 -155.205 147.045 -154.875 ;
        RECT 146.715 -156.565 147.045 -156.235 ;
        RECT 146.715 -157.925 147.045 -157.595 ;
        RECT 146.715 -159.285 147.045 -158.955 ;
        RECT 146.715 -160.645 147.045 -160.315 ;
        RECT 146.715 -162.005 147.045 -161.675 ;
        RECT 146.715 -163.365 147.045 -163.035 ;
        RECT 146.715 -164.725 147.045 -164.395 ;
        RECT 146.715 -166.085 147.045 -165.755 ;
        RECT 146.715 -167.445 147.045 -167.115 ;
        RECT 146.715 -168.805 147.045 -168.475 ;
        RECT 146.715 -170.165 147.045 -169.835 ;
        RECT 146.715 -171.525 147.045 -171.195 ;
        RECT 146.715 -172.885 147.045 -172.555 ;
        RECT 146.715 -174.245 147.045 -173.915 ;
        RECT 146.715 -175.605 147.045 -175.275 ;
        RECT 146.715 -176.965 147.045 -176.635 ;
        RECT 146.715 -178.325 147.045 -177.995 ;
        RECT 146.715 -180.57 147.045 -179.44 ;
        RECT 146.72 -180.685 147.04 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 148.075 241.32 148.405 242.45 ;
        RECT 148.075 239.195 148.405 239.525 ;
        RECT 148.075 237.835 148.405 238.165 ;
        RECT 148.08 237.16 148.4 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 148.075 -1.525 148.405 -1.195 ;
        RECT 148.075 -2.885 148.405 -2.555 ;
        RECT 148.08 -3.56 148.4 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 148.075 -91.285 148.405 -90.955 ;
        RECT 148.075 -92.645 148.405 -92.315 ;
        RECT 148.075 -94.005 148.405 -93.675 ;
        RECT 148.075 -95.365 148.405 -95.035 ;
        RECT 148.075 -96.725 148.405 -96.395 ;
        RECT 148.075 -98.085 148.405 -97.755 ;
        RECT 148.075 -99.445 148.405 -99.115 ;
        RECT 148.075 -100.805 148.405 -100.475 ;
        RECT 148.075 -102.165 148.405 -101.835 ;
        RECT 148.075 -103.525 148.405 -103.195 ;
        RECT 148.075 -104.885 148.405 -104.555 ;
        RECT 148.075 -106.245 148.405 -105.915 ;
        RECT 148.075 -107.605 148.405 -107.275 ;
        RECT 148.075 -108.965 148.405 -108.635 ;
        RECT 148.075 -110.325 148.405 -109.995 ;
        RECT 148.075 -111.685 148.405 -111.355 ;
        RECT 148.075 -113.045 148.405 -112.715 ;
        RECT 148.075 -114.405 148.405 -114.075 ;
        RECT 148.075 -115.765 148.405 -115.435 ;
        RECT 148.075 -117.125 148.405 -116.795 ;
        RECT 148.075 -118.485 148.405 -118.155 ;
        RECT 148.075 -119.845 148.405 -119.515 ;
        RECT 148.075 -121.205 148.405 -120.875 ;
        RECT 148.075 -122.565 148.405 -122.235 ;
        RECT 148.075 -123.925 148.405 -123.595 ;
        RECT 148.075 -125.285 148.405 -124.955 ;
        RECT 148.075 -126.645 148.405 -126.315 ;
        RECT 148.075 -128.005 148.405 -127.675 ;
        RECT 148.075 -129.365 148.405 -129.035 ;
        RECT 148.075 -130.725 148.405 -130.395 ;
        RECT 148.075 -132.085 148.405 -131.755 ;
        RECT 148.075 -133.445 148.405 -133.115 ;
        RECT 148.075 -134.805 148.405 -134.475 ;
        RECT 148.075 -136.165 148.405 -135.835 ;
        RECT 148.075 -137.525 148.405 -137.195 ;
        RECT 148.075 -138.885 148.405 -138.555 ;
        RECT 148.075 -140.245 148.405 -139.915 ;
        RECT 148.075 -141.605 148.405 -141.275 ;
        RECT 148.075 -142.965 148.405 -142.635 ;
        RECT 148.075 -144.325 148.405 -143.995 ;
        RECT 148.075 -145.685 148.405 -145.355 ;
        RECT 148.075 -147.045 148.405 -146.715 ;
        RECT 148.075 -148.405 148.405 -148.075 ;
        RECT 148.075 -149.765 148.405 -149.435 ;
        RECT 148.075 -151.125 148.405 -150.795 ;
        RECT 148.075 -152.485 148.405 -152.155 ;
        RECT 148.075 -153.845 148.405 -153.515 ;
        RECT 148.075 -155.205 148.405 -154.875 ;
        RECT 148.075 -156.565 148.405 -156.235 ;
        RECT 148.075 -157.925 148.405 -157.595 ;
        RECT 148.075 -159.285 148.405 -158.955 ;
        RECT 148.075 -160.645 148.405 -160.315 ;
        RECT 148.075 -162.005 148.405 -161.675 ;
        RECT 148.075 -163.365 148.405 -163.035 ;
        RECT 148.075 -164.725 148.405 -164.395 ;
        RECT 148.075 -166.085 148.405 -165.755 ;
        RECT 148.075 -167.445 148.405 -167.115 ;
        RECT 148.075 -168.805 148.405 -168.475 ;
        RECT 148.075 -170.165 148.405 -169.835 ;
        RECT 148.075 -171.525 148.405 -171.195 ;
        RECT 148.075 -172.885 148.405 -172.555 ;
        RECT 148.075 -174.245 148.405 -173.915 ;
        RECT 148.075 -175.605 148.405 -175.275 ;
        RECT 148.075 -176.965 148.405 -176.635 ;
        RECT 148.075 -178.325 148.405 -177.995 ;
        RECT 148.075 -180.57 148.405 -179.44 ;
        RECT 148.08 -180.685 148.4 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 149.435 241.32 149.765 242.45 ;
        RECT 149.435 239.195 149.765 239.525 ;
        RECT 149.435 237.835 149.765 238.165 ;
        RECT 149.44 237.16 149.76 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 149.435 -95.365 149.765 -95.035 ;
        RECT 149.435 -96.725 149.765 -96.395 ;
        RECT 149.435 -98.085 149.765 -97.755 ;
        RECT 149.435 -99.445 149.765 -99.115 ;
        RECT 149.435 -100.805 149.765 -100.475 ;
        RECT 149.435 -102.165 149.765 -101.835 ;
        RECT 149.435 -103.525 149.765 -103.195 ;
        RECT 149.435 -104.885 149.765 -104.555 ;
        RECT 149.435 -106.245 149.765 -105.915 ;
        RECT 149.435 -107.605 149.765 -107.275 ;
        RECT 149.435 -108.965 149.765 -108.635 ;
        RECT 149.435 -110.325 149.765 -109.995 ;
        RECT 149.435 -111.685 149.765 -111.355 ;
        RECT 149.435 -113.045 149.765 -112.715 ;
        RECT 149.435 -114.405 149.765 -114.075 ;
        RECT 149.435 -115.765 149.765 -115.435 ;
        RECT 149.435 -117.125 149.765 -116.795 ;
        RECT 149.435 -118.485 149.765 -118.155 ;
        RECT 149.435 -119.845 149.765 -119.515 ;
        RECT 149.435 -121.205 149.765 -120.875 ;
        RECT 149.435 -122.565 149.765 -122.235 ;
        RECT 149.435 -123.925 149.765 -123.595 ;
        RECT 149.435 -125.285 149.765 -124.955 ;
        RECT 149.435 -126.645 149.765 -126.315 ;
        RECT 149.435 -128.005 149.765 -127.675 ;
        RECT 149.435 -129.365 149.765 -129.035 ;
        RECT 149.435 -130.725 149.765 -130.395 ;
        RECT 149.435 -132.085 149.765 -131.755 ;
        RECT 149.435 -133.445 149.765 -133.115 ;
        RECT 149.435 -134.805 149.765 -134.475 ;
        RECT 149.435 -136.165 149.765 -135.835 ;
        RECT 149.435 -137.525 149.765 -137.195 ;
        RECT 149.435 -138.885 149.765 -138.555 ;
        RECT 149.435 -140.245 149.765 -139.915 ;
        RECT 149.435 -141.605 149.765 -141.275 ;
        RECT 149.435 -142.965 149.765 -142.635 ;
        RECT 149.435 -144.325 149.765 -143.995 ;
        RECT 149.435 -145.685 149.765 -145.355 ;
        RECT 149.435 -147.045 149.765 -146.715 ;
        RECT 149.435 -148.405 149.765 -148.075 ;
        RECT 149.435 -149.765 149.765 -149.435 ;
        RECT 149.435 -151.125 149.765 -150.795 ;
        RECT 149.435 -152.485 149.765 -152.155 ;
        RECT 149.435 -153.845 149.765 -153.515 ;
        RECT 149.435 -155.205 149.765 -154.875 ;
        RECT 149.435 -156.565 149.765 -156.235 ;
        RECT 149.435 -157.925 149.765 -157.595 ;
        RECT 149.435 -159.285 149.765 -158.955 ;
        RECT 149.435 -160.645 149.765 -160.315 ;
        RECT 149.435 -162.005 149.765 -161.675 ;
        RECT 149.435 -163.365 149.765 -163.035 ;
        RECT 149.435 -164.725 149.765 -164.395 ;
        RECT 149.435 -166.085 149.765 -165.755 ;
        RECT 149.435 -167.445 149.765 -167.115 ;
        RECT 149.435 -168.805 149.765 -168.475 ;
        RECT 149.435 -170.165 149.765 -169.835 ;
        RECT 149.435 -171.525 149.765 -171.195 ;
        RECT 149.435 -172.885 149.765 -172.555 ;
        RECT 149.435 -174.245 149.765 -173.915 ;
        RECT 149.435 -175.605 149.765 -175.275 ;
        RECT 149.435 -176.965 149.765 -176.635 ;
        RECT 149.435 -178.325 149.765 -177.995 ;
        RECT 149.435 -180.57 149.765 -179.44 ;
        RECT 149.44 -180.685 149.76 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 149.71 -94.075 150.04 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 150.795 241.32 151.125 242.45 ;
        RECT 150.795 239.195 151.125 239.525 ;
        RECT 150.795 237.835 151.125 238.165 ;
        RECT 150.8 237.16 151.12 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 150.795 -1.525 151.125 -1.195 ;
        RECT 150.795 -2.885 151.125 -2.555 ;
        RECT 150.8 -3.56 151.12 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 152.155 241.32 152.485 242.45 ;
        RECT 152.155 239.195 152.485 239.525 ;
        RECT 152.155 237.835 152.485 238.165 ;
        RECT 152.16 237.16 152.48 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 152.155 -1.525 152.485 -1.195 ;
        RECT 152.155 -2.885 152.485 -2.555 ;
        RECT 152.16 -3.56 152.48 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 153.515 241.32 153.845 242.45 ;
        RECT 153.515 239.195 153.845 239.525 ;
        RECT 153.515 237.835 153.845 238.165 ;
        RECT 153.52 237.16 153.84 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 153.515 -1.525 153.845 -1.195 ;
        RECT 153.515 -2.885 153.845 -2.555 ;
        RECT 153.52 -3.56 153.84 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 154.875 241.32 155.205 242.45 ;
        RECT 154.875 239.195 155.205 239.525 ;
        RECT 154.875 237.835 155.205 238.165 ;
        RECT 154.88 237.16 155.2 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 154.875 -95.365 155.205 -95.035 ;
        RECT 154.875 -96.725 155.205 -96.395 ;
        RECT 154.875 -98.085 155.205 -97.755 ;
        RECT 154.875 -99.445 155.205 -99.115 ;
        RECT 154.875 -100.805 155.205 -100.475 ;
        RECT 154.875 -102.165 155.205 -101.835 ;
        RECT 154.875 -103.525 155.205 -103.195 ;
        RECT 154.875 -104.885 155.205 -104.555 ;
        RECT 154.875 -106.245 155.205 -105.915 ;
        RECT 154.875 -107.605 155.205 -107.275 ;
        RECT 154.875 -108.965 155.205 -108.635 ;
        RECT 154.875 -110.325 155.205 -109.995 ;
        RECT 154.875 -111.685 155.205 -111.355 ;
        RECT 154.875 -113.045 155.205 -112.715 ;
        RECT 154.875 -114.405 155.205 -114.075 ;
        RECT 154.875 -115.765 155.205 -115.435 ;
        RECT 154.875 -117.125 155.205 -116.795 ;
        RECT 154.875 -118.485 155.205 -118.155 ;
        RECT 154.875 -119.845 155.205 -119.515 ;
        RECT 154.875 -121.205 155.205 -120.875 ;
        RECT 154.875 -122.565 155.205 -122.235 ;
        RECT 154.875 -123.925 155.205 -123.595 ;
        RECT 154.875 -125.285 155.205 -124.955 ;
        RECT 154.875 -126.645 155.205 -126.315 ;
        RECT 154.875 -128.005 155.205 -127.675 ;
        RECT 154.875 -129.365 155.205 -129.035 ;
        RECT 154.875 -130.725 155.205 -130.395 ;
        RECT 154.875 -132.085 155.205 -131.755 ;
        RECT 154.875 -133.445 155.205 -133.115 ;
        RECT 154.875 -134.805 155.205 -134.475 ;
        RECT 154.875 -136.165 155.205 -135.835 ;
        RECT 154.875 -137.525 155.205 -137.195 ;
        RECT 154.875 -138.885 155.205 -138.555 ;
        RECT 154.875 -140.245 155.205 -139.915 ;
        RECT 154.875 -141.605 155.205 -141.275 ;
        RECT 154.875 -142.965 155.205 -142.635 ;
        RECT 154.875 -144.325 155.205 -143.995 ;
        RECT 154.875 -145.685 155.205 -145.355 ;
        RECT 154.875 -147.045 155.205 -146.715 ;
        RECT 154.875 -148.405 155.205 -148.075 ;
        RECT 154.875 -149.765 155.205 -149.435 ;
        RECT 154.875 -151.125 155.205 -150.795 ;
        RECT 154.875 -152.485 155.205 -152.155 ;
        RECT 154.875 -153.845 155.205 -153.515 ;
        RECT 154.875 -155.205 155.205 -154.875 ;
        RECT 154.875 -156.565 155.205 -156.235 ;
        RECT 154.875 -157.925 155.205 -157.595 ;
        RECT 154.875 -159.285 155.205 -158.955 ;
        RECT 154.875 -160.645 155.205 -160.315 ;
        RECT 154.875 -162.005 155.205 -161.675 ;
        RECT 154.875 -163.365 155.205 -163.035 ;
        RECT 154.875 -164.725 155.205 -164.395 ;
        RECT 154.875 -166.085 155.205 -165.755 ;
        RECT 154.875 -167.445 155.205 -167.115 ;
        RECT 154.875 -168.805 155.205 -168.475 ;
        RECT 154.875 -170.165 155.205 -169.835 ;
        RECT 154.875 -171.525 155.205 -171.195 ;
        RECT 154.875 -172.885 155.205 -172.555 ;
        RECT 154.875 -174.245 155.205 -173.915 ;
        RECT 154.875 -175.605 155.205 -175.275 ;
        RECT 154.875 -176.965 155.205 -176.635 ;
        RECT 154.875 -178.325 155.205 -177.995 ;
        RECT 154.875 -180.57 155.205 -179.44 ;
        RECT 154.88 -180.685 155.2 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 155.81 -94.075 156.14 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 156.235 241.32 156.565 242.45 ;
        RECT 156.235 239.195 156.565 239.525 ;
        RECT 156.235 237.835 156.565 238.165 ;
        RECT 156.24 237.16 156.56 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 157.595 241.32 157.925 242.45 ;
        RECT 157.595 239.195 157.925 239.525 ;
        RECT 157.595 237.835 157.925 238.165 ;
        RECT 157.6 237.16 157.92 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 157.595 -1.525 157.925 -1.195 ;
        RECT 157.595 -2.885 157.925 -2.555 ;
        RECT 157.6 -3.56 157.92 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 158.955 241.32 159.285 242.45 ;
        RECT 158.955 239.195 159.285 239.525 ;
        RECT 158.955 237.835 159.285 238.165 ;
        RECT 158.96 237.16 159.28 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 158.955 -1.525 159.285 -1.195 ;
        RECT 158.955 -2.885 159.285 -2.555 ;
        RECT 158.96 -3.56 159.28 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 158.955 -91.285 159.285 -90.955 ;
        RECT 158.955 -92.645 159.285 -92.315 ;
        RECT 158.955 -94.005 159.285 -93.675 ;
        RECT 158.955 -95.365 159.285 -95.035 ;
        RECT 158.955 -96.725 159.285 -96.395 ;
        RECT 158.955 -98.085 159.285 -97.755 ;
        RECT 158.955 -99.445 159.285 -99.115 ;
        RECT 158.955 -100.805 159.285 -100.475 ;
        RECT 158.955 -102.165 159.285 -101.835 ;
        RECT 158.955 -103.525 159.285 -103.195 ;
        RECT 158.955 -104.885 159.285 -104.555 ;
        RECT 158.955 -106.245 159.285 -105.915 ;
        RECT 158.955 -107.605 159.285 -107.275 ;
        RECT 158.955 -108.965 159.285 -108.635 ;
        RECT 158.955 -110.325 159.285 -109.995 ;
        RECT 158.955 -111.685 159.285 -111.355 ;
        RECT 158.955 -113.045 159.285 -112.715 ;
        RECT 158.955 -114.405 159.285 -114.075 ;
        RECT 158.955 -115.765 159.285 -115.435 ;
        RECT 158.955 -117.125 159.285 -116.795 ;
        RECT 158.955 -118.485 159.285 -118.155 ;
        RECT 158.955 -119.845 159.285 -119.515 ;
        RECT 158.955 -121.205 159.285 -120.875 ;
        RECT 158.955 -122.565 159.285 -122.235 ;
        RECT 158.955 -123.925 159.285 -123.595 ;
        RECT 158.955 -125.285 159.285 -124.955 ;
        RECT 158.955 -126.645 159.285 -126.315 ;
        RECT 158.955 -128.005 159.285 -127.675 ;
        RECT 158.955 -129.365 159.285 -129.035 ;
        RECT 158.955 -130.725 159.285 -130.395 ;
        RECT 158.955 -132.085 159.285 -131.755 ;
        RECT 158.955 -133.445 159.285 -133.115 ;
        RECT 158.955 -134.805 159.285 -134.475 ;
        RECT 158.955 -136.165 159.285 -135.835 ;
        RECT 158.955 -137.525 159.285 -137.195 ;
        RECT 158.955 -138.885 159.285 -138.555 ;
        RECT 158.955 -140.245 159.285 -139.915 ;
        RECT 158.955 -141.605 159.285 -141.275 ;
        RECT 158.955 -142.965 159.285 -142.635 ;
        RECT 158.955 -144.325 159.285 -143.995 ;
        RECT 158.955 -145.685 159.285 -145.355 ;
        RECT 158.955 -147.045 159.285 -146.715 ;
        RECT 158.955 -148.405 159.285 -148.075 ;
        RECT 158.955 -149.765 159.285 -149.435 ;
        RECT 158.955 -151.125 159.285 -150.795 ;
        RECT 158.955 -152.485 159.285 -152.155 ;
        RECT 158.955 -153.845 159.285 -153.515 ;
        RECT 158.955 -155.205 159.285 -154.875 ;
        RECT 158.955 -156.565 159.285 -156.235 ;
        RECT 158.955 -157.925 159.285 -157.595 ;
        RECT 158.955 -159.285 159.285 -158.955 ;
        RECT 158.955 -160.645 159.285 -160.315 ;
        RECT 158.955 -162.005 159.285 -161.675 ;
        RECT 158.955 -163.365 159.285 -163.035 ;
        RECT 158.955 -164.725 159.285 -164.395 ;
        RECT 158.955 -166.085 159.285 -165.755 ;
        RECT 158.955 -167.445 159.285 -167.115 ;
        RECT 158.955 -168.805 159.285 -168.475 ;
        RECT 158.955 -170.165 159.285 -169.835 ;
        RECT 158.955 -171.525 159.285 -171.195 ;
        RECT 158.955 -172.885 159.285 -172.555 ;
        RECT 158.955 -174.245 159.285 -173.915 ;
        RECT 158.955 -175.605 159.285 -175.275 ;
        RECT 158.955 -176.965 159.285 -176.635 ;
        RECT 158.955 -178.325 159.285 -177.995 ;
        RECT 158.955 -180.57 159.285 -179.44 ;
        RECT 158.96 -180.685 159.28 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 160.315 241.32 160.645 242.45 ;
        RECT 160.315 239.195 160.645 239.525 ;
        RECT 160.315 237.835 160.645 238.165 ;
        RECT 160.32 237.16 160.64 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 160.315 -1.525 160.645 -1.195 ;
        RECT 160.315 -2.885 160.645 -2.555 ;
        RECT 160.32 -3.56 160.64 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 160.315 -91.285 160.645 -90.955 ;
        RECT 160.315 -92.645 160.645 -92.315 ;
        RECT 160.315 -94.005 160.645 -93.675 ;
        RECT 160.315 -95.365 160.645 -95.035 ;
        RECT 160.315 -96.725 160.645 -96.395 ;
        RECT 160.315 -98.085 160.645 -97.755 ;
        RECT 160.315 -99.445 160.645 -99.115 ;
        RECT 160.315 -100.805 160.645 -100.475 ;
        RECT 160.315 -102.165 160.645 -101.835 ;
        RECT 160.315 -103.525 160.645 -103.195 ;
        RECT 160.315 -104.885 160.645 -104.555 ;
        RECT 160.315 -106.245 160.645 -105.915 ;
        RECT 160.315 -107.605 160.645 -107.275 ;
        RECT 160.315 -108.965 160.645 -108.635 ;
        RECT 160.315 -110.325 160.645 -109.995 ;
        RECT 160.315 -111.685 160.645 -111.355 ;
        RECT 160.315 -113.045 160.645 -112.715 ;
        RECT 160.315 -114.405 160.645 -114.075 ;
        RECT 160.315 -115.765 160.645 -115.435 ;
        RECT 160.315 -117.125 160.645 -116.795 ;
        RECT 160.315 -118.485 160.645 -118.155 ;
        RECT 160.315 -119.845 160.645 -119.515 ;
        RECT 160.315 -121.205 160.645 -120.875 ;
        RECT 160.315 -122.565 160.645 -122.235 ;
        RECT 160.315 -123.925 160.645 -123.595 ;
        RECT 160.315 -125.285 160.645 -124.955 ;
        RECT 160.315 -126.645 160.645 -126.315 ;
        RECT 160.315 -128.005 160.645 -127.675 ;
        RECT 160.315 -129.365 160.645 -129.035 ;
        RECT 160.315 -130.725 160.645 -130.395 ;
        RECT 160.315 -132.085 160.645 -131.755 ;
        RECT 160.315 -133.445 160.645 -133.115 ;
        RECT 160.315 -134.805 160.645 -134.475 ;
        RECT 160.315 -136.165 160.645 -135.835 ;
        RECT 160.315 -137.525 160.645 -137.195 ;
        RECT 160.315 -138.885 160.645 -138.555 ;
        RECT 160.315 -140.245 160.645 -139.915 ;
        RECT 160.315 -141.605 160.645 -141.275 ;
        RECT 160.315 -142.965 160.645 -142.635 ;
        RECT 160.315 -144.325 160.645 -143.995 ;
        RECT 160.315 -145.685 160.645 -145.355 ;
        RECT 160.315 -147.045 160.645 -146.715 ;
        RECT 160.315 -148.405 160.645 -148.075 ;
        RECT 160.315 -149.765 160.645 -149.435 ;
        RECT 160.315 -151.125 160.645 -150.795 ;
        RECT 160.315 -152.485 160.645 -152.155 ;
        RECT 160.315 -153.845 160.645 -153.515 ;
        RECT 160.315 -155.205 160.645 -154.875 ;
        RECT 160.315 -156.565 160.645 -156.235 ;
        RECT 160.315 -157.925 160.645 -157.595 ;
        RECT 160.315 -159.285 160.645 -158.955 ;
        RECT 160.315 -160.645 160.645 -160.315 ;
        RECT 160.315 -162.005 160.645 -161.675 ;
        RECT 160.315 -163.365 160.645 -163.035 ;
        RECT 160.315 -164.725 160.645 -164.395 ;
        RECT 160.315 -166.085 160.645 -165.755 ;
        RECT 160.315 -167.445 160.645 -167.115 ;
        RECT 160.315 -168.805 160.645 -168.475 ;
        RECT 160.315 -170.165 160.645 -169.835 ;
        RECT 160.315 -171.525 160.645 -171.195 ;
        RECT 160.315 -172.885 160.645 -172.555 ;
        RECT 160.315 -174.245 160.645 -173.915 ;
        RECT 160.315 -175.605 160.645 -175.275 ;
        RECT 160.315 -176.965 160.645 -176.635 ;
        RECT 160.315 -178.325 160.645 -177.995 ;
        RECT 160.315 -180.57 160.645 -179.44 ;
        RECT 160.32 -180.685 160.64 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 161.675 241.32 162.005 242.45 ;
        RECT 161.675 239.195 162.005 239.525 ;
        RECT 161.675 237.835 162.005 238.165 ;
        RECT 161.68 237.16 162 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 161.675 -95.365 162.005 -95.035 ;
        RECT 161.675 -96.725 162.005 -96.395 ;
        RECT 161.675 -98.085 162.005 -97.755 ;
        RECT 161.675 -99.445 162.005 -99.115 ;
        RECT 161.675 -100.805 162.005 -100.475 ;
        RECT 161.675 -102.165 162.005 -101.835 ;
        RECT 161.675 -103.525 162.005 -103.195 ;
        RECT 161.675 -104.885 162.005 -104.555 ;
        RECT 161.675 -106.245 162.005 -105.915 ;
        RECT 161.675 -107.605 162.005 -107.275 ;
        RECT 161.675 -108.965 162.005 -108.635 ;
        RECT 161.675 -110.325 162.005 -109.995 ;
        RECT 161.675 -111.685 162.005 -111.355 ;
        RECT 161.675 -113.045 162.005 -112.715 ;
        RECT 161.675 -114.405 162.005 -114.075 ;
        RECT 161.675 -115.765 162.005 -115.435 ;
        RECT 161.675 -117.125 162.005 -116.795 ;
        RECT 161.675 -118.485 162.005 -118.155 ;
        RECT 161.675 -119.845 162.005 -119.515 ;
        RECT 161.675 -121.205 162.005 -120.875 ;
        RECT 161.675 -122.565 162.005 -122.235 ;
        RECT 161.675 -123.925 162.005 -123.595 ;
        RECT 161.675 -125.285 162.005 -124.955 ;
        RECT 161.675 -126.645 162.005 -126.315 ;
        RECT 161.675 -128.005 162.005 -127.675 ;
        RECT 161.675 -129.365 162.005 -129.035 ;
        RECT 161.675 -130.725 162.005 -130.395 ;
        RECT 161.675 -132.085 162.005 -131.755 ;
        RECT 161.675 -133.445 162.005 -133.115 ;
        RECT 161.675 -134.805 162.005 -134.475 ;
        RECT 161.675 -136.165 162.005 -135.835 ;
        RECT 161.675 -137.525 162.005 -137.195 ;
        RECT 161.675 -138.885 162.005 -138.555 ;
        RECT 161.675 -140.245 162.005 -139.915 ;
        RECT 161.675 -141.605 162.005 -141.275 ;
        RECT 161.675 -142.965 162.005 -142.635 ;
        RECT 161.675 -144.325 162.005 -143.995 ;
        RECT 161.675 -145.685 162.005 -145.355 ;
        RECT 161.675 -147.045 162.005 -146.715 ;
        RECT 161.675 -148.405 162.005 -148.075 ;
        RECT 161.675 -149.765 162.005 -149.435 ;
        RECT 161.675 -151.125 162.005 -150.795 ;
        RECT 161.675 -152.485 162.005 -152.155 ;
        RECT 161.675 -153.845 162.005 -153.515 ;
        RECT 161.675 -155.205 162.005 -154.875 ;
        RECT 161.675 -156.565 162.005 -156.235 ;
        RECT 161.675 -157.925 162.005 -157.595 ;
        RECT 161.675 -159.285 162.005 -158.955 ;
        RECT 161.675 -160.645 162.005 -160.315 ;
        RECT 161.675 -162.005 162.005 -161.675 ;
        RECT 161.675 -163.365 162.005 -163.035 ;
        RECT 161.675 -164.725 162.005 -164.395 ;
        RECT 161.675 -166.085 162.005 -165.755 ;
        RECT 161.675 -167.445 162.005 -167.115 ;
        RECT 161.675 -168.805 162.005 -168.475 ;
        RECT 161.675 -170.165 162.005 -169.835 ;
        RECT 161.675 -171.525 162.005 -171.195 ;
        RECT 161.675 -172.885 162.005 -172.555 ;
        RECT 161.675 -174.245 162.005 -173.915 ;
        RECT 161.675 -175.605 162.005 -175.275 ;
        RECT 161.675 -176.965 162.005 -176.635 ;
        RECT 161.675 -178.325 162.005 -177.995 ;
        RECT 161.675 -180.57 162.005 -179.44 ;
        RECT 161.68 -180.685 162 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 161.91 -94.075 162.24 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 163.035 241.32 163.365 242.45 ;
        RECT 163.035 239.195 163.365 239.525 ;
        RECT 163.035 237.835 163.365 238.165 ;
        RECT 163.04 237.16 163.36 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 163.035 -1.525 163.365 -1.195 ;
        RECT 163.035 -2.885 163.365 -2.555 ;
        RECT 163.04 -3.56 163.36 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 164.395 241.32 164.725 242.45 ;
        RECT 164.395 239.195 164.725 239.525 ;
        RECT 164.395 237.835 164.725 238.165 ;
        RECT 164.4 237.16 164.72 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 164.395 -1.525 164.725 -1.195 ;
        RECT 164.395 -2.885 164.725 -2.555 ;
        RECT 164.4 -3.56 164.72 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 165.755 241.32 166.085 242.45 ;
        RECT 165.755 239.195 166.085 239.525 ;
        RECT 165.755 237.835 166.085 238.165 ;
        RECT 165.76 237.16 166.08 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 165.755 -1.525 166.085 -1.195 ;
        RECT 165.755 -2.885 166.085 -2.555 ;
        RECT 165.76 -3.56 166.08 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 165.755 -91.285 166.085 -90.955 ;
        RECT 165.755 -92.645 166.085 -92.315 ;
        RECT 165.755 -94.005 166.085 -93.675 ;
        RECT 165.755 -95.365 166.085 -95.035 ;
        RECT 165.755 -96.725 166.085 -96.395 ;
        RECT 165.755 -98.085 166.085 -97.755 ;
        RECT 165.755 -99.445 166.085 -99.115 ;
        RECT 165.755 -100.805 166.085 -100.475 ;
        RECT 165.755 -102.165 166.085 -101.835 ;
        RECT 165.755 -103.525 166.085 -103.195 ;
        RECT 165.755 -104.885 166.085 -104.555 ;
        RECT 165.755 -106.245 166.085 -105.915 ;
        RECT 165.755 -107.605 166.085 -107.275 ;
        RECT 165.755 -108.965 166.085 -108.635 ;
        RECT 165.755 -110.325 166.085 -109.995 ;
        RECT 165.755 -111.685 166.085 -111.355 ;
        RECT 165.755 -113.045 166.085 -112.715 ;
        RECT 165.755 -114.405 166.085 -114.075 ;
        RECT 165.755 -115.765 166.085 -115.435 ;
        RECT 165.755 -117.125 166.085 -116.795 ;
        RECT 165.755 -118.485 166.085 -118.155 ;
        RECT 165.755 -119.845 166.085 -119.515 ;
        RECT 165.755 -121.205 166.085 -120.875 ;
        RECT 165.755 -122.565 166.085 -122.235 ;
        RECT 165.755 -123.925 166.085 -123.595 ;
        RECT 165.755 -125.285 166.085 -124.955 ;
        RECT 165.755 -126.645 166.085 -126.315 ;
        RECT 165.755 -128.005 166.085 -127.675 ;
        RECT 165.755 -129.365 166.085 -129.035 ;
        RECT 165.755 -130.725 166.085 -130.395 ;
        RECT 165.755 -132.085 166.085 -131.755 ;
        RECT 165.755 -133.445 166.085 -133.115 ;
        RECT 165.755 -134.805 166.085 -134.475 ;
        RECT 165.755 -136.165 166.085 -135.835 ;
        RECT 165.755 -137.525 166.085 -137.195 ;
        RECT 165.755 -138.885 166.085 -138.555 ;
        RECT 165.755 -140.245 166.085 -139.915 ;
        RECT 165.755 -141.605 166.085 -141.275 ;
        RECT 165.755 -142.965 166.085 -142.635 ;
        RECT 165.755 -144.325 166.085 -143.995 ;
        RECT 165.755 -145.685 166.085 -145.355 ;
        RECT 165.755 -147.045 166.085 -146.715 ;
        RECT 165.755 -148.405 166.085 -148.075 ;
        RECT 165.755 -149.765 166.085 -149.435 ;
        RECT 165.755 -151.125 166.085 -150.795 ;
        RECT 165.755 -152.485 166.085 -152.155 ;
        RECT 165.755 -153.845 166.085 -153.515 ;
        RECT 165.755 -155.205 166.085 -154.875 ;
        RECT 165.755 -156.565 166.085 -156.235 ;
        RECT 165.755 -157.925 166.085 -157.595 ;
        RECT 165.755 -159.285 166.085 -158.955 ;
        RECT 165.755 -160.645 166.085 -160.315 ;
        RECT 165.755 -162.005 166.085 -161.675 ;
        RECT 165.755 -163.365 166.085 -163.035 ;
        RECT 165.755 -164.725 166.085 -164.395 ;
        RECT 165.755 -166.085 166.085 -165.755 ;
        RECT 165.755 -167.445 166.085 -167.115 ;
        RECT 165.755 -168.805 166.085 -168.475 ;
        RECT 165.755 -170.165 166.085 -169.835 ;
        RECT 165.755 -171.525 166.085 -171.195 ;
        RECT 165.755 -172.885 166.085 -172.555 ;
        RECT 165.755 -174.245 166.085 -173.915 ;
        RECT 165.755 -175.605 166.085 -175.275 ;
        RECT 165.755 -176.965 166.085 -176.635 ;
        RECT 165.755 -178.325 166.085 -177.995 ;
        RECT 165.755 -180.57 166.085 -179.44 ;
        RECT 165.76 -180.685 166.08 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 167.115 241.32 167.445 242.45 ;
        RECT 167.115 239.195 167.445 239.525 ;
        RECT 167.115 237.835 167.445 238.165 ;
        RECT 167.12 237.16 167.44 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 167.115 -95.365 167.445 -95.035 ;
        RECT 167.115 -96.725 167.445 -96.395 ;
        RECT 167.115 -98.085 167.445 -97.755 ;
        RECT 167.115 -99.445 167.445 -99.115 ;
        RECT 167.115 -100.805 167.445 -100.475 ;
        RECT 167.115 -102.165 167.445 -101.835 ;
        RECT 167.115 -103.525 167.445 -103.195 ;
        RECT 167.115 -104.885 167.445 -104.555 ;
        RECT 167.115 -106.245 167.445 -105.915 ;
        RECT 167.115 -107.605 167.445 -107.275 ;
        RECT 167.115 -108.965 167.445 -108.635 ;
        RECT 167.115 -110.325 167.445 -109.995 ;
        RECT 167.115 -111.685 167.445 -111.355 ;
        RECT 167.115 -113.045 167.445 -112.715 ;
        RECT 167.115 -114.405 167.445 -114.075 ;
        RECT 167.115 -115.765 167.445 -115.435 ;
        RECT 167.115 -117.125 167.445 -116.795 ;
        RECT 167.115 -118.485 167.445 -118.155 ;
        RECT 167.115 -119.845 167.445 -119.515 ;
        RECT 167.115 -121.205 167.445 -120.875 ;
        RECT 167.115 -122.565 167.445 -122.235 ;
        RECT 167.115 -123.925 167.445 -123.595 ;
        RECT 167.115 -125.285 167.445 -124.955 ;
        RECT 167.115 -126.645 167.445 -126.315 ;
        RECT 167.115 -128.005 167.445 -127.675 ;
        RECT 167.115 -129.365 167.445 -129.035 ;
        RECT 167.115 -130.725 167.445 -130.395 ;
        RECT 167.115 -132.085 167.445 -131.755 ;
        RECT 167.115 -133.445 167.445 -133.115 ;
        RECT 167.115 -134.805 167.445 -134.475 ;
        RECT 167.115 -136.165 167.445 -135.835 ;
        RECT 167.115 -137.525 167.445 -137.195 ;
        RECT 167.115 -138.885 167.445 -138.555 ;
        RECT 167.115 -140.245 167.445 -139.915 ;
        RECT 167.115 -141.605 167.445 -141.275 ;
        RECT 167.115 -142.965 167.445 -142.635 ;
        RECT 167.115 -144.325 167.445 -143.995 ;
        RECT 167.115 -145.685 167.445 -145.355 ;
        RECT 167.115 -147.045 167.445 -146.715 ;
        RECT 167.115 -148.405 167.445 -148.075 ;
        RECT 167.115 -149.765 167.445 -149.435 ;
        RECT 167.115 -151.125 167.445 -150.795 ;
        RECT 167.115 -152.485 167.445 -152.155 ;
        RECT 167.115 -153.845 167.445 -153.515 ;
        RECT 167.115 -155.205 167.445 -154.875 ;
        RECT 167.115 -156.565 167.445 -156.235 ;
        RECT 167.115 -157.925 167.445 -157.595 ;
        RECT 167.115 -159.285 167.445 -158.955 ;
        RECT 167.115 -160.645 167.445 -160.315 ;
        RECT 167.115 -162.005 167.445 -161.675 ;
        RECT 167.115 -163.365 167.445 -163.035 ;
        RECT 167.115 -164.725 167.445 -164.395 ;
        RECT 167.115 -166.085 167.445 -165.755 ;
        RECT 167.115 -167.445 167.445 -167.115 ;
        RECT 167.115 -168.805 167.445 -168.475 ;
        RECT 167.115 -170.165 167.445 -169.835 ;
        RECT 167.115 -171.525 167.445 -171.195 ;
        RECT 167.115 -172.885 167.445 -172.555 ;
        RECT 167.115 -174.245 167.445 -173.915 ;
        RECT 167.115 -175.605 167.445 -175.275 ;
        RECT 167.115 -176.965 167.445 -176.635 ;
        RECT 167.115 -178.325 167.445 -177.995 ;
        RECT 167.115 -180.57 167.445 -179.44 ;
        RECT 167.12 -180.685 167.44 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 168.01 -94.075 168.34 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 168.475 241.32 168.805 242.45 ;
        RECT 168.475 239.195 168.805 239.525 ;
        RECT 168.475 237.835 168.805 238.165 ;
        RECT 168.48 237.16 168.8 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 169.835 241.32 170.165 242.45 ;
        RECT 169.835 239.195 170.165 239.525 ;
        RECT 169.835 237.835 170.165 238.165 ;
        RECT 169.84 237.16 170.16 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 169.835 -1.525 170.165 -1.195 ;
        RECT 169.835 -2.885 170.165 -2.555 ;
        RECT 169.84 -3.56 170.16 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 171.195 241.32 171.525 242.45 ;
        RECT 171.195 239.195 171.525 239.525 ;
        RECT 171.195 237.835 171.525 238.165 ;
        RECT 171.2 237.16 171.52 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 171.195 -1.525 171.525 -1.195 ;
        RECT 171.195 -2.885 171.525 -2.555 ;
        RECT 171.2 -3.56 171.52 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 171.195 -91.285 171.525 -90.955 ;
        RECT 171.195 -92.645 171.525 -92.315 ;
        RECT 171.195 -94.005 171.525 -93.675 ;
        RECT 171.195 -95.365 171.525 -95.035 ;
        RECT 171.195 -96.725 171.525 -96.395 ;
        RECT 171.195 -98.085 171.525 -97.755 ;
        RECT 171.195 -99.445 171.525 -99.115 ;
        RECT 171.195 -100.805 171.525 -100.475 ;
        RECT 171.195 -102.165 171.525 -101.835 ;
        RECT 171.195 -103.525 171.525 -103.195 ;
        RECT 171.195 -104.885 171.525 -104.555 ;
        RECT 171.195 -106.245 171.525 -105.915 ;
        RECT 171.195 -107.605 171.525 -107.275 ;
        RECT 171.195 -108.965 171.525 -108.635 ;
        RECT 171.195 -110.325 171.525 -109.995 ;
        RECT 171.195 -111.685 171.525 -111.355 ;
        RECT 171.195 -113.045 171.525 -112.715 ;
        RECT 171.195 -114.405 171.525 -114.075 ;
        RECT 171.195 -115.765 171.525 -115.435 ;
        RECT 171.195 -117.125 171.525 -116.795 ;
        RECT 171.195 -118.485 171.525 -118.155 ;
        RECT 171.195 -119.845 171.525 -119.515 ;
        RECT 171.195 -121.205 171.525 -120.875 ;
        RECT 171.195 -122.565 171.525 -122.235 ;
        RECT 171.195 -123.925 171.525 -123.595 ;
        RECT 171.195 -125.285 171.525 -124.955 ;
        RECT 171.195 -126.645 171.525 -126.315 ;
        RECT 171.195 -128.005 171.525 -127.675 ;
        RECT 171.195 -129.365 171.525 -129.035 ;
        RECT 171.195 -130.725 171.525 -130.395 ;
        RECT 171.195 -132.085 171.525 -131.755 ;
        RECT 171.195 -133.445 171.525 -133.115 ;
        RECT 171.195 -134.805 171.525 -134.475 ;
        RECT 171.195 -136.165 171.525 -135.835 ;
        RECT 171.195 -137.525 171.525 -137.195 ;
        RECT 171.195 -138.885 171.525 -138.555 ;
        RECT 171.195 -140.245 171.525 -139.915 ;
        RECT 171.195 -141.605 171.525 -141.275 ;
        RECT 171.195 -142.965 171.525 -142.635 ;
        RECT 171.195 -144.325 171.525 -143.995 ;
        RECT 171.195 -145.685 171.525 -145.355 ;
        RECT 171.195 -147.045 171.525 -146.715 ;
        RECT 171.195 -148.405 171.525 -148.075 ;
        RECT 171.195 -149.765 171.525 -149.435 ;
        RECT 171.195 -151.125 171.525 -150.795 ;
        RECT 171.195 -152.485 171.525 -152.155 ;
        RECT 171.195 -153.845 171.525 -153.515 ;
        RECT 171.195 -155.205 171.525 -154.875 ;
        RECT 171.195 -156.565 171.525 -156.235 ;
        RECT 171.195 -157.925 171.525 -157.595 ;
        RECT 171.195 -159.285 171.525 -158.955 ;
        RECT 171.195 -160.645 171.525 -160.315 ;
        RECT 171.195 -162.005 171.525 -161.675 ;
        RECT 171.195 -163.365 171.525 -163.035 ;
        RECT 171.195 -164.725 171.525 -164.395 ;
        RECT 171.195 -166.085 171.525 -165.755 ;
        RECT 171.195 -167.445 171.525 -167.115 ;
        RECT 171.195 -168.805 171.525 -168.475 ;
        RECT 171.195 -170.165 171.525 -169.835 ;
        RECT 171.195 -171.525 171.525 -171.195 ;
        RECT 171.195 -172.885 171.525 -172.555 ;
        RECT 171.195 -174.245 171.525 -173.915 ;
        RECT 171.195 -175.605 171.525 -175.275 ;
        RECT 171.195 -176.965 171.525 -176.635 ;
        RECT 171.195 -178.325 171.525 -177.995 ;
        RECT 171.195 -180.57 171.525 -179.44 ;
        RECT 171.2 -180.685 171.52 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 172.555 241.32 172.885 242.45 ;
        RECT 172.555 239.195 172.885 239.525 ;
        RECT 172.555 237.835 172.885 238.165 ;
        RECT 172.56 237.16 172.88 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 172.555 -1.525 172.885 -1.195 ;
        RECT 172.555 -2.885 172.885 -2.555 ;
        RECT 172.56 -3.56 172.88 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 172.56 -180.685 172.88 -90.955 ;
        RECT 172.555 -91.285 172.885 -90.955 ;
        RECT 172.555 -92.645 172.885 -92.315 ;
        RECT 172.555 -94.005 172.885 -93.675 ;
        RECT 172.555 -95.365 172.885 -95.035 ;
        RECT 172.555 -96.725 172.885 -96.395 ;
        RECT 172.555 -98.085 172.885 -97.755 ;
        RECT 172.555 -99.445 172.885 -99.115 ;
        RECT 172.555 -100.805 172.885 -100.475 ;
        RECT 172.555 -102.165 172.885 -101.835 ;
        RECT 172.555 -103.525 172.885 -103.195 ;
        RECT 172.555 -104.885 172.885 -104.555 ;
        RECT 172.555 -106.245 172.885 -105.915 ;
        RECT 172.555 -107.605 172.885 -107.275 ;
        RECT 172.555 -108.965 172.885 -108.635 ;
        RECT 172.555 -110.325 172.885 -109.995 ;
        RECT 172.555 -111.685 172.885 -111.355 ;
        RECT 172.555 -113.045 172.885 -112.715 ;
        RECT 172.555 -114.405 172.885 -114.075 ;
        RECT 172.555 -115.765 172.885 -115.435 ;
        RECT 172.555 -117.125 172.885 -116.795 ;
        RECT 172.555 -118.485 172.885 -118.155 ;
        RECT 172.555 -119.845 172.885 -119.515 ;
        RECT 172.555 -121.205 172.885 -120.875 ;
        RECT 172.555 -122.565 172.885 -122.235 ;
        RECT 172.555 -123.925 172.885 -123.595 ;
        RECT 172.555 -125.285 172.885 -124.955 ;
        RECT 172.555 -126.645 172.885 -126.315 ;
        RECT 172.555 -128.005 172.885 -127.675 ;
        RECT 172.555 -129.365 172.885 -129.035 ;
        RECT 172.555 -130.725 172.885 -130.395 ;
        RECT 172.555 -132.085 172.885 -131.755 ;
        RECT 172.555 -133.445 172.885 -133.115 ;
        RECT 172.555 -134.805 172.885 -134.475 ;
        RECT 172.555 -136.165 172.885 -135.835 ;
        RECT 172.555 -137.525 172.885 -137.195 ;
        RECT 172.555 -138.885 172.885 -138.555 ;
        RECT 172.555 -140.245 172.885 -139.915 ;
        RECT 172.555 -141.605 172.885 -141.275 ;
        RECT 172.555 -142.965 172.885 -142.635 ;
        RECT 172.555 -144.325 172.885 -143.995 ;
        RECT 172.555 -145.685 172.885 -145.355 ;
        RECT 172.555 -147.045 172.885 -146.715 ;
        RECT 172.555 -148.405 172.885 -148.075 ;
        RECT 172.555 -149.765 172.885 -149.435 ;
        RECT 172.555 -151.125 172.885 -150.795 ;
        RECT 172.555 -152.485 172.885 -152.155 ;
        RECT 172.555 -153.845 172.885 -153.515 ;
        RECT 172.555 -155.205 172.885 -154.875 ;
        RECT 172.555 -156.565 172.885 -156.235 ;
        RECT 172.555 -157.925 172.885 -157.595 ;
        RECT 172.555 -159.285 172.885 -158.955 ;
        RECT 172.555 -160.645 172.885 -160.315 ;
        RECT 172.555 -162.005 172.885 -161.675 ;
        RECT 172.555 -163.365 172.885 -163.035 ;
        RECT 172.555 -164.725 172.885 -164.395 ;
        RECT 172.555 -166.085 172.885 -165.755 ;
        RECT 172.555 -167.445 172.885 -167.115 ;
        RECT 172.555 -168.805 172.885 -168.475 ;
        RECT 172.555 -170.165 172.885 -169.835 ;
        RECT 172.555 -171.525 172.885 -171.195 ;
        RECT 172.555 -172.885 172.885 -172.555 ;
        RECT 172.555 -174.245 172.885 -173.915 ;
        RECT 172.555 -175.605 172.885 -175.275 ;
        RECT 172.555 -176.965 172.885 -176.635 ;
        RECT 172.555 -178.325 172.885 -177.995 ;
        RECT 172.555 -180.57 172.885 -179.44 ;
    END
    PORT
      LAYER met3 ;
        RECT 100.475 241.32 100.805 242.45 ;
        RECT 100.475 239.195 100.805 239.525 ;
        RECT 100.475 237.835 100.805 238.165 ;
        RECT 100.48 237.16 100.8 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 100.475 -95.365 100.805 -95.035 ;
        RECT 100.475 -96.725 100.805 -96.395 ;
        RECT 100.475 -98.085 100.805 -97.755 ;
        RECT 100.475 -99.445 100.805 -99.115 ;
        RECT 100.475 -100.805 100.805 -100.475 ;
        RECT 100.475 -102.165 100.805 -101.835 ;
        RECT 100.475 -103.525 100.805 -103.195 ;
        RECT 100.475 -104.885 100.805 -104.555 ;
        RECT 100.475 -106.245 100.805 -105.915 ;
        RECT 100.475 -107.605 100.805 -107.275 ;
        RECT 100.475 -108.965 100.805 -108.635 ;
        RECT 100.475 -110.325 100.805 -109.995 ;
        RECT 100.475 -111.685 100.805 -111.355 ;
        RECT 100.475 -113.045 100.805 -112.715 ;
        RECT 100.475 -114.405 100.805 -114.075 ;
        RECT 100.475 -115.765 100.805 -115.435 ;
        RECT 100.475 -117.125 100.805 -116.795 ;
        RECT 100.475 -118.485 100.805 -118.155 ;
        RECT 100.475 -119.845 100.805 -119.515 ;
        RECT 100.475 -121.205 100.805 -120.875 ;
        RECT 100.475 -122.565 100.805 -122.235 ;
        RECT 100.475 -123.925 100.805 -123.595 ;
        RECT 100.475 -125.285 100.805 -124.955 ;
        RECT 100.475 -126.645 100.805 -126.315 ;
        RECT 100.475 -128.005 100.805 -127.675 ;
        RECT 100.475 -129.365 100.805 -129.035 ;
        RECT 100.475 -130.725 100.805 -130.395 ;
        RECT 100.475 -132.085 100.805 -131.755 ;
        RECT 100.475 -133.445 100.805 -133.115 ;
        RECT 100.475 -134.805 100.805 -134.475 ;
        RECT 100.475 -136.165 100.805 -135.835 ;
        RECT 100.475 -137.525 100.805 -137.195 ;
        RECT 100.475 -138.885 100.805 -138.555 ;
        RECT 100.475 -140.245 100.805 -139.915 ;
        RECT 100.475 -141.605 100.805 -141.275 ;
        RECT 100.475 -142.965 100.805 -142.635 ;
        RECT 100.475 -144.325 100.805 -143.995 ;
        RECT 100.475 -145.685 100.805 -145.355 ;
        RECT 100.475 -147.045 100.805 -146.715 ;
        RECT 100.475 -148.405 100.805 -148.075 ;
        RECT 100.475 -149.765 100.805 -149.435 ;
        RECT 100.475 -151.125 100.805 -150.795 ;
        RECT 100.475 -152.485 100.805 -152.155 ;
        RECT 100.475 -153.845 100.805 -153.515 ;
        RECT 100.475 -155.205 100.805 -154.875 ;
        RECT 100.475 -156.565 100.805 -156.235 ;
        RECT 100.475 -157.925 100.805 -157.595 ;
        RECT 100.475 -159.285 100.805 -158.955 ;
        RECT 100.475 -160.645 100.805 -160.315 ;
        RECT 100.475 -162.005 100.805 -161.675 ;
        RECT 100.475 -163.365 100.805 -163.035 ;
        RECT 100.475 -164.725 100.805 -164.395 ;
        RECT 100.475 -166.085 100.805 -165.755 ;
        RECT 100.475 -167.445 100.805 -167.115 ;
        RECT 100.475 -168.805 100.805 -168.475 ;
        RECT 100.475 -170.165 100.805 -169.835 ;
        RECT 100.475 -171.525 100.805 -171.195 ;
        RECT 100.475 -172.885 100.805 -172.555 ;
        RECT 100.475 -174.245 100.805 -173.915 ;
        RECT 100.475 -175.605 100.805 -175.275 ;
        RECT 100.475 -176.965 100.805 -176.635 ;
        RECT 100.475 -178.325 100.805 -177.995 ;
        RECT 100.475 -180.57 100.805 -179.44 ;
        RECT 100.48 -180.685 100.8 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 100.91 -94.075 101.24 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 101.835 241.32 102.165 242.45 ;
        RECT 101.835 239.195 102.165 239.525 ;
        RECT 101.835 237.835 102.165 238.165 ;
        RECT 101.84 237.16 102.16 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 101.835 -1.525 102.165 -1.195 ;
        RECT 101.835 -2.885 102.165 -2.555 ;
        RECT 101.84 -3.56 102.16 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 103.195 241.32 103.525 242.45 ;
        RECT 103.195 239.195 103.525 239.525 ;
        RECT 103.195 237.835 103.525 238.165 ;
        RECT 103.2 237.16 103.52 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 103.195 -1.525 103.525 -1.195 ;
        RECT 103.195 -2.885 103.525 -2.555 ;
        RECT 103.2 -3.56 103.52 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 104.555 241.32 104.885 242.45 ;
        RECT 104.555 239.195 104.885 239.525 ;
        RECT 104.555 237.835 104.885 238.165 ;
        RECT 104.56 237.16 104.88 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 104.555 -1.525 104.885 -1.195 ;
        RECT 104.555 -2.885 104.885 -2.555 ;
        RECT 104.56 -3.56 104.88 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 105.915 241.32 106.245 242.45 ;
        RECT 105.915 239.195 106.245 239.525 ;
        RECT 105.915 237.835 106.245 238.165 ;
        RECT 105.92 237.16 106.24 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 105.915 -95.365 106.245 -95.035 ;
        RECT 105.915 -96.725 106.245 -96.395 ;
        RECT 105.915 -98.085 106.245 -97.755 ;
        RECT 105.915 -99.445 106.245 -99.115 ;
        RECT 105.915 -100.805 106.245 -100.475 ;
        RECT 105.915 -102.165 106.245 -101.835 ;
        RECT 105.915 -103.525 106.245 -103.195 ;
        RECT 105.915 -104.885 106.245 -104.555 ;
        RECT 105.915 -106.245 106.245 -105.915 ;
        RECT 105.915 -107.605 106.245 -107.275 ;
        RECT 105.915 -108.965 106.245 -108.635 ;
        RECT 105.915 -110.325 106.245 -109.995 ;
        RECT 105.915 -111.685 106.245 -111.355 ;
        RECT 105.915 -113.045 106.245 -112.715 ;
        RECT 105.915 -114.405 106.245 -114.075 ;
        RECT 105.915 -115.765 106.245 -115.435 ;
        RECT 105.915 -117.125 106.245 -116.795 ;
        RECT 105.915 -118.485 106.245 -118.155 ;
        RECT 105.915 -119.845 106.245 -119.515 ;
        RECT 105.915 -121.205 106.245 -120.875 ;
        RECT 105.915 -122.565 106.245 -122.235 ;
        RECT 105.915 -123.925 106.245 -123.595 ;
        RECT 105.915 -125.285 106.245 -124.955 ;
        RECT 105.915 -126.645 106.245 -126.315 ;
        RECT 105.915 -128.005 106.245 -127.675 ;
        RECT 105.915 -129.365 106.245 -129.035 ;
        RECT 105.915 -130.725 106.245 -130.395 ;
        RECT 105.915 -132.085 106.245 -131.755 ;
        RECT 105.915 -133.445 106.245 -133.115 ;
        RECT 105.915 -134.805 106.245 -134.475 ;
        RECT 105.915 -136.165 106.245 -135.835 ;
        RECT 105.915 -137.525 106.245 -137.195 ;
        RECT 105.915 -138.885 106.245 -138.555 ;
        RECT 105.915 -140.245 106.245 -139.915 ;
        RECT 105.915 -141.605 106.245 -141.275 ;
        RECT 105.915 -142.965 106.245 -142.635 ;
        RECT 105.915 -144.325 106.245 -143.995 ;
        RECT 105.915 -145.685 106.245 -145.355 ;
        RECT 105.915 -147.045 106.245 -146.715 ;
        RECT 105.915 -148.405 106.245 -148.075 ;
        RECT 105.915 -149.765 106.245 -149.435 ;
        RECT 105.915 -151.125 106.245 -150.795 ;
        RECT 105.915 -152.485 106.245 -152.155 ;
        RECT 105.915 -153.845 106.245 -153.515 ;
        RECT 105.915 -155.205 106.245 -154.875 ;
        RECT 105.915 -156.565 106.245 -156.235 ;
        RECT 105.915 -157.925 106.245 -157.595 ;
        RECT 105.915 -159.285 106.245 -158.955 ;
        RECT 105.915 -160.645 106.245 -160.315 ;
        RECT 105.915 -162.005 106.245 -161.675 ;
        RECT 105.915 -163.365 106.245 -163.035 ;
        RECT 105.915 -164.725 106.245 -164.395 ;
        RECT 105.915 -166.085 106.245 -165.755 ;
        RECT 105.915 -167.445 106.245 -167.115 ;
        RECT 105.915 -168.805 106.245 -168.475 ;
        RECT 105.915 -170.165 106.245 -169.835 ;
        RECT 105.915 -171.525 106.245 -171.195 ;
        RECT 105.915 -172.885 106.245 -172.555 ;
        RECT 105.915 -174.245 106.245 -173.915 ;
        RECT 105.915 -175.605 106.245 -175.275 ;
        RECT 105.915 -176.965 106.245 -176.635 ;
        RECT 105.915 -178.325 106.245 -177.995 ;
        RECT 105.915 -180.57 106.245 -179.44 ;
        RECT 105.92 -180.685 106.24 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 107.01 -94.075 107.34 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 107.275 241.32 107.605 242.45 ;
        RECT 107.275 239.195 107.605 239.525 ;
        RECT 107.275 237.835 107.605 238.165 ;
        RECT 107.28 237.16 107.6 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 108.635 241.32 108.965 242.45 ;
        RECT 108.635 239.195 108.965 239.525 ;
        RECT 108.635 237.835 108.965 238.165 ;
        RECT 108.64 237.16 108.96 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 108.635 -1.525 108.965 -1.195 ;
        RECT 108.635 -2.885 108.965 -2.555 ;
        RECT 108.64 -3.56 108.96 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 109.995 241.32 110.325 242.45 ;
        RECT 109.995 239.195 110.325 239.525 ;
        RECT 109.995 237.835 110.325 238.165 ;
        RECT 110 237.16 110.32 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 109.995 -1.525 110.325 -1.195 ;
        RECT 109.995 -2.885 110.325 -2.555 ;
        RECT 110 -3.56 110.32 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 111.355 241.32 111.685 242.45 ;
        RECT 111.355 239.195 111.685 239.525 ;
        RECT 111.355 237.835 111.685 238.165 ;
        RECT 111.36 237.16 111.68 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 111.355 -1.525 111.685 -1.195 ;
        RECT 111.355 -2.885 111.685 -2.555 ;
        RECT 111.36 -3.56 111.68 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 111.355 -91.285 111.685 -90.955 ;
        RECT 111.355 -92.645 111.685 -92.315 ;
        RECT 111.355 -94.005 111.685 -93.675 ;
        RECT 111.355 -95.365 111.685 -95.035 ;
        RECT 111.355 -96.725 111.685 -96.395 ;
        RECT 111.355 -98.085 111.685 -97.755 ;
        RECT 111.355 -99.445 111.685 -99.115 ;
        RECT 111.355 -100.805 111.685 -100.475 ;
        RECT 111.355 -102.165 111.685 -101.835 ;
        RECT 111.355 -103.525 111.685 -103.195 ;
        RECT 111.355 -104.885 111.685 -104.555 ;
        RECT 111.355 -106.245 111.685 -105.915 ;
        RECT 111.355 -107.605 111.685 -107.275 ;
        RECT 111.355 -108.965 111.685 -108.635 ;
        RECT 111.355 -110.325 111.685 -109.995 ;
        RECT 111.355 -111.685 111.685 -111.355 ;
        RECT 111.355 -113.045 111.685 -112.715 ;
        RECT 111.355 -114.405 111.685 -114.075 ;
        RECT 111.355 -115.765 111.685 -115.435 ;
        RECT 111.355 -117.125 111.685 -116.795 ;
        RECT 111.355 -118.485 111.685 -118.155 ;
        RECT 111.355 -119.845 111.685 -119.515 ;
        RECT 111.355 -121.205 111.685 -120.875 ;
        RECT 111.355 -122.565 111.685 -122.235 ;
        RECT 111.355 -123.925 111.685 -123.595 ;
        RECT 111.355 -125.285 111.685 -124.955 ;
        RECT 111.355 -126.645 111.685 -126.315 ;
        RECT 111.355 -128.005 111.685 -127.675 ;
        RECT 111.355 -129.365 111.685 -129.035 ;
        RECT 111.355 -130.725 111.685 -130.395 ;
        RECT 111.355 -132.085 111.685 -131.755 ;
        RECT 111.355 -133.445 111.685 -133.115 ;
        RECT 111.355 -134.805 111.685 -134.475 ;
        RECT 111.355 -136.165 111.685 -135.835 ;
        RECT 111.355 -137.525 111.685 -137.195 ;
        RECT 111.355 -138.885 111.685 -138.555 ;
        RECT 111.355 -140.245 111.685 -139.915 ;
        RECT 111.355 -141.605 111.685 -141.275 ;
        RECT 111.355 -142.965 111.685 -142.635 ;
        RECT 111.355 -144.325 111.685 -143.995 ;
        RECT 111.355 -145.685 111.685 -145.355 ;
        RECT 111.355 -147.045 111.685 -146.715 ;
        RECT 111.355 -148.405 111.685 -148.075 ;
        RECT 111.355 -149.765 111.685 -149.435 ;
        RECT 111.355 -151.125 111.685 -150.795 ;
        RECT 111.355 -152.485 111.685 -152.155 ;
        RECT 111.355 -153.845 111.685 -153.515 ;
        RECT 111.355 -155.205 111.685 -154.875 ;
        RECT 111.355 -156.565 111.685 -156.235 ;
        RECT 111.355 -157.925 111.685 -157.595 ;
        RECT 111.355 -159.285 111.685 -158.955 ;
        RECT 111.355 -160.645 111.685 -160.315 ;
        RECT 111.355 -162.005 111.685 -161.675 ;
        RECT 111.355 -163.365 111.685 -163.035 ;
        RECT 111.355 -164.725 111.685 -164.395 ;
        RECT 111.355 -166.085 111.685 -165.755 ;
        RECT 111.355 -167.445 111.685 -167.115 ;
        RECT 111.355 -168.805 111.685 -168.475 ;
        RECT 111.355 -170.165 111.685 -169.835 ;
        RECT 111.355 -171.525 111.685 -171.195 ;
        RECT 111.355 -172.885 111.685 -172.555 ;
        RECT 111.355 -174.245 111.685 -173.915 ;
        RECT 111.355 -175.605 111.685 -175.275 ;
        RECT 111.355 -176.965 111.685 -176.635 ;
        RECT 111.355 -178.325 111.685 -177.995 ;
        RECT 111.355 -180.57 111.685 -179.44 ;
        RECT 111.36 -180.685 111.68 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 112.715 241.32 113.045 242.45 ;
        RECT 112.715 239.195 113.045 239.525 ;
        RECT 112.715 237.835 113.045 238.165 ;
        RECT 112.72 237.16 113.04 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 112.715 -95.365 113.045 -95.035 ;
        RECT 112.715 -96.725 113.045 -96.395 ;
        RECT 112.715 -98.085 113.045 -97.755 ;
        RECT 112.715 -99.445 113.045 -99.115 ;
        RECT 112.715 -100.805 113.045 -100.475 ;
        RECT 112.715 -102.165 113.045 -101.835 ;
        RECT 112.715 -103.525 113.045 -103.195 ;
        RECT 112.715 -104.885 113.045 -104.555 ;
        RECT 112.715 -106.245 113.045 -105.915 ;
        RECT 112.715 -107.605 113.045 -107.275 ;
        RECT 112.715 -108.965 113.045 -108.635 ;
        RECT 112.715 -110.325 113.045 -109.995 ;
        RECT 112.715 -111.685 113.045 -111.355 ;
        RECT 112.715 -113.045 113.045 -112.715 ;
        RECT 112.715 -114.405 113.045 -114.075 ;
        RECT 112.715 -115.765 113.045 -115.435 ;
        RECT 112.715 -117.125 113.045 -116.795 ;
        RECT 112.715 -118.485 113.045 -118.155 ;
        RECT 112.715 -119.845 113.045 -119.515 ;
        RECT 112.715 -121.205 113.045 -120.875 ;
        RECT 112.715 -122.565 113.045 -122.235 ;
        RECT 112.715 -123.925 113.045 -123.595 ;
        RECT 112.715 -125.285 113.045 -124.955 ;
        RECT 112.715 -126.645 113.045 -126.315 ;
        RECT 112.715 -128.005 113.045 -127.675 ;
        RECT 112.715 -129.365 113.045 -129.035 ;
        RECT 112.715 -130.725 113.045 -130.395 ;
        RECT 112.715 -132.085 113.045 -131.755 ;
        RECT 112.715 -133.445 113.045 -133.115 ;
        RECT 112.715 -134.805 113.045 -134.475 ;
        RECT 112.715 -136.165 113.045 -135.835 ;
        RECT 112.715 -137.525 113.045 -137.195 ;
        RECT 112.715 -138.885 113.045 -138.555 ;
        RECT 112.715 -140.245 113.045 -139.915 ;
        RECT 112.715 -141.605 113.045 -141.275 ;
        RECT 112.715 -142.965 113.045 -142.635 ;
        RECT 112.715 -144.325 113.045 -143.995 ;
        RECT 112.715 -145.685 113.045 -145.355 ;
        RECT 112.715 -147.045 113.045 -146.715 ;
        RECT 112.715 -148.405 113.045 -148.075 ;
        RECT 112.715 -149.765 113.045 -149.435 ;
        RECT 112.715 -151.125 113.045 -150.795 ;
        RECT 112.715 -152.485 113.045 -152.155 ;
        RECT 112.715 -153.845 113.045 -153.515 ;
        RECT 112.715 -155.205 113.045 -154.875 ;
        RECT 112.715 -156.565 113.045 -156.235 ;
        RECT 112.715 -157.925 113.045 -157.595 ;
        RECT 112.715 -159.285 113.045 -158.955 ;
        RECT 112.715 -160.645 113.045 -160.315 ;
        RECT 112.715 -162.005 113.045 -161.675 ;
        RECT 112.715 -163.365 113.045 -163.035 ;
        RECT 112.715 -164.725 113.045 -164.395 ;
        RECT 112.715 -166.085 113.045 -165.755 ;
        RECT 112.715 -167.445 113.045 -167.115 ;
        RECT 112.715 -168.805 113.045 -168.475 ;
        RECT 112.715 -170.165 113.045 -169.835 ;
        RECT 112.715 -171.525 113.045 -171.195 ;
        RECT 112.715 -172.885 113.045 -172.555 ;
        RECT 112.715 -174.245 113.045 -173.915 ;
        RECT 112.715 -175.605 113.045 -175.275 ;
        RECT 112.715 -176.965 113.045 -176.635 ;
        RECT 112.715 -178.325 113.045 -177.995 ;
        RECT 112.715 -180.57 113.045 -179.44 ;
        RECT 112.72 -180.685 113.04 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 113.11 -94.075 113.44 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 114.075 241.32 114.405 242.45 ;
        RECT 114.075 239.195 114.405 239.525 ;
        RECT 114.075 237.835 114.405 238.165 ;
        RECT 114.08 237.16 114.4 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 114.075 -1.525 114.405 -1.195 ;
        RECT 114.075 -2.885 114.405 -2.555 ;
        RECT 114.08 -3.56 114.4 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 115.435 241.32 115.765 242.45 ;
        RECT 115.435 239.195 115.765 239.525 ;
        RECT 115.435 237.835 115.765 238.165 ;
        RECT 115.44 237.16 115.76 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 115.435 -1.525 115.765 -1.195 ;
        RECT 115.435 -2.885 115.765 -2.555 ;
        RECT 115.44 -3.56 115.76 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 116.795 241.32 117.125 242.45 ;
        RECT 116.795 239.195 117.125 239.525 ;
        RECT 116.795 237.835 117.125 238.165 ;
        RECT 116.8 237.16 117.12 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 116.795 -1.525 117.125 -1.195 ;
        RECT 116.795 -2.885 117.125 -2.555 ;
        RECT 116.8 -3.56 117.12 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 116.795 -91.285 117.125 -90.955 ;
        RECT 116.795 -92.645 117.125 -92.315 ;
        RECT 116.795 -94.005 117.125 -93.675 ;
        RECT 116.795 -95.365 117.125 -95.035 ;
        RECT 116.795 -96.725 117.125 -96.395 ;
        RECT 116.795 -98.085 117.125 -97.755 ;
        RECT 116.795 -99.445 117.125 -99.115 ;
        RECT 116.795 -100.805 117.125 -100.475 ;
        RECT 116.795 -102.165 117.125 -101.835 ;
        RECT 116.795 -103.525 117.125 -103.195 ;
        RECT 116.795 -104.885 117.125 -104.555 ;
        RECT 116.795 -106.245 117.125 -105.915 ;
        RECT 116.795 -107.605 117.125 -107.275 ;
        RECT 116.795 -108.965 117.125 -108.635 ;
        RECT 116.795 -110.325 117.125 -109.995 ;
        RECT 116.795 -111.685 117.125 -111.355 ;
        RECT 116.795 -113.045 117.125 -112.715 ;
        RECT 116.795 -114.405 117.125 -114.075 ;
        RECT 116.795 -115.765 117.125 -115.435 ;
        RECT 116.795 -117.125 117.125 -116.795 ;
        RECT 116.795 -118.485 117.125 -118.155 ;
        RECT 116.795 -119.845 117.125 -119.515 ;
        RECT 116.795 -121.205 117.125 -120.875 ;
        RECT 116.795 -122.565 117.125 -122.235 ;
        RECT 116.795 -123.925 117.125 -123.595 ;
        RECT 116.795 -125.285 117.125 -124.955 ;
        RECT 116.795 -126.645 117.125 -126.315 ;
        RECT 116.795 -128.005 117.125 -127.675 ;
        RECT 116.795 -129.365 117.125 -129.035 ;
        RECT 116.795 -130.725 117.125 -130.395 ;
        RECT 116.795 -132.085 117.125 -131.755 ;
        RECT 116.795 -133.445 117.125 -133.115 ;
        RECT 116.795 -134.805 117.125 -134.475 ;
        RECT 116.795 -136.165 117.125 -135.835 ;
        RECT 116.795 -137.525 117.125 -137.195 ;
        RECT 116.795 -138.885 117.125 -138.555 ;
        RECT 116.795 -140.245 117.125 -139.915 ;
        RECT 116.795 -141.605 117.125 -141.275 ;
        RECT 116.795 -142.965 117.125 -142.635 ;
        RECT 116.795 -144.325 117.125 -143.995 ;
        RECT 116.795 -145.685 117.125 -145.355 ;
        RECT 116.795 -147.045 117.125 -146.715 ;
        RECT 116.795 -148.405 117.125 -148.075 ;
        RECT 116.795 -149.765 117.125 -149.435 ;
        RECT 116.795 -151.125 117.125 -150.795 ;
        RECT 116.795 -152.485 117.125 -152.155 ;
        RECT 116.795 -153.845 117.125 -153.515 ;
        RECT 116.795 -155.205 117.125 -154.875 ;
        RECT 116.795 -156.565 117.125 -156.235 ;
        RECT 116.795 -157.925 117.125 -157.595 ;
        RECT 116.795 -159.285 117.125 -158.955 ;
        RECT 116.795 -160.645 117.125 -160.315 ;
        RECT 116.795 -162.005 117.125 -161.675 ;
        RECT 116.795 -163.365 117.125 -163.035 ;
        RECT 116.795 -164.725 117.125 -164.395 ;
        RECT 116.795 -166.085 117.125 -165.755 ;
        RECT 116.795 -167.445 117.125 -167.115 ;
        RECT 116.795 -168.805 117.125 -168.475 ;
        RECT 116.795 -170.165 117.125 -169.835 ;
        RECT 116.795 -171.525 117.125 -171.195 ;
        RECT 116.795 -172.885 117.125 -172.555 ;
        RECT 116.795 -174.245 117.125 -173.915 ;
        RECT 116.795 -175.605 117.125 -175.275 ;
        RECT 116.795 -176.965 117.125 -176.635 ;
        RECT 116.795 -178.325 117.125 -177.995 ;
        RECT 116.795 -180.57 117.125 -179.44 ;
        RECT 116.8 -180.685 117.12 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 118.155 241.32 118.485 242.45 ;
        RECT 118.155 239.195 118.485 239.525 ;
        RECT 118.155 237.835 118.485 238.165 ;
        RECT 118.16 237.16 118.48 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 118.155 -95.365 118.485 -95.035 ;
        RECT 118.155 -96.725 118.485 -96.395 ;
        RECT 118.155 -98.085 118.485 -97.755 ;
        RECT 118.155 -99.445 118.485 -99.115 ;
        RECT 118.155 -100.805 118.485 -100.475 ;
        RECT 118.155 -102.165 118.485 -101.835 ;
        RECT 118.155 -103.525 118.485 -103.195 ;
        RECT 118.155 -104.885 118.485 -104.555 ;
        RECT 118.155 -106.245 118.485 -105.915 ;
        RECT 118.155 -107.605 118.485 -107.275 ;
        RECT 118.155 -108.965 118.485 -108.635 ;
        RECT 118.155 -110.325 118.485 -109.995 ;
        RECT 118.155 -111.685 118.485 -111.355 ;
        RECT 118.155 -113.045 118.485 -112.715 ;
        RECT 118.155 -114.405 118.485 -114.075 ;
        RECT 118.155 -115.765 118.485 -115.435 ;
        RECT 118.155 -117.125 118.485 -116.795 ;
        RECT 118.155 -118.485 118.485 -118.155 ;
        RECT 118.155 -119.845 118.485 -119.515 ;
        RECT 118.155 -121.205 118.485 -120.875 ;
        RECT 118.155 -122.565 118.485 -122.235 ;
        RECT 118.155 -123.925 118.485 -123.595 ;
        RECT 118.155 -125.285 118.485 -124.955 ;
        RECT 118.155 -126.645 118.485 -126.315 ;
        RECT 118.155 -128.005 118.485 -127.675 ;
        RECT 118.155 -129.365 118.485 -129.035 ;
        RECT 118.155 -130.725 118.485 -130.395 ;
        RECT 118.155 -132.085 118.485 -131.755 ;
        RECT 118.155 -133.445 118.485 -133.115 ;
        RECT 118.155 -134.805 118.485 -134.475 ;
        RECT 118.155 -136.165 118.485 -135.835 ;
        RECT 118.155 -137.525 118.485 -137.195 ;
        RECT 118.155 -138.885 118.485 -138.555 ;
        RECT 118.155 -140.245 118.485 -139.915 ;
        RECT 118.155 -141.605 118.485 -141.275 ;
        RECT 118.155 -142.965 118.485 -142.635 ;
        RECT 118.155 -144.325 118.485 -143.995 ;
        RECT 118.155 -145.685 118.485 -145.355 ;
        RECT 118.155 -147.045 118.485 -146.715 ;
        RECT 118.155 -148.405 118.485 -148.075 ;
        RECT 118.155 -149.765 118.485 -149.435 ;
        RECT 118.155 -151.125 118.485 -150.795 ;
        RECT 118.155 -152.485 118.485 -152.155 ;
        RECT 118.155 -153.845 118.485 -153.515 ;
        RECT 118.155 -155.205 118.485 -154.875 ;
        RECT 118.155 -156.565 118.485 -156.235 ;
        RECT 118.155 -157.925 118.485 -157.595 ;
        RECT 118.155 -159.285 118.485 -158.955 ;
        RECT 118.155 -160.645 118.485 -160.315 ;
        RECT 118.155 -162.005 118.485 -161.675 ;
        RECT 118.155 -163.365 118.485 -163.035 ;
        RECT 118.155 -164.725 118.485 -164.395 ;
        RECT 118.155 -166.085 118.485 -165.755 ;
        RECT 118.155 -167.445 118.485 -167.115 ;
        RECT 118.155 -168.805 118.485 -168.475 ;
        RECT 118.155 -170.165 118.485 -169.835 ;
        RECT 118.155 -171.525 118.485 -171.195 ;
        RECT 118.155 -172.885 118.485 -172.555 ;
        RECT 118.155 -174.245 118.485 -173.915 ;
        RECT 118.155 -175.605 118.485 -175.275 ;
        RECT 118.155 -176.965 118.485 -176.635 ;
        RECT 118.155 -178.325 118.485 -177.995 ;
        RECT 118.155 -180.57 118.485 -179.44 ;
        RECT 118.16 -180.685 118.48 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 119.21 -94.075 119.54 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 119.515 241.32 119.845 242.45 ;
        RECT 119.515 239.195 119.845 239.525 ;
        RECT 119.515 237.835 119.845 238.165 ;
        RECT 119.52 237.16 119.84 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 120.875 241.32 121.205 242.45 ;
        RECT 120.875 239.195 121.205 239.525 ;
        RECT 120.875 237.835 121.205 238.165 ;
        RECT 120.88 237.16 121.2 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 120.875 -1.525 121.205 -1.195 ;
        RECT 120.875 -2.885 121.205 -2.555 ;
        RECT 120.88 -3.56 121.2 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 122.235 241.32 122.565 242.45 ;
        RECT 122.235 239.195 122.565 239.525 ;
        RECT 122.235 237.835 122.565 238.165 ;
        RECT 122.24 237.16 122.56 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 122.235 -1.525 122.565 -1.195 ;
        RECT 122.235 -2.885 122.565 -2.555 ;
        RECT 122.24 -3.56 122.56 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 123.595 241.32 123.925 242.45 ;
        RECT 123.595 239.195 123.925 239.525 ;
        RECT 123.595 237.835 123.925 238.165 ;
        RECT 123.6 237.16 123.92 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 123.595 -1.525 123.925 -1.195 ;
        RECT 123.595 -2.885 123.925 -2.555 ;
        RECT 123.6 -3.56 123.92 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 123.595 -91.285 123.925 -90.955 ;
        RECT 123.595 -92.645 123.925 -92.315 ;
        RECT 123.595 -94.005 123.925 -93.675 ;
        RECT 123.595 -95.365 123.925 -95.035 ;
        RECT 123.595 -96.725 123.925 -96.395 ;
        RECT 123.595 -98.085 123.925 -97.755 ;
        RECT 123.595 -99.445 123.925 -99.115 ;
        RECT 123.595 -100.805 123.925 -100.475 ;
        RECT 123.595 -102.165 123.925 -101.835 ;
        RECT 123.595 -103.525 123.925 -103.195 ;
        RECT 123.595 -104.885 123.925 -104.555 ;
        RECT 123.595 -106.245 123.925 -105.915 ;
        RECT 123.595 -107.605 123.925 -107.275 ;
        RECT 123.595 -108.965 123.925 -108.635 ;
        RECT 123.595 -110.325 123.925 -109.995 ;
        RECT 123.595 -111.685 123.925 -111.355 ;
        RECT 123.595 -113.045 123.925 -112.715 ;
        RECT 123.595 -114.405 123.925 -114.075 ;
        RECT 123.595 -115.765 123.925 -115.435 ;
        RECT 123.595 -117.125 123.925 -116.795 ;
        RECT 123.595 -118.485 123.925 -118.155 ;
        RECT 123.595 -119.845 123.925 -119.515 ;
        RECT 123.595 -121.205 123.925 -120.875 ;
        RECT 123.595 -122.565 123.925 -122.235 ;
        RECT 123.595 -123.925 123.925 -123.595 ;
        RECT 123.595 -125.285 123.925 -124.955 ;
        RECT 123.595 -126.645 123.925 -126.315 ;
        RECT 123.595 -128.005 123.925 -127.675 ;
        RECT 123.595 -129.365 123.925 -129.035 ;
        RECT 123.595 -130.725 123.925 -130.395 ;
        RECT 123.595 -132.085 123.925 -131.755 ;
        RECT 123.595 -133.445 123.925 -133.115 ;
        RECT 123.595 -134.805 123.925 -134.475 ;
        RECT 123.595 -136.165 123.925 -135.835 ;
        RECT 123.595 -137.525 123.925 -137.195 ;
        RECT 123.595 -138.885 123.925 -138.555 ;
        RECT 123.595 -140.245 123.925 -139.915 ;
        RECT 123.595 -141.605 123.925 -141.275 ;
        RECT 123.595 -142.965 123.925 -142.635 ;
        RECT 123.595 -144.325 123.925 -143.995 ;
        RECT 123.595 -145.685 123.925 -145.355 ;
        RECT 123.595 -147.045 123.925 -146.715 ;
        RECT 123.595 -148.405 123.925 -148.075 ;
        RECT 123.595 -149.765 123.925 -149.435 ;
        RECT 123.595 -151.125 123.925 -150.795 ;
        RECT 123.595 -152.485 123.925 -152.155 ;
        RECT 123.595 -153.845 123.925 -153.515 ;
        RECT 123.595 -155.205 123.925 -154.875 ;
        RECT 123.595 -156.565 123.925 -156.235 ;
        RECT 123.595 -157.925 123.925 -157.595 ;
        RECT 123.595 -159.285 123.925 -158.955 ;
        RECT 123.595 -160.645 123.925 -160.315 ;
        RECT 123.595 -162.005 123.925 -161.675 ;
        RECT 123.595 -163.365 123.925 -163.035 ;
        RECT 123.595 -164.725 123.925 -164.395 ;
        RECT 123.595 -166.085 123.925 -165.755 ;
        RECT 123.595 -167.445 123.925 -167.115 ;
        RECT 123.595 -168.805 123.925 -168.475 ;
        RECT 123.595 -170.165 123.925 -169.835 ;
        RECT 123.595 -171.525 123.925 -171.195 ;
        RECT 123.595 -172.885 123.925 -172.555 ;
        RECT 123.595 -174.245 123.925 -173.915 ;
        RECT 123.595 -175.605 123.925 -175.275 ;
        RECT 123.595 -176.965 123.925 -176.635 ;
        RECT 123.595 -178.325 123.925 -177.995 ;
        RECT 123.595 -180.57 123.925 -179.44 ;
        RECT 123.6 -180.685 123.92 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 124.955 241.32 125.285 242.45 ;
        RECT 124.955 239.195 125.285 239.525 ;
        RECT 124.955 237.835 125.285 238.165 ;
        RECT 124.96 237.16 125.28 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 124.955 -95.365 125.285 -95.035 ;
        RECT 124.955 -96.725 125.285 -96.395 ;
        RECT 124.955 -98.085 125.285 -97.755 ;
        RECT 124.955 -99.445 125.285 -99.115 ;
        RECT 124.955 -100.805 125.285 -100.475 ;
        RECT 124.955 -102.165 125.285 -101.835 ;
        RECT 124.955 -103.525 125.285 -103.195 ;
        RECT 124.955 -104.885 125.285 -104.555 ;
        RECT 124.955 -106.245 125.285 -105.915 ;
        RECT 124.955 -107.605 125.285 -107.275 ;
        RECT 124.955 -108.965 125.285 -108.635 ;
        RECT 124.955 -110.325 125.285 -109.995 ;
        RECT 124.955 -111.685 125.285 -111.355 ;
        RECT 124.955 -113.045 125.285 -112.715 ;
        RECT 124.955 -114.405 125.285 -114.075 ;
        RECT 124.955 -115.765 125.285 -115.435 ;
        RECT 124.955 -117.125 125.285 -116.795 ;
        RECT 124.955 -118.485 125.285 -118.155 ;
        RECT 124.955 -119.845 125.285 -119.515 ;
        RECT 124.955 -121.205 125.285 -120.875 ;
        RECT 124.955 -122.565 125.285 -122.235 ;
        RECT 124.955 -123.925 125.285 -123.595 ;
        RECT 124.955 -125.285 125.285 -124.955 ;
        RECT 124.955 -126.645 125.285 -126.315 ;
        RECT 124.955 -128.005 125.285 -127.675 ;
        RECT 124.955 -129.365 125.285 -129.035 ;
        RECT 124.955 -130.725 125.285 -130.395 ;
        RECT 124.955 -132.085 125.285 -131.755 ;
        RECT 124.955 -133.445 125.285 -133.115 ;
        RECT 124.955 -134.805 125.285 -134.475 ;
        RECT 124.955 -136.165 125.285 -135.835 ;
        RECT 124.955 -137.525 125.285 -137.195 ;
        RECT 124.955 -138.885 125.285 -138.555 ;
        RECT 124.955 -140.245 125.285 -139.915 ;
        RECT 124.955 -141.605 125.285 -141.275 ;
        RECT 124.955 -142.965 125.285 -142.635 ;
        RECT 124.955 -144.325 125.285 -143.995 ;
        RECT 124.955 -145.685 125.285 -145.355 ;
        RECT 124.955 -147.045 125.285 -146.715 ;
        RECT 124.955 -148.405 125.285 -148.075 ;
        RECT 124.955 -149.765 125.285 -149.435 ;
        RECT 124.955 -151.125 125.285 -150.795 ;
        RECT 124.955 -152.485 125.285 -152.155 ;
        RECT 124.955 -153.845 125.285 -153.515 ;
        RECT 124.955 -155.205 125.285 -154.875 ;
        RECT 124.955 -156.565 125.285 -156.235 ;
        RECT 124.955 -157.925 125.285 -157.595 ;
        RECT 124.955 -159.285 125.285 -158.955 ;
        RECT 124.955 -160.645 125.285 -160.315 ;
        RECT 124.955 -162.005 125.285 -161.675 ;
        RECT 124.955 -163.365 125.285 -163.035 ;
        RECT 124.955 -164.725 125.285 -164.395 ;
        RECT 124.955 -166.085 125.285 -165.755 ;
        RECT 124.955 -167.445 125.285 -167.115 ;
        RECT 124.955 -168.805 125.285 -168.475 ;
        RECT 124.955 -170.165 125.285 -169.835 ;
        RECT 124.955 -171.525 125.285 -171.195 ;
        RECT 124.955 -172.885 125.285 -172.555 ;
        RECT 124.955 -174.245 125.285 -173.915 ;
        RECT 124.955 -175.605 125.285 -175.275 ;
        RECT 124.955 -176.965 125.285 -176.635 ;
        RECT 124.955 -178.325 125.285 -177.995 ;
        RECT 124.955 -180.57 125.285 -179.44 ;
        RECT 124.96 -180.685 125.28 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 125.31 -94.075 125.64 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 126.315 241.32 126.645 242.45 ;
        RECT 126.315 239.195 126.645 239.525 ;
        RECT 126.315 237.835 126.645 238.165 ;
        RECT 126.32 237.16 126.64 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 126.315 -1.525 126.645 -1.195 ;
        RECT 126.315 -2.885 126.645 -2.555 ;
        RECT 126.32 -3.56 126.64 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 127.675 241.32 128.005 242.45 ;
        RECT 127.675 239.195 128.005 239.525 ;
        RECT 127.675 237.835 128.005 238.165 ;
        RECT 127.68 237.16 128 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 127.675 -1.525 128.005 -1.195 ;
        RECT 127.675 -2.885 128.005 -2.555 ;
        RECT 127.68 -3.56 128 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.035 241.32 129.365 242.45 ;
        RECT 129.035 239.195 129.365 239.525 ;
        RECT 129.035 237.835 129.365 238.165 ;
        RECT 129.04 237.16 129.36 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.035 -1.525 129.365 -1.195 ;
        RECT 129.035 -2.885 129.365 -2.555 ;
        RECT 129.04 -3.56 129.36 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.035 -91.285 129.365 -90.955 ;
        RECT 129.035 -92.645 129.365 -92.315 ;
        RECT 129.035 -94.005 129.365 -93.675 ;
        RECT 129.035 -95.365 129.365 -95.035 ;
        RECT 129.035 -96.725 129.365 -96.395 ;
        RECT 129.035 -98.085 129.365 -97.755 ;
        RECT 129.035 -99.445 129.365 -99.115 ;
        RECT 129.035 -100.805 129.365 -100.475 ;
        RECT 129.035 -102.165 129.365 -101.835 ;
        RECT 129.035 -103.525 129.365 -103.195 ;
        RECT 129.035 -104.885 129.365 -104.555 ;
        RECT 129.035 -106.245 129.365 -105.915 ;
        RECT 129.035 -107.605 129.365 -107.275 ;
        RECT 129.035 -108.965 129.365 -108.635 ;
        RECT 129.035 -110.325 129.365 -109.995 ;
        RECT 129.035 -111.685 129.365 -111.355 ;
        RECT 129.035 -113.045 129.365 -112.715 ;
        RECT 129.035 -114.405 129.365 -114.075 ;
        RECT 129.035 -115.765 129.365 -115.435 ;
        RECT 129.035 -117.125 129.365 -116.795 ;
        RECT 129.035 -118.485 129.365 -118.155 ;
        RECT 129.035 -119.845 129.365 -119.515 ;
        RECT 129.035 -121.205 129.365 -120.875 ;
        RECT 129.035 -122.565 129.365 -122.235 ;
        RECT 129.035 -123.925 129.365 -123.595 ;
        RECT 129.035 -125.285 129.365 -124.955 ;
        RECT 129.035 -126.645 129.365 -126.315 ;
        RECT 129.035 -128.005 129.365 -127.675 ;
        RECT 129.035 -129.365 129.365 -129.035 ;
        RECT 129.035 -130.725 129.365 -130.395 ;
        RECT 129.035 -132.085 129.365 -131.755 ;
        RECT 129.035 -133.445 129.365 -133.115 ;
        RECT 129.035 -134.805 129.365 -134.475 ;
        RECT 129.035 -136.165 129.365 -135.835 ;
        RECT 129.035 -137.525 129.365 -137.195 ;
        RECT 129.035 -138.885 129.365 -138.555 ;
        RECT 129.035 -140.245 129.365 -139.915 ;
        RECT 129.035 -141.605 129.365 -141.275 ;
        RECT 129.035 -142.965 129.365 -142.635 ;
        RECT 129.035 -144.325 129.365 -143.995 ;
        RECT 129.035 -145.685 129.365 -145.355 ;
        RECT 129.035 -147.045 129.365 -146.715 ;
        RECT 129.035 -148.405 129.365 -148.075 ;
        RECT 129.035 -149.765 129.365 -149.435 ;
        RECT 129.035 -151.125 129.365 -150.795 ;
        RECT 129.035 -152.485 129.365 -152.155 ;
        RECT 129.035 -153.845 129.365 -153.515 ;
        RECT 129.035 -155.205 129.365 -154.875 ;
        RECT 129.035 -156.565 129.365 -156.235 ;
        RECT 129.035 -157.925 129.365 -157.595 ;
        RECT 129.035 -159.285 129.365 -158.955 ;
        RECT 129.035 -160.645 129.365 -160.315 ;
        RECT 129.035 -162.005 129.365 -161.675 ;
        RECT 129.035 -163.365 129.365 -163.035 ;
        RECT 129.035 -164.725 129.365 -164.395 ;
        RECT 129.035 -166.085 129.365 -165.755 ;
        RECT 129.035 -167.445 129.365 -167.115 ;
        RECT 129.035 -168.805 129.365 -168.475 ;
        RECT 129.035 -170.165 129.365 -169.835 ;
        RECT 129.035 -171.525 129.365 -171.195 ;
        RECT 129.035 -172.885 129.365 -172.555 ;
        RECT 129.035 -174.245 129.365 -173.915 ;
        RECT 129.035 -175.605 129.365 -175.275 ;
        RECT 129.035 -176.965 129.365 -176.635 ;
        RECT 129.035 -178.325 129.365 -177.995 ;
        RECT 129.035 -180.57 129.365 -179.44 ;
        RECT 129.04 -180.685 129.36 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 130.395 241.32 130.725 242.45 ;
        RECT 130.395 239.195 130.725 239.525 ;
        RECT 130.395 237.835 130.725 238.165 ;
        RECT 130.4 237.16 130.72 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 130.395 -95.365 130.725 -95.035 ;
        RECT 130.395 -96.725 130.725 -96.395 ;
        RECT 130.395 -98.085 130.725 -97.755 ;
        RECT 130.395 -99.445 130.725 -99.115 ;
        RECT 130.395 -100.805 130.725 -100.475 ;
        RECT 130.395 -102.165 130.725 -101.835 ;
        RECT 130.395 -103.525 130.725 -103.195 ;
        RECT 130.395 -104.885 130.725 -104.555 ;
        RECT 130.395 -106.245 130.725 -105.915 ;
        RECT 130.395 -107.605 130.725 -107.275 ;
        RECT 130.395 -108.965 130.725 -108.635 ;
        RECT 130.395 -110.325 130.725 -109.995 ;
        RECT 130.395 -111.685 130.725 -111.355 ;
        RECT 130.395 -113.045 130.725 -112.715 ;
        RECT 130.395 -114.405 130.725 -114.075 ;
        RECT 130.395 -115.765 130.725 -115.435 ;
        RECT 130.395 -117.125 130.725 -116.795 ;
        RECT 130.395 -118.485 130.725 -118.155 ;
        RECT 130.395 -119.845 130.725 -119.515 ;
        RECT 130.395 -121.205 130.725 -120.875 ;
        RECT 130.395 -122.565 130.725 -122.235 ;
        RECT 130.395 -123.925 130.725 -123.595 ;
        RECT 130.395 -125.285 130.725 -124.955 ;
        RECT 130.395 -126.645 130.725 -126.315 ;
        RECT 130.395 -128.005 130.725 -127.675 ;
        RECT 130.395 -129.365 130.725 -129.035 ;
        RECT 130.395 -130.725 130.725 -130.395 ;
        RECT 130.395 -132.085 130.725 -131.755 ;
        RECT 130.395 -133.445 130.725 -133.115 ;
        RECT 130.395 -134.805 130.725 -134.475 ;
        RECT 130.395 -136.165 130.725 -135.835 ;
        RECT 130.395 -137.525 130.725 -137.195 ;
        RECT 130.395 -138.885 130.725 -138.555 ;
        RECT 130.395 -140.245 130.725 -139.915 ;
        RECT 130.395 -141.605 130.725 -141.275 ;
        RECT 130.395 -142.965 130.725 -142.635 ;
        RECT 130.395 -144.325 130.725 -143.995 ;
        RECT 130.395 -145.685 130.725 -145.355 ;
        RECT 130.395 -147.045 130.725 -146.715 ;
        RECT 130.395 -148.405 130.725 -148.075 ;
        RECT 130.395 -149.765 130.725 -149.435 ;
        RECT 130.395 -151.125 130.725 -150.795 ;
        RECT 130.395 -152.485 130.725 -152.155 ;
        RECT 130.395 -153.845 130.725 -153.515 ;
        RECT 130.395 -155.205 130.725 -154.875 ;
        RECT 130.395 -156.565 130.725 -156.235 ;
        RECT 130.395 -157.925 130.725 -157.595 ;
        RECT 130.395 -159.285 130.725 -158.955 ;
        RECT 130.395 -160.645 130.725 -160.315 ;
        RECT 130.395 -162.005 130.725 -161.675 ;
        RECT 130.395 -163.365 130.725 -163.035 ;
        RECT 130.395 -164.725 130.725 -164.395 ;
        RECT 130.395 -166.085 130.725 -165.755 ;
        RECT 130.395 -167.445 130.725 -167.115 ;
        RECT 130.395 -168.805 130.725 -168.475 ;
        RECT 130.395 -170.165 130.725 -169.835 ;
        RECT 130.395 -171.525 130.725 -171.195 ;
        RECT 130.395 -172.885 130.725 -172.555 ;
        RECT 130.395 -174.245 130.725 -173.915 ;
        RECT 130.395 -175.605 130.725 -175.275 ;
        RECT 130.395 -176.965 130.725 -176.635 ;
        RECT 130.395 -178.325 130.725 -177.995 ;
        RECT 130.395 -180.57 130.725 -179.44 ;
        RECT 130.4 -180.685 130.72 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 131.41 -94.075 131.74 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 131.755 241.32 132.085 242.45 ;
        RECT 131.755 239.195 132.085 239.525 ;
        RECT 131.755 237.835 132.085 238.165 ;
        RECT 131.76 237.16 132.08 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 133.115 241.32 133.445 242.45 ;
        RECT 133.115 239.195 133.445 239.525 ;
        RECT 133.115 237.835 133.445 238.165 ;
        RECT 133.12 237.16 133.44 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 133.115 -1.525 133.445 -1.195 ;
        RECT 133.115 -2.885 133.445 -2.555 ;
        RECT 133.12 -3.56 133.44 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 134.475 241.32 134.805 242.45 ;
        RECT 134.475 239.195 134.805 239.525 ;
        RECT 134.475 237.835 134.805 238.165 ;
        RECT 134.48 237.16 134.8 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 134.475 -1.525 134.805 -1.195 ;
        RECT 134.475 -2.885 134.805 -2.555 ;
        RECT 134.48 -3.56 134.8 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 134.475 -91.285 134.805 -90.955 ;
        RECT 134.475 -92.645 134.805 -92.315 ;
        RECT 134.475 -94.005 134.805 -93.675 ;
        RECT 134.475 -95.365 134.805 -95.035 ;
        RECT 134.475 -96.725 134.805 -96.395 ;
        RECT 134.475 -98.085 134.805 -97.755 ;
        RECT 134.475 -99.445 134.805 -99.115 ;
        RECT 134.475 -100.805 134.805 -100.475 ;
        RECT 134.475 -102.165 134.805 -101.835 ;
        RECT 134.475 -103.525 134.805 -103.195 ;
        RECT 134.475 -104.885 134.805 -104.555 ;
        RECT 134.475 -106.245 134.805 -105.915 ;
        RECT 134.475 -107.605 134.805 -107.275 ;
        RECT 134.475 -108.965 134.805 -108.635 ;
        RECT 134.475 -110.325 134.805 -109.995 ;
        RECT 134.475 -111.685 134.805 -111.355 ;
        RECT 134.475 -113.045 134.805 -112.715 ;
        RECT 134.475 -114.405 134.805 -114.075 ;
        RECT 134.475 -115.765 134.805 -115.435 ;
        RECT 134.475 -117.125 134.805 -116.795 ;
        RECT 134.475 -118.485 134.805 -118.155 ;
        RECT 134.475 -119.845 134.805 -119.515 ;
        RECT 134.475 -121.205 134.805 -120.875 ;
        RECT 134.475 -122.565 134.805 -122.235 ;
        RECT 134.475 -123.925 134.805 -123.595 ;
        RECT 134.475 -125.285 134.805 -124.955 ;
        RECT 134.475 -126.645 134.805 -126.315 ;
        RECT 134.475 -128.005 134.805 -127.675 ;
        RECT 134.475 -129.365 134.805 -129.035 ;
        RECT 134.475 -130.725 134.805 -130.395 ;
        RECT 134.475 -132.085 134.805 -131.755 ;
        RECT 134.475 -133.445 134.805 -133.115 ;
        RECT 134.475 -134.805 134.805 -134.475 ;
        RECT 134.475 -136.165 134.805 -135.835 ;
        RECT 134.475 -137.525 134.805 -137.195 ;
        RECT 134.475 -138.885 134.805 -138.555 ;
        RECT 134.475 -140.245 134.805 -139.915 ;
        RECT 134.475 -141.605 134.805 -141.275 ;
        RECT 134.475 -142.965 134.805 -142.635 ;
        RECT 134.475 -144.325 134.805 -143.995 ;
        RECT 134.475 -145.685 134.805 -145.355 ;
        RECT 134.475 -147.045 134.805 -146.715 ;
        RECT 134.475 -148.405 134.805 -148.075 ;
        RECT 134.475 -149.765 134.805 -149.435 ;
        RECT 134.475 -151.125 134.805 -150.795 ;
        RECT 134.475 -152.485 134.805 -152.155 ;
        RECT 134.475 -153.845 134.805 -153.515 ;
        RECT 134.475 -155.205 134.805 -154.875 ;
        RECT 134.475 -156.565 134.805 -156.235 ;
        RECT 134.475 -157.925 134.805 -157.595 ;
        RECT 134.475 -159.285 134.805 -158.955 ;
        RECT 134.475 -160.645 134.805 -160.315 ;
        RECT 134.475 -162.005 134.805 -161.675 ;
        RECT 134.475 -163.365 134.805 -163.035 ;
        RECT 134.475 -164.725 134.805 -164.395 ;
        RECT 134.475 -166.085 134.805 -165.755 ;
        RECT 134.475 -167.445 134.805 -167.115 ;
        RECT 134.475 -168.805 134.805 -168.475 ;
        RECT 134.475 -170.165 134.805 -169.835 ;
        RECT 134.475 -171.525 134.805 -171.195 ;
        RECT 134.475 -172.885 134.805 -172.555 ;
        RECT 134.475 -174.245 134.805 -173.915 ;
        RECT 134.475 -175.605 134.805 -175.275 ;
        RECT 134.475 -176.965 134.805 -176.635 ;
        RECT 134.475 -178.325 134.805 -177.995 ;
        RECT 134.475 -180.57 134.805 -179.44 ;
        RECT 134.48 -180.685 134.8 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 135.835 241.32 136.165 242.45 ;
        RECT 135.835 239.195 136.165 239.525 ;
        RECT 135.835 237.835 136.165 238.165 ;
        RECT 135.84 237.16 136.16 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 135.835 -1.525 136.165 -1.195 ;
        RECT 135.835 -2.885 136.165 -2.555 ;
        RECT 135.84 -3.56 136.16 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 135.835 -91.285 136.165 -90.955 ;
        RECT 135.835 -92.645 136.165 -92.315 ;
        RECT 135.835 -94.005 136.165 -93.675 ;
        RECT 135.835 -95.365 136.165 -95.035 ;
        RECT 135.835 -96.725 136.165 -96.395 ;
        RECT 135.835 -98.085 136.165 -97.755 ;
        RECT 135.835 -99.445 136.165 -99.115 ;
        RECT 135.835 -100.805 136.165 -100.475 ;
        RECT 135.835 -102.165 136.165 -101.835 ;
        RECT 135.835 -103.525 136.165 -103.195 ;
        RECT 135.835 -104.885 136.165 -104.555 ;
        RECT 135.835 -106.245 136.165 -105.915 ;
        RECT 135.835 -107.605 136.165 -107.275 ;
        RECT 135.835 -108.965 136.165 -108.635 ;
        RECT 135.835 -110.325 136.165 -109.995 ;
        RECT 135.835 -111.685 136.165 -111.355 ;
        RECT 135.835 -113.045 136.165 -112.715 ;
        RECT 135.835 -114.405 136.165 -114.075 ;
        RECT 135.835 -115.765 136.165 -115.435 ;
        RECT 135.835 -117.125 136.165 -116.795 ;
        RECT 135.835 -118.485 136.165 -118.155 ;
        RECT 135.835 -119.845 136.165 -119.515 ;
        RECT 135.835 -121.205 136.165 -120.875 ;
        RECT 135.835 -122.565 136.165 -122.235 ;
        RECT 135.835 -123.925 136.165 -123.595 ;
        RECT 135.835 -125.285 136.165 -124.955 ;
        RECT 135.835 -126.645 136.165 -126.315 ;
        RECT 135.835 -128.005 136.165 -127.675 ;
        RECT 135.835 -129.365 136.165 -129.035 ;
        RECT 135.835 -130.725 136.165 -130.395 ;
        RECT 135.835 -132.085 136.165 -131.755 ;
        RECT 135.835 -133.445 136.165 -133.115 ;
        RECT 135.835 -134.805 136.165 -134.475 ;
        RECT 135.835 -136.165 136.165 -135.835 ;
        RECT 135.835 -137.525 136.165 -137.195 ;
        RECT 135.835 -138.885 136.165 -138.555 ;
        RECT 135.835 -140.245 136.165 -139.915 ;
        RECT 135.835 -141.605 136.165 -141.275 ;
        RECT 135.835 -142.965 136.165 -142.635 ;
        RECT 135.835 -144.325 136.165 -143.995 ;
        RECT 135.835 -145.685 136.165 -145.355 ;
        RECT 135.835 -147.045 136.165 -146.715 ;
        RECT 135.835 -148.405 136.165 -148.075 ;
        RECT 135.835 -149.765 136.165 -149.435 ;
        RECT 135.835 -151.125 136.165 -150.795 ;
        RECT 135.835 -152.485 136.165 -152.155 ;
        RECT 135.835 -153.845 136.165 -153.515 ;
        RECT 135.835 -155.205 136.165 -154.875 ;
        RECT 135.835 -156.565 136.165 -156.235 ;
        RECT 135.835 -157.925 136.165 -157.595 ;
        RECT 135.835 -159.285 136.165 -158.955 ;
        RECT 135.835 -160.645 136.165 -160.315 ;
        RECT 135.835 -162.005 136.165 -161.675 ;
        RECT 135.835 -163.365 136.165 -163.035 ;
        RECT 135.835 -164.725 136.165 -164.395 ;
        RECT 135.835 -166.085 136.165 -165.755 ;
        RECT 135.835 -167.445 136.165 -167.115 ;
        RECT 135.835 -168.805 136.165 -168.475 ;
        RECT 135.835 -170.165 136.165 -169.835 ;
        RECT 135.835 -171.525 136.165 -171.195 ;
        RECT 135.835 -172.885 136.165 -172.555 ;
        RECT 135.835 -174.245 136.165 -173.915 ;
        RECT 135.835 -175.605 136.165 -175.275 ;
        RECT 135.835 -176.965 136.165 -176.635 ;
        RECT 135.835 -178.325 136.165 -177.995 ;
        RECT 135.835 -180.57 136.165 -179.44 ;
        RECT 135.84 -180.685 136.16 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 137.195 241.32 137.525 242.45 ;
        RECT 137.195 239.195 137.525 239.525 ;
        RECT 137.195 237.835 137.525 238.165 ;
        RECT 137.2 237.16 137.52 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 137.195 -157.925 137.525 -157.595 ;
        RECT 137.195 -159.285 137.525 -158.955 ;
        RECT 137.195 -160.645 137.525 -160.315 ;
        RECT 137.195 -162.005 137.525 -161.675 ;
        RECT 137.195 -163.365 137.525 -163.035 ;
        RECT 137.195 -164.725 137.525 -164.395 ;
        RECT 137.195 -166.085 137.525 -165.755 ;
        RECT 137.195 -167.445 137.525 -167.115 ;
        RECT 137.195 -168.805 137.525 -168.475 ;
        RECT 137.195 -170.165 137.525 -169.835 ;
        RECT 137.195 -171.525 137.525 -171.195 ;
        RECT 137.195 -172.885 137.525 -172.555 ;
        RECT 137.195 -174.245 137.525 -173.915 ;
        RECT 137.195 -175.605 137.525 -175.275 ;
        RECT 137.195 -176.965 137.525 -176.635 ;
        RECT 137.195 -178.325 137.525 -177.995 ;
        RECT 137.195 -180.57 137.525 -179.44 ;
        RECT 137.2 -180.685 137.52 -95.035 ;
        RECT 137.195 -95.365 137.525 -95.035 ;
        RECT 137.195 -96.725 137.525 -96.395 ;
        RECT 137.195 -98.085 137.525 -97.755 ;
        RECT 137.195 -99.445 137.525 -99.115 ;
        RECT 137.195 -100.805 137.525 -100.475 ;
        RECT 137.195 -102.165 137.525 -101.835 ;
        RECT 137.195 -103.525 137.525 -103.195 ;
        RECT 137.195 -104.885 137.525 -104.555 ;
        RECT 137.195 -106.245 137.525 -105.915 ;
        RECT 137.195 -107.605 137.525 -107.275 ;
        RECT 137.195 -108.965 137.525 -108.635 ;
        RECT 137.195 -110.325 137.525 -109.995 ;
        RECT 137.195 -111.685 137.525 -111.355 ;
        RECT 137.195 -113.045 137.525 -112.715 ;
        RECT 137.195 -114.405 137.525 -114.075 ;
        RECT 137.195 -115.765 137.525 -115.435 ;
        RECT 137.195 -117.125 137.525 -116.795 ;
        RECT 137.195 -118.485 137.525 -118.155 ;
        RECT 137.195 -119.845 137.525 -119.515 ;
        RECT 137.195 -121.205 137.525 -120.875 ;
        RECT 137.195 -122.565 137.525 -122.235 ;
        RECT 137.195 -123.925 137.525 -123.595 ;
        RECT 137.195 -125.285 137.525 -124.955 ;
        RECT 137.195 -126.645 137.525 -126.315 ;
        RECT 137.195 -128.005 137.525 -127.675 ;
        RECT 137.195 -129.365 137.525 -129.035 ;
        RECT 137.195 -130.725 137.525 -130.395 ;
        RECT 137.195 -132.085 137.525 -131.755 ;
        RECT 137.195 -133.445 137.525 -133.115 ;
        RECT 137.195 -134.805 137.525 -134.475 ;
        RECT 137.195 -136.165 137.525 -135.835 ;
        RECT 137.195 -137.525 137.525 -137.195 ;
        RECT 137.195 -138.885 137.525 -138.555 ;
        RECT 137.195 -140.245 137.525 -139.915 ;
        RECT 137.195 -141.605 137.525 -141.275 ;
        RECT 137.195 -142.965 137.525 -142.635 ;
        RECT 137.195 -144.325 137.525 -143.995 ;
        RECT 137.195 -145.685 137.525 -145.355 ;
        RECT 137.195 -147.045 137.525 -146.715 ;
        RECT 137.195 -148.405 137.525 -148.075 ;
        RECT 137.195 -149.765 137.525 -149.435 ;
        RECT 137.195 -151.125 137.525 -150.795 ;
        RECT 137.195 -152.485 137.525 -152.155 ;
        RECT 137.195 -153.845 137.525 -153.515 ;
        RECT 137.195 -155.205 137.525 -154.875 ;
        RECT 137.195 -156.565 137.525 -156.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.195 241.32 69.525 242.45 ;
        RECT 69.195 239.195 69.525 239.525 ;
        RECT 69.195 237.835 69.525 238.165 ;
        RECT 69.2 237.16 69.52 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.195 -95.365 69.525 -95.035 ;
        RECT 69.195 -96.725 69.525 -96.395 ;
        RECT 69.195 -98.085 69.525 -97.755 ;
        RECT 69.195 -99.445 69.525 -99.115 ;
        RECT 69.195 -100.805 69.525 -100.475 ;
        RECT 69.195 -102.165 69.525 -101.835 ;
        RECT 69.195 -103.525 69.525 -103.195 ;
        RECT 69.195 -104.885 69.525 -104.555 ;
        RECT 69.195 -106.245 69.525 -105.915 ;
        RECT 69.195 -107.605 69.525 -107.275 ;
        RECT 69.195 -108.965 69.525 -108.635 ;
        RECT 69.195 -110.325 69.525 -109.995 ;
        RECT 69.195 -111.685 69.525 -111.355 ;
        RECT 69.195 -113.045 69.525 -112.715 ;
        RECT 69.195 -114.405 69.525 -114.075 ;
        RECT 69.195 -115.765 69.525 -115.435 ;
        RECT 69.195 -117.125 69.525 -116.795 ;
        RECT 69.195 -118.485 69.525 -118.155 ;
        RECT 69.195 -119.845 69.525 -119.515 ;
        RECT 69.195 -121.205 69.525 -120.875 ;
        RECT 69.195 -122.565 69.525 -122.235 ;
        RECT 69.195 -123.925 69.525 -123.595 ;
        RECT 69.195 -125.285 69.525 -124.955 ;
        RECT 69.195 -126.645 69.525 -126.315 ;
        RECT 69.195 -128.005 69.525 -127.675 ;
        RECT 69.195 -129.365 69.525 -129.035 ;
        RECT 69.195 -130.725 69.525 -130.395 ;
        RECT 69.195 -132.085 69.525 -131.755 ;
        RECT 69.195 -133.445 69.525 -133.115 ;
        RECT 69.195 -134.805 69.525 -134.475 ;
        RECT 69.195 -136.165 69.525 -135.835 ;
        RECT 69.195 -137.525 69.525 -137.195 ;
        RECT 69.195 -138.885 69.525 -138.555 ;
        RECT 69.195 -140.245 69.525 -139.915 ;
        RECT 69.195 -141.605 69.525 -141.275 ;
        RECT 69.195 -142.965 69.525 -142.635 ;
        RECT 69.195 -144.325 69.525 -143.995 ;
        RECT 69.195 -145.685 69.525 -145.355 ;
        RECT 69.195 -147.045 69.525 -146.715 ;
        RECT 69.195 -148.405 69.525 -148.075 ;
        RECT 69.195 -149.765 69.525 -149.435 ;
        RECT 69.195 -151.125 69.525 -150.795 ;
        RECT 69.195 -152.485 69.525 -152.155 ;
        RECT 69.195 -153.845 69.525 -153.515 ;
        RECT 69.195 -155.205 69.525 -154.875 ;
        RECT 69.195 -156.565 69.525 -156.235 ;
        RECT 69.195 -157.925 69.525 -157.595 ;
        RECT 69.195 -159.285 69.525 -158.955 ;
        RECT 69.195 -160.645 69.525 -160.315 ;
        RECT 69.195 -162.005 69.525 -161.675 ;
        RECT 69.195 -163.365 69.525 -163.035 ;
        RECT 69.195 -164.725 69.525 -164.395 ;
        RECT 69.195 -166.085 69.525 -165.755 ;
        RECT 69.195 -167.445 69.525 -167.115 ;
        RECT 69.195 -168.805 69.525 -168.475 ;
        RECT 69.195 -170.165 69.525 -169.835 ;
        RECT 69.195 -171.525 69.525 -171.195 ;
        RECT 69.195 -172.885 69.525 -172.555 ;
        RECT 69.195 -174.245 69.525 -173.915 ;
        RECT 69.195 -175.605 69.525 -175.275 ;
        RECT 69.195 -176.965 69.525 -176.635 ;
        RECT 69.195 -178.325 69.525 -177.995 ;
        RECT 69.195 -180.57 69.525 -179.44 ;
        RECT 69.2 -180.685 69.52 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.41 -94.075 70.74 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.555 241.32 70.885 242.45 ;
        RECT 70.555 239.195 70.885 239.525 ;
        RECT 70.555 237.835 70.885 238.165 ;
        RECT 70.56 237.16 70.88 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915 241.32 72.245 242.45 ;
        RECT 71.915 239.195 72.245 239.525 ;
        RECT 71.915 237.835 72.245 238.165 ;
        RECT 71.92 237.16 72.24 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915 -1.525 72.245 -1.195 ;
        RECT 71.915 -2.885 72.245 -2.555 ;
        RECT 71.92 -3.56 72.24 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915 -91.285 72.245 -90.955 ;
        RECT 71.915 -92.645 72.245 -92.315 ;
        RECT 71.915 -94.005 72.245 -93.675 ;
        RECT 71.915 -95.365 72.245 -95.035 ;
        RECT 71.915 -96.725 72.245 -96.395 ;
        RECT 71.915 -98.085 72.245 -97.755 ;
        RECT 71.915 -99.445 72.245 -99.115 ;
        RECT 71.915 -100.805 72.245 -100.475 ;
        RECT 71.915 -102.165 72.245 -101.835 ;
        RECT 71.915 -103.525 72.245 -103.195 ;
        RECT 71.915 -104.885 72.245 -104.555 ;
        RECT 71.915 -106.245 72.245 -105.915 ;
        RECT 71.915 -107.605 72.245 -107.275 ;
        RECT 71.915 -108.965 72.245 -108.635 ;
        RECT 71.915 -110.325 72.245 -109.995 ;
        RECT 71.915 -111.685 72.245 -111.355 ;
        RECT 71.915 -113.045 72.245 -112.715 ;
        RECT 71.915 -114.405 72.245 -114.075 ;
        RECT 71.915 -115.765 72.245 -115.435 ;
        RECT 71.915 -117.125 72.245 -116.795 ;
        RECT 71.915 -118.485 72.245 -118.155 ;
        RECT 71.915 -119.845 72.245 -119.515 ;
        RECT 71.915 -121.205 72.245 -120.875 ;
        RECT 71.915 -122.565 72.245 -122.235 ;
        RECT 71.915 -123.925 72.245 -123.595 ;
        RECT 71.915 -125.285 72.245 -124.955 ;
        RECT 71.915 -126.645 72.245 -126.315 ;
        RECT 71.915 -128.005 72.245 -127.675 ;
        RECT 71.915 -129.365 72.245 -129.035 ;
        RECT 71.915 -130.725 72.245 -130.395 ;
        RECT 71.915 -132.085 72.245 -131.755 ;
        RECT 71.915 -133.445 72.245 -133.115 ;
        RECT 71.915 -134.805 72.245 -134.475 ;
        RECT 71.915 -136.165 72.245 -135.835 ;
        RECT 71.915 -137.525 72.245 -137.195 ;
        RECT 71.915 -138.885 72.245 -138.555 ;
        RECT 71.915 -140.245 72.245 -139.915 ;
        RECT 71.915 -141.605 72.245 -141.275 ;
        RECT 71.915 -142.965 72.245 -142.635 ;
        RECT 71.915 -144.325 72.245 -143.995 ;
        RECT 71.915 -145.685 72.245 -145.355 ;
        RECT 71.915 -147.045 72.245 -146.715 ;
        RECT 71.915 -148.405 72.245 -148.075 ;
        RECT 71.915 -149.765 72.245 -149.435 ;
        RECT 71.915 -151.125 72.245 -150.795 ;
        RECT 71.915 -152.485 72.245 -152.155 ;
        RECT 71.915 -153.845 72.245 -153.515 ;
        RECT 71.915 -155.205 72.245 -154.875 ;
        RECT 71.915 -156.565 72.245 -156.235 ;
        RECT 71.915 -157.925 72.245 -157.595 ;
        RECT 71.915 -159.285 72.245 -158.955 ;
        RECT 71.915 -160.645 72.245 -160.315 ;
        RECT 71.915 -162.005 72.245 -161.675 ;
        RECT 71.915 -163.365 72.245 -163.035 ;
        RECT 71.915 -164.725 72.245 -164.395 ;
        RECT 71.915 -166.085 72.245 -165.755 ;
        RECT 71.915 -167.445 72.245 -167.115 ;
        RECT 71.915 -168.805 72.245 -168.475 ;
        RECT 71.915 -170.165 72.245 -169.835 ;
        RECT 71.915 -171.525 72.245 -171.195 ;
        RECT 71.915 -172.885 72.245 -172.555 ;
        RECT 71.915 -174.245 72.245 -173.915 ;
        RECT 71.915 -175.605 72.245 -175.275 ;
        RECT 71.915 -176.965 72.245 -176.635 ;
        RECT 71.915 -178.325 72.245 -177.995 ;
        RECT 71.915 -180.57 72.245 -179.44 ;
        RECT 71.92 -180.685 72.24 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.275 241.32 73.605 242.45 ;
        RECT 73.275 239.195 73.605 239.525 ;
        RECT 73.275 237.835 73.605 238.165 ;
        RECT 73.28 237.16 73.6 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.275 -1.525 73.605 -1.195 ;
        RECT 73.275 -2.885 73.605 -2.555 ;
        RECT 73.28 -3.56 73.6 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.635 241.32 74.965 242.45 ;
        RECT 74.635 239.195 74.965 239.525 ;
        RECT 74.635 237.835 74.965 238.165 ;
        RECT 74.64 237.16 74.96 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.635 -1.525 74.965 -1.195 ;
        RECT 74.635 -2.885 74.965 -2.555 ;
        RECT 74.64 -3.56 74.96 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.635 -91.285 74.965 -90.955 ;
        RECT 74.635 -92.645 74.965 -92.315 ;
        RECT 74.635 -94.005 74.965 -93.675 ;
        RECT 74.635 -95.365 74.965 -95.035 ;
        RECT 74.635 -96.725 74.965 -96.395 ;
        RECT 74.635 -98.085 74.965 -97.755 ;
        RECT 74.635 -99.445 74.965 -99.115 ;
        RECT 74.635 -100.805 74.965 -100.475 ;
        RECT 74.635 -102.165 74.965 -101.835 ;
        RECT 74.635 -103.525 74.965 -103.195 ;
        RECT 74.635 -104.885 74.965 -104.555 ;
        RECT 74.635 -106.245 74.965 -105.915 ;
        RECT 74.635 -107.605 74.965 -107.275 ;
        RECT 74.635 -108.965 74.965 -108.635 ;
        RECT 74.635 -110.325 74.965 -109.995 ;
        RECT 74.635 -111.685 74.965 -111.355 ;
        RECT 74.635 -113.045 74.965 -112.715 ;
        RECT 74.635 -114.405 74.965 -114.075 ;
        RECT 74.635 -115.765 74.965 -115.435 ;
        RECT 74.635 -117.125 74.965 -116.795 ;
        RECT 74.635 -118.485 74.965 -118.155 ;
        RECT 74.635 -119.845 74.965 -119.515 ;
        RECT 74.635 -121.205 74.965 -120.875 ;
        RECT 74.635 -122.565 74.965 -122.235 ;
        RECT 74.635 -123.925 74.965 -123.595 ;
        RECT 74.635 -125.285 74.965 -124.955 ;
        RECT 74.635 -126.645 74.965 -126.315 ;
        RECT 74.635 -128.005 74.965 -127.675 ;
        RECT 74.635 -129.365 74.965 -129.035 ;
        RECT 74.635 -130.725 74.965 -130.395 ;
        RECT 74.635 -132.085 74.965 -131.755 ;
        RECT 74.635 -133.445 74.965 -133.115 ;
        RECT 74.635 -134.805 74.965 -134.475 ;
        RECT 74.635 -136.165 74.965 -135.835 ;
        RECT 74.635 -137.525 74.965 -137.195 ;
        RECT 74.635 -138.885 74.965 -138.555 ;
        RECT 74.635 -140.245 74.965 -139.915 ;
        RECT 74.635 -141.605 74.965 -141.275 ;
        RECT 74.635 -142.965 74.965 -142.635 ;
        RECT 74.635 -144.325 74.965 -143.995 ;
        RECT 74.635 -145.685 74.965 -145.355 ;
        RECT 74.635 -147.045 74.965 -146.715 ;
        RECT 74.635 -148.405 74.965 -148.075 ;
        RECT 74.635 -149.765 74.965 -149.435 ;
        RECT 74.635 -151.125 74.965 -150.795 ;
        RECT 74.635 -152.485 74.965 -152.155 ;
        RECT 74.635 -153.845 74.965 -153.515 ;
        RECT 74.635 -155.205 74.965 -154.875 ;
        RECT 74.635 -156.565 74.965 -156.235 ;
        RECT 74.635 -157.925 74.965 -157.595 ;
        RECT 74.635 -159.285 74.965 -158.955 ;
        RECT 74.635 -160.645 74.965 -160.315 ;
        RECT 74.635 -162.005 74.965 -161.675 ;
        RECT 74.635 -163.365 74.965 -163.035 ;
        RECT 74.635 -164.725 74.965 -164.395 ;
        RECT 74.635 -166.085 74.965 -165.755 ;
        RECT 74.635 -167.445 74.965 -167.115 ;
        RECT 74.635 -168.805 74.965 -168.475 ;
        RECT 74.635 -170.165 74.965 -169.835 ;
        RECT 74.635 -171.525 74.965 -171.195 ;
        RECT 74.635 -172.885 74.965 -172.555 ;
        RECT 74.635 -174.245 74.965 -173.915 ;
        RECT 74.635 -175.605 74.965 -175.275 ;
        RECT 74.635 -176.965 74.965 -176.635 ;
        RECT 74.635 -178.325 74.965 -177.995 ;
        RECT 74.635 -180.57 74.965 -179.44 ;
        RECT 74.64 -180.685 74.96 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 75.995 241.32 76.325 242.45 ;
        RECT 75.995 239.195 76.325 239.525 ;
        RECT 75.995 237.835 76.325 238.165 ;
        RECT 76 237.16 76.32 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 75.995 -95.365 76.325 -95.035 ;
        RECT 75.995 -96.725 76.325 -96.395 ;
        RECT 75.995 -98.085 76.325 -97.755 ;
        RECT 75.995 -99.445 76.325 -99.115 ;
        RECT 75.995 -100.805 76.325 -100.475 ;
        RECT 75.995 -102.165 76.325 -101.835 ;
        RECT 75.995 -103.525 76.325 -103.195 ;
        RECT 75.995 -104.885 76.325 -104.555 ;
        RECT 75.995 -106.245 76.325 -105.915 ;
        RECT 75.995 -107.605 76.325 -107.275 ;
        RECT 75.995 -108.965 76.325 -108.635 ;
        RECT 75.995 -110.325 76.325 -109.995 ;
        RECT 75.995 -111.685 76.325 -111.355 ;
        RECT 75.995 -113.045 76.325 -112.715 ;
        RECT 75.995 -114.405 76.325 -114.075 ;
        RECT 75.995 -115.765 76.325 -115.435 ;
        RECT 75.995 -117.125 76.325 -116.795 ;
        RECT 75.995 -118.485 76.325 -118.155 ;
        RECT 75.995 -119.845 76.325 -119.515 ;
        RECT 75.995 -121.205 76.325 -120.875 ;
        RECT 75.995 -122.565 76.325 -122.235 ;
        RECT 75.995 -123.925 76.325 -123.595 ;
        RECT 75.995 -125.285 76.325 -124.955 ;
        RECT 75.995 -126.645 76.325 -126.315 ;
        RECT 75.995 -128.005 76.325 -127.675 ;
        RECT 75.995 -129.365 76.325 -129.035 ;
        RECT 75.995 -130.725 76.325 -130.395 ;
        RECT 75.995 -132.085 76.325 -131.755 ;
        RECT 75.995 -133.445 76.325 -133.115 ;
        RECT 75.995 -134.805 76.325 -134.475 ;
        RECT 75.995 -136.165 76.325 -135.835 ;
        RECT 75.995 -137.525 76.325 -137.195 ;
        RECT 75.995 -138.885 76.325 -138.555 ;
        RECT 75.995 -140.245 76.325 -139.915 ;
        RECT 75.995 -141.605 76.325 -141.275 ;
        RECT 75.995 -142.965 76.325 -142.635 ;
        RECT 75.995 -144.325 76.325 -143.995 ;
        RECT 75.995 -145.685 76.325 -145.355 ;
        RECT 75.995 -147.045 76.325 -146.715 ;
        RECT 75.995 -148.405 76.325 -148.075 ;
        RECT 75.995 -149.765 76.325 -149.435 ;
        RECT 75.995 -151.125 76.325 -150.795 ;
        RECT 75.995 -152.485 76.325 -152.155 ;
        RECT 75.995 -153.845 76.325 -153.515 ;
        RECT 75.995 -155.205 76.325 -154.875 ;
        RECT 75.995 -156.565 76.325 -156.235 ;
        RECT 75.995 -157.925 76.325 -157.595 ;
        RECT 75.995 -159.285 76.325 -158.955 ;
        RECT 75.995 -160.645 76.325 -160.315 ;
        RECT 75.995 -162.005 76.325 -161.675 ;
        RECT 75.995 -163.365 76.325 -163.035 ;
        RECT 75.995 -164.725 76.325 -164.395 ;
        RECT 75.995 -166.085 76.325 -165.755 ;
        RECT 75.995 -167.445 76.325 -167.115 ;
        RECT 75.995 -168.805 76.325 -168.475 ;
        RECT 75.995 -170.165 76.325 -169.835 ;
        RECT 75.995 -171.525 76.325 -171.195 ;
        RECT 75.995 -172.885 76.325 -172.555 ;
        RECT 75.995 -174.245 76.325 -173.915 ;
        RECT 75.995 -175.605 76.325 -175.275 ;
        RECT 75.995 -176.965 76.325 -176.635 ;
        RECT 75.995 -178.325 76.325 -177.995 ;
        RECT 75.995 -180.57 76.325 -179.44 ;
        RECT 76 -180.685 76.32 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 76.51 -94.075 76.84 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 77.355 241.32 77.685 242.45 ;
        RECT 77.355 239.195 77.685 239.525 ;
        RECT 77.355 237.835 77.685 238.165 ;
        RECT 77.36 237.16 77.68 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 77.355 -1.525 77.685 -1.195 ;
        RECT 77.355 -2.885 77.685 -2.555 ;
        RECT 77.36 -3.56 77.68 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 78.715 241.32 79.045 242.45 ;
        RECT 78.715 239.195 79.045 239.525 ;
        RECT 78.715 237.835 79.045 238.165 ;
        RECT 78.72 237.16 79.04 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 78.715 -1.525 79.045 -1.195 ;
        RECT 78.715 -2.885 79.045 -2.555 ;
        RECT 78.72 -3.56 79.04 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 80.075 241.32 80.405 242.45 ;
        RECT 80.075 239.195 80.405 239.525 ;
        RECT 80.075 237.835 80.405 238.165 ;
        RECT 80.08 237.16 80.4 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 80.075 -1.525 80.405 -1.195 ;
        RECT 80.075 -2.885 80.405 -2.555 ;
        RECT 80.08 -3.56 80.4 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 80.075 -91.285 80.405 -90.955 ;
        RECT 80.075 -92.645 80.405 -92.315 ;
        RECT 80.075 -94.005 80.405 -93.675 ;
        RECT 80.075 -95.365 80.405 -95.035 ;
        RECT 80.075 -96.725 80.405 -96.395 ;
        RECT 80.075 -98.085 80.405 -97.755 ;
        RECT 80.075 -99.445 80.405 -99.115 ;
        RECT 80.075 -100.805 80.405 -100.475 ;
        RECT 80.075 -102.165 80.405 -101.835 ;
        RECT 80.075 -103.525 80.405 -103.195 ;
        RECT 80.075 -104.885 80.405 -104.555 ;
        RECT 80.075 -106.245 80.405 -105.915 ;
        RECT 80.075 -107.605 80.405 -107.275 ;
        RECT 80.075 -108.965 80.405 -108.635 ;
        RECT 80.075 -110.325 80.405 -109.995 ;
        RECT 80.075 -111.685 80.405 -111.355 ;
        RECT 80.075 -113.045 80.405 -112.715 ;
        RECT 80.075 -114.405 80.405 -114.075 ;
        RECT 80.075 -115.765 80.405 -115.435 ;
        RECT 80.075 -117.125 80.405 -116.795 ;
        RECT 80.075 -118.485 80.405 -118.155 ;
        RECT 80.075 -119.845 80.405 -119.515 ;
        RECT 80.075 -121.205 80.405 -120.875 ;
        RECT 80.075 -122.565 80.405 -122.235 ;
        RECT 80.075 -123.925 80.405 -123.595 ;
        RECT 80.075 -125.285 80.405 -124.955 ;
        RECT 80.075 -126.645 80.405 -126.315 ;
        RECT 80.075 -128.005 80.405 -127.675 ;
        RECT 80.075 -129.365 80.405 -129.035 ;
        RECT 80.075 -130.725 80.405 -130.395 ;
        RECT 80.075 -132.085 80.405 -131.755 ;
        RECT 80.075 -133.445 80.405 -133.115 ;
        RECT 80.075 -134.805 80.405 -134.475 ;
        RECT 80.075 -136.165 80.405 -135.835 ;
        RECT 80.075 -137.525 80.405 -137.195 ;
        RECT 80.075 -138.885 80.405 -138.555 ;
        RECT 80.075 -140.245 80.405 -139.915 ;
        RECT 80.075 -141.605 80.405 -141.275 ;
        RECT 80.075 -142.965 80.405 -142.635 ;
        RECT 80.075 -144.325 80.405 -143.995 ;
        RECT 80.075 -145.685 80.405 -145.355 ;
        RECT 80.075 -147.045 80.405 -146.715 ;
        RECT 80.075 -148.405 80.405 -148.075 ;
        RECT 80.075 -149.765 80.405 -149.435 ;
        RECT 80.075 -151.125 80.405 -150.795 ;
        RECT 80.075 -152.485 80.405 -152.155 ;
        RECT 80.075 -153.845 80.405 -153.515 ;
        RECT 80.075 -155.205 80.405 -154.875 ;
        RECT 80.075 -156.565 80.405 -156.235 ;
        RECT 80.075 -157.925 80.405 -157.595 ;
        RECT 80.075 -159.285 80.405 -158.955 ;
        RECT 80.075 -160.645 80.405 -160.315 ;
        RECT 80.075 -162.005 80.405 -161.675 ;
        RECT 80.075 -163.365 80.405 -163.035 ;
        RECT 80.075 -164.725 80.405 -164.395 ;
        RECT 80.075 -166.085 80.405 -165.755 ;
        RECT 80.075 -167.445 80.405 -167.115 ;
        RECT 80.075 -168.805 80.405 -168.475 ;
        RECT 80.075 -170.165 80.405 -169.835 ;
        RECT 80.075 -171.525 80.405 -171.195 ;
        RECT 80.075 -172.885 80.405 -172.555 ;
        RECT 80.075 -174.245 80.405 -173.915 ;
        RECT 80.075 -175.605 80.405 -175.275 ;
        RECT 80.075 -176.965 80.405 -176.635 ;
        RECT 80.075 -178.325 80.405 -177.995 ;
        RECT 80.075 -180.57 80.405 -179.44 ;
        RECT 80.08 -180.685 80.4 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 81.435 241.32 81.765 242.45 ;
        RECT 81.435 239.195 81.765 239.525 ;
        RECT 81.435 237.835 81.765 238.165 ;
        RECT 81.44 237.16 81.76 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 81.435 -95.365 81.765 -95.035 ;
        RECT 81.435 -96.725 81.765 -96.395 ;
        RECT 81.435 -98.085 81.765 -97.755 ;
        RECT 81.435 -99.445 81.765 -99.115 ;
        RECT 81.435 -100.805 81.765 -100.475 ;
        RECT 81.435 -102.165 81.765 -101.835 ;
        RECT 81.435 -103.525 81.765 -103.195 ;
        RECT 81.435 -104.885 81.765 -104.555 ;
        RECT 81.435 -106.245 81.765 -105.915 ;
        RECT 81.435 -107.605 81.765 -107.275 ;
        RECT 81.435 -108.965 81.765 -108.635 ;
        RECT 81.435 -110.325 81.765 -109.995 ;
        RECT 81.435 -111.685 81.765 -111.355 ;
        RECT 81.435 -113.045 81.765 -112.715 ;
        RECT 81.435 -114.405 81.765 -114.075 ;
        RECT 81.435 -115.765 81.765 -115.435 ;
        RECT 81.435 -117.125 81.765 -116.795 ;
        RECT 81.435 -118.485 81.765 -118.155 ;
        RECT 81.435 -119.845 81.765 -119.515 ;
        RECT 81.435 -121.205 81.765 -120.875 ;
        RECT 81.435 -122.565 81.765 -122.235 ;
        RECT 81.435 -123.925 81.765 -123.595 ;
        RECT 81.435 -125.285 81.765 -124.955 ;
        RECT 81.435 -126.645 81.765 -126.315 ;
        RECT 81.435 -128.005 81.765 -127.675 ;
        RECT 81.435 -129.365 81.765 -129.035 ;
        RECT 81.435 -130.725 81.765 -130.395 ;
        RECT 81.435 -132.085 81.765 -131.755 ;
        RECT 81.435 -133.445 81.765 -133.115 ;
        RECT 81.435 -134.805 81.765 -134.475 ;
        RECT 81.435 -136.165 81.765 -135.835 ;
        RECT 81.435 -137.525 81.765 -137.195 ;
        RECT 81.435 -138.885 81.765 -138.555 ;
        RECT 81.435 -140.245 81.765 -139.915 ;
        RECT 81.435 -141.605 81.765 -141.275 ;
        RECT 81.435 -142.965 81.765 -142.635 ;
        RECT 81.435 -144.325 81.765 -143.995 ;
        RECT 81.435 -145.685 81.765 -145.355 ;
        RECT 81.435 -147.045 81.765 -146.715 ;
        RECT 81.435 -148.405 81.765 -148.075 ;
        RECT 81.435 -149.765 81.765 -149.435 ;
        RECT 81.435 -151.125 81.765 -150.795 ;
        RECT 81.435 -152.485 81.765 -152.155 ;
        RECT 81.435 -153.845 81.765 -153.515 ;
        RECT 81.435 -155.205 81.765 -154.875 ;
        RECT 81.435 -156.565 81.765 -156.235 ;
        RECT 81.435 -157.925 81.765 -157.595 ;
        RECT 81.435 -159.285 81.765 -158.955 ;
        RECT 81.435 -160.645 81.765 -160.315 ;
        RECT 81.435 -162.005 81.765 -161.675 ;
        RECT 81.435 -163.365 81.765 -163.035 ;
        RECT 81.435 -164.725 81.765 -164.395 ;
        RECT 81.435 -166.085 81.765 -165.755 ;
        RECT 81.435 -167.445 81.765 -167.115 ;
        RECT 81.435 -168.805 81.765 -168.475 ;
        RECT 81.435 -170.165 81.765 -169.835 ;
        RECT 81.435 -171.525 81.765 -171.195 ;
        RECT 81.435 -172.885 81.765 -172.555 ;
        RECT 81.435 -174.245 81.765 -173.915 ;
        RECT 81.435 -175.605 81.765 -175.275 ;
        RECT 81.435 -176.965 81.765 -176.635 ;
        RECT 81.435 -178.325 81.765 -177.995 ;
        RECT 81.435 -180.57 81.765 -179.44 ;
        RECT 81.44 -180.685 81.76 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 82.61 -94.075 82.94 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 82.795 241.32 83.125 242.45 ;
        RECT 82.795 239.195 83.125 239.525 ;
        RECT 82.795 237.835 83.125 238.165 ;
        RECT 82.8 237.16 83.12 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 84.155 241.32 84.485 242.45 ;
        RECT 84.155 239.195 84.485 239.525 ;
        RECT 84.155 237.835 84.485 238.165 ;
        RECT 84.16 237.16 84.48 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 84.155 -1.525 84.485 -1.195 ;
        RECT 84.155 -2.885 84.485 -2.555 ;
        RECT 84.16 -3.56 84.48 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 84.155 -91.285 84.485 -90.955 ;
        RECT 84.155 -92.645 84.485 -92.315 ;
        RECT 84.155 -94.005 84.485 -93.675 ;
        RECT 84.155 -95.365 84.485 -95.035 ;
        RECT 84.155 -96.725 84.485 -96.395 ;
        RECT 84.155 -98.085 84.485 -97.755 ;
        RECT 84.155 -99.445 84.485 -99.115 ;
        RECT 84.155 -100.805 84.485 -100.475 ;
        RECT 84.155 -102.165 84.485 -101.835 ;
        RECT 84.155 -103.525 84.485 -103.195 ;
        RECT 84.155 -104.885 84.485 -104.555 ;
        RECT 84.155 -106.245 84.485 -105.915 ;
        RECT 84.155 -107.605 84.485 -107.275 ;
        RECT 84.155 -108.965 84.485 -108.635 ;
        RECT 84.155 -110.325 84.485 -109.995 ;
        RECT 84.155 -111.685 84.485 -111.355 ;
        RECT 84.155 -113.045 84.485 -112.715 ;
        RECT 84.155 -114.405 84.485 -114.075 ;
        RECT 84.155 -115.765 84.485 -115.435 ;
        RECT 84.155 -117.125 84.485 -116.795 ;
        RECT 84.155 -118.485 84.485 -118.155 ;
        RECT 84.155 -119.845 84.485 -119.515 ;
        RECT 84.155 -121.205 84.485 -120.875 ;
        RECT 84.155 -122.565 84.485 -122.235 ;
        RECT 84.155 -123.925 84.485 -123.595 ;
        RECT 84.155 -125.285 84.485 -124.955 ;
        RECT 84.155 -126.645 84.485 -126.315 ;
        RECT 84.155 -128.005 84.485 -127.675 ;
        RECT 84.155 -129.365 84.485 -129.035 ;
        RECT 84.155 -130.725 84.485 -130.395 ;
        RECT 84.155 -132.085 84.485 -131.755 ;
        RECT 84.155 -133.445 84.485 -133.115 ;
        RECT 84.155 -134.805 84.485 -134.475 ;
        RECT 84.155 -136.165 84.485 -135.835 ;
        RECT 84.155 -137.525 84.485 -137.195 ;
        RECT 84.155 -138.885 84.485 -138.555 ;
        RECT 84.155 -140.245 84.485 -139.915 ;
        RECT 84.155 -141.605 84.485 -141.275 ;
        RECT 84.155 -142.965 84.485 -142.635 ;
        RECT 84.155 -144.325 84.485 -143.995 ;
        RECT 84.155 -145.685 84.485 -145.355 ;
        RECT 84.155 -147.045 84.485 -146.715 ;
        RECT 84.155 -148.405 84.485 -148.075 ;
        RECT 84.155 -149.765 84.485 -149.435 ;
        RECT 84.155 -151.125 84.485 -150.795 ;
        RECT 84.155 -152.485 84.485 -152.155 ;
        RECT 84.155 -153.845 84.485 -153.515 ;
        RECT 84.155 -155.205 84.485 -154.875 ;
        RECT 84.155 -156.565 84.485 -156.235 ;
        RECT 84.155 -157.925 84.485 -157.595 ;
        RECT 84.155 -159.285 84.485 -158.955 ;
        RECT 84.155 -160.645 84.485 -160.315 ;
        RECT 84.155 -162.005 84.485 -161.675 ;
        RECT 84.155 -163.365 84.485 -163.035 ;
        RECT 84.155 -164.725 84.485 -164.395 ;
        RECT 84.155 -166.085 84.485 -165.755 ;
        RECT 84.155 -167.445 84.485 -167.115 ;
        RECT 84.155 -168.805 84.485 -168.475 ;
        RECT 84.155 -170.165 84.485 -169.835 ;
        RECT 84.155 -171.525 84.485 -171.195 ;
        RECT 84.155 -172.885 84.485 -172.555 ;
        RECT 84.155 -174.245 84.485 -173.915 ;
        RECT 84.155 -175.605 84.485 -175.275 ;
        RECT 84.155 -176.965 84.485 -176.635 ;
        RECT 84.155 -178.325 84.485 -177.995 ;
        RECT 84.155 -180.57 84.485 -179.44 ;
        RECT 84.16 -180.685 84.48 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 85.515 241.32 85.845 242.45 ;
        RECT 85.515 239.195 85.845 239.525 ;
        RECT 85.515 237.835 85.845 238.165 ;
        RECT 85.52 237.16 85.84 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 85.515 -1.525 85.845 -1.195 ;
        RECT 85.515 -2.885 85.845 -2.555 ;
        RECT 85.52 -3.56 85.84 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 86.875 241.32 87.205 242.45 ;
        RECT 86.875 239.195 87.205 239.525 ;
        RECT 86.875 237.835 87.205 238.165 ;
        RECT 86.88 237.16 87.2 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 86.875 -1.525 87.205 -1.195 ;
        RECT 86.875 -2.885 87.205 -2.555 ;
        RECT 86.88 -3.56 87.2 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 86.875 -91.285 87.205 -90.955 ;
        RECT 86.875 -92.645 87.205 -92.315 ;
        RECT 86.875 -94.005 87.205 -93.675 ;
        RECT 86.875 -95.365 87.205 -95.035 ;
        RECT 86.875 -96.725 87.205 -96.395 ;
        RECT 86.875 -98.085 87.205 -97.755 ;
        RECT 86.875 -99.445 87.205 -99.115 ;
        RECT 86.875 -100.805 87.205 -100.475 ;
        RECT 86.875 -102.165 87.205 -101.835 ;
        RECT 86.875 -103.525 87.205 -103.195 ;
        RECT 86.875 -104.885 87.205 -104.555 ;
        RECT 86.875 -106.245 87.205 -105.915 ;
        RECT 86.875 -107.605 87.205 -107.275 ;
        RECT 86.875 -108.965 87.205 -108.635 ;
        RECT 86.875 -110.325 87.205 -109.995 ;
        RECT 86.875 -111.685 87.205 -111.355 ;
        RECT 86.875 -113.045 87.205 -112.715 ;
        RECT 86.875 -114.405 87.205 -114.075 ;
        RECT 86.875 -115.765 87.205 -115.435 ;
        RECT 86.875 -117.125 87.205 -116.795 ;
        RECT 86.875 -118.485 87.205 -118.155 ;
        RECT 86.875 -119.845 87.205 -119.515 ;
        RECT 86.875 -121.205 87.205 -120.875 ;
        RECT 86.875 -122.565 87.205 -122.235 ;
        RECT 86.875 -123.925 87.205 -123.595 ;
        RECT 86.875 -125.285 87.205 -124.955 ;
        RECT 86.875 -126.645 87.205 -126.315 ;
        RECT 86.875 -128.005 87.205 -127.675 ;
        RECT 86.875 -129.365 87.205 -129.035 ;
        RECT 86.875 -130.725 87.205 -130.395 ;
        RECT 86.875 -132.085 87.205 -131.755 ;
        RECT 86.875 -133.445 87.205 -133.115 ;
        RECT 86.875 -134.805 87.205 -134.475 ;
        RECT 86.875 -136.165 87.205 -135.835 ;
        RECT 86.875 -137.525 87.205 -137.195 ;
        RECT 86.875 -138.885 87.205 -138.555 ;
        RECT 86.875 -140.245 87.205 -139.915 ;
        RECT 86.875 -141.605 87.205 -141.275 ;
        RECT 86.875 -142.965 87.205 -142.635 ;
        RECT 86.875 -144.325 87.205 -143.995 ;
        RECT 86.875 -145.685 87.205 -145.355 ;
        RECT 86.875 -147.045 87.205 -146.715 ;
        RECT 86.875 -148.405 87.205 -148.075 ;
        RECT 86.875 -149.765 87.205 -149.435 ;
        RECT 86.875 -151.125 87.205 -150.795 ;
        RECT 86.875 -152.485 87.205 -152.155 ;
        RECT 86.875 -153.845 87.205 -153.515 ;
        RECT 86.875 -155.205 87.205 -154.875 ;
        RECT 86.875 -156.565 87.205 -156.235 ;
        RECT 86.875 -157.925 87.205 -157.595 ;
        RECT 86.875 -159.285 87.205 -158.955 ;
        RECT 86.875 -160.645 87.205 -160.315 ;
        RECT 86.875 -162.005 87.205 -161.675 ;
        RECT 86.875 -163.365 87.205 -163.035 ;
        RECT 86.875 -164.725 87.205 -164.395 ;
        RECT 86.875 -166.085 87.205 -165.755 ;
        RECT 86.875 -167.445 87.205 -167.115 ;
        RECT 86.875 -168.805 87.205 -168.475 ;
        RECT 86.875 -170.165 87.205 -169.835 ;
        RECT 86.875 -171.525 87.205 -171.195 ;
        RECT 86.875 -172.885 87.205 -172.555 ;
        RECT 86.875 -174.245 87.205 -173.915 ;
        RECT 86.875 -175.605 87.205 -175.275 ;
        RECT 86.875 -176.965 87.205 -176.635 ;
        RECT 86.875 -178.325 87.205 -177.995 ;
        RECT 86.875 -180.57 87.205 -179.44 ;
        RECT 86.88 -180.685 87.2 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 88.235 241.32 88.565 242.45 ;
        RECT 88.235 239.195 88.565 239.525 ;
        RECT 88.235 237.835 88.565 238.165 ;
        RECT 88.24 237.16 88.56 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 88.235 -95.365 88.565 -95.035 ;
        RECT 88.235 -96.725 88.565 -96.395 ;
        RECT 88.235 -98.085 88.565 -97.755 ;
        RECT 88.235 -99.445 88.565 -99.115 ;
        RECT 88.235 -100.805 88.565 -100.475 ;
        RECT 88.235 -102.165 88.565 -101.835 ;
        RECT 88.235 -103.525 88.565 -103.195 ;
        RECT 88.235 -104.885 88.565 -104.555 ;
        RECT 88.235 -106.245 88.565 -105.915 ;
        RECT 88.235 -107.605 88.565 -107.275 ;
        RECT 88.235 -108.965 88.565 -108.635 ;
        RECT 88.235 -110.325 88.565 -109.995 ;
        RECT 88.235 -111.685 88.565 -111.355 ;
        RECT 88.235 -113.045 88.565 -112.715 ;
        RECT 88.235 -114.405 88.565 -114.075 ;
        RECT 88.235 -115.765 88.565 -115.435 ;
        RECT 88.235 -117.125 88.565 -116.795 ;
        RECT 88.235 -118.485 88.565 -118.155 ;
        RECT 88.235 -119.845 88.565 -119.515 ;
        RECT 88.235 -121.205 88.565 -120.875 ;
        RECT 88.235 -122.565 88.565 -122.235 ;
        RECT 88.235 -123.925 88.565 -123.595 ;
        RECT 88.235 -125.285 88.565 -124.955 ;
        RECT 88.235 -126.645 88.565 -126.315 ;
        RECT 88.235 -128.005 88.565 -127.675 ;
        RECT 88.235 -129.365 88.565 -129.035 ;
        RECT 88.235 -130.725 88.565 -130.395 ;
        RECT 88.235 -132.085 88.565 -131.755 ;
        RECT 88.235 -133.445 88.565 -133.115 ;
        RECT 88.235 -134.805 88.565 -134.475 ;
        RECT 88.235 -136.165 88.565 -135.835 ;
        RECT 88.235 -137.525 88.565 -137.195 ;
        RECT 88.235 -138.885 88.565 -138.555 ;
        RECT 88.235 -140.245 88.565 -139.915 ;
        RECT 88.235 -141.605 88.565 -141.275 ;
        RECT 88.235 -142.965 88.565 -142.635 ;
        RECT 88.235 -144.325 88.565 -143.995 ;
        RECT 88.235 -145.685 88.565 -145.355 ;
        RECT 88.235 -147.045 88.565 -146.715 ;
        RECT 88.235 -148.405 88.565 -148.075 ;
        RECT 88.235 -149.765 88.565 -149.435 ;
        RECT 88.235 -151.125 88.565 -150.795 ;
        RECT 88.235 -152.485 88.565 -152.155 ;
        RECT 88.235 -153.845 88.565 -153.515 ;
        RECT 88.235 -155.205 88.565 -154.875 ;
        RECT 88.235 -156.565 88.565 -156.235 ;
        RECT 88.235 -157.925 88.565 -157.595 ;
        RECT 88.235 -159.285 88.565 -158.955 ;
        RECT 88.235 -160.645 88.565 -160.315 ;
        RECT 88.235 -162.005 88.565 -161.675 ;
        RECT 88.235 -163.365 88.565 -163.035 ;
        RECT 88.235 -164.725 88.565 -164.395 ;
        RECT 88.235 -166.085 88.565 -165.755 ;
        RECT 88.235 -167.445 88.565 -167.115 ;
        RECT 88.235 -168.805 88.565 -168.475 ;
        RECT 88.235 -170.165 88.565 -169.835 ;
        RECT 88.235 -171.525 88.565 -171.195 ;
        RECT 88.235 -172.885 88.565 -172.555 ;
        RECT 88.235 -174.245 88.565 -173.915 ;
        RECT 88.235 -175.605 88.565 -175.275 ;
        RECT 88.235 -176.965 88.565 -176.635 ;
        RECT 88.235 -178.325 88.565 -177.995 ;
        RECT 88.235 -180.57 88.565 -179.44 ;
        RECT 88.24 -180.685 88.56 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 88.71 -94.075 89.04 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 89.595 241.32 89.925 242.45 ;
        RECT 89.595 239.195 89.925 239.525 ;
        RECT 89.595 237.835 89.925 238.165 ;
        RECT 89.6 237.16 89.92 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 89.595 -1.525 89.925 -1.195 ;
        RECT 89.595 -2.885 89.925 -2.555 ;
        RECT 89.6 -3.56 89.92 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 90.955 241.32 91.285 242.45 ;
        RECT 90.955 239.195 91.285 239.525 ;
        RECT 90.955 237.835 91.285 238.165 ;
        RECT 90.96 237.16 91.28 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 90.955 -1.525 91.285 -1.195 ;
        RECT 90.955 -2.885 91.285 -2.555 ;
        RECT 90.96 -3.56 91.28 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 92.315 241.32 92.645 242.45 ;
        RECT 92.315 239.195 92.645 239.525 ;
        RECT 92.315 237.835 92.645 238.165 ;
        RECT 92.32 237.16 92.64 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 92.315 -1.525 92.645 -1.195 ;
        RECT 92.315 -2.885 92.645 -2.555 ;
        RECT 92.32 -3.56 92.64 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 92.315 -91.285 92.645 -90.955 ;
        RECT 92.315 -92.645 92.645 -92.315 ;
        RECT 92.315 -94.005 92.645 -93.675 ;
        RECT 92.315 -95.365 92.645 -95.035 ;
        RECT 92.315 -96.725 92.645 -96.395 ;
        RECT 92.315 -98.085 92.645 -97.755 ;
        RECT 92.315 -99.445 92.645 -99.115 ;
        RECT 92.315 -100.805 92.645 -100.475 ;
        RECT 92.315 -102.165 92.645 -101.835 ;
        RECT 92.315 -103.525 92.645 -103.195 ;
        RECT 92.315 -104.885 92.645 -104.555 ;
        RECT 92.315 -106.245 92.645 -105.915 ;
        RECT 92.315 -107.605 92.645 -107.275 ;
        RECT 92.315 -108.965 92.645 -108.635 ;
        RECT 92.315 -110.325 92.645 -109.995 ;
        RECT 92.315 -111.685 92.645 -111.355 ;
        RECT 92.315 -113.045 92.645 -112.715 ;
        RECT 92.315 -114.405 92.645 -114.075 ;
        RECT 92.315 -115.765 92.645 -115.435 ;
        RECT 92.315 -117.125 92.645 -116.795 ;
        RECT 92.315 -118.485 92.645 -118.155 ;
        RECT 92.315 -119.845 92.645 -119.515 ;
        RECT 92.315 -121.205 92.645 -120.875 ;
        RECT 92.315 -122.565 92.645 -122.235 ;
        RECT 92.315 -123.925 92.645 -123.595 ;
        RECT 92.315 -125.285 92.645 -124.955 ;
        RECT 92.315 -126.645 92.645 -126.315 ;
        RECT 92.315 -128.005 92.645 -127.675 ;
        RECT 92.315 -129.365 92.645 -129.035 ;
        RECT 92.315 -130.725 92.645 -130.395 ;
        RECT 92.315 -132.085 92.645 -131.755 ;
        RECT 92.315 -133.445 92.645 -133.115 ;
        RECT 92.315 -134.805 92.645 -134.475 ;
        RECT 92.315 -136.165 92.645 -135.835 ;
        RECT 92.315 -137.525 92.645 -137.195 ;
        RECT 92.315 -138.885 92.645 -138.555 ;
        RECT 92.315 -140.245 92.645 -139.915 ;
        RECT 92.315 -141.605 92.645 -141.275 ;
        RECT 92.315 -142.965 92.645 -142.635 ;
        RECT 92.315 -144.325 92.645 -143.995 ;
        RECT 92.315 -145.685 92.645 -145.355 ;
        RECT 92.315 -147.045 92.645 -146.715 ;
        RECT 92.315 -148.405 92.645 -148.075 ;
        RECT 92.315 -149.765 92.645 -149.435 ;
        RECT 92.315 -151.125 92.645 -150.795 ;
        RECT 92.315 -152.485 92.645 -152.155 ;
        RECT 92.315 -153.845 92.645 -153.515 ;
        RECT 92.315 -155.205 92.645 -154.875 ;
        RECT 92.315 -156.565 92.645 -156.235 ;
        RECT 92.315 -157.925 92.645 -157.595 ;
        RECT 92.315 -159.285 92.645 -158.955 ;
        RECT 92.315 -160.645 92.645 -160.315 ;
        RECT 92.315 -162.005 92.645 -161.675 ;
        RECT 92.315 -163.365 92.645 -163.035 ;
        RECT 92.315 -164.725 92.645 -164.395 ;
        RECT 92.315 -166.085 92.645 -165.755 ;
        RECT 92.315 -167.445 92.645 -167.115 ;
        RECT 92.315 -168.805 92.645 -168.475 ;
        RECT 92.315 -170.165 92.645 -169.835 ;
        RECT 92.315 -171.525 92.645 -171.195 ;
        RECT 92.315 -172.885 92.645 -172.555 ;
        RECT 92.315 -174.245 92.645 -173.915 ;
        RECT 92.315 -175.605 92.645 -175.275 ;
        RECT 92.315 -176.965 92.645 -176.635 ;
        RECT 92.315 -178.325 92.645 -177.995 ;
        RECT 92.315 -180.57 92.645 -179.44 ;
        RECT 92.32 -180.685 92.64 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 93.675 241.32 94.005 242.45 ;
        RECT 93.675 239.195 94.005 239.525 ;
        RECT 93.675 237.835 94.005 238.165 ;
        RECT 93.68 237.16 94 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 93.675 -95.365 94.005 -95.035 ;
        RECT 93.675 -96.725 94.005 -96.395 ;
        RECT 93.675 -98.085 94.005 -97.755 ;
        RECT 93.675 -99.445 94.005 -99.115 ;
        RECT 93.675 -100.805 94.005 -100.475 ;
        RECT 93.675 -102.165 94.005 -101.835 ;
        RECT 93.675 -103.525 94.005 -103.195 ;
        RECT 93.675 -104.885 94.005 -104.555 ;
        RECT 93.675 -106.245 94.005 -105.915 ;
        RECT 93.675 -107.605 94.005 -107.275 ;
        RECT 93.675 -108.965 94.005 -108.635 ;
        RECT 93.675 -110.325 94.005 -109.995 ;
        RECT 93.675 -111.685 94.005 -111.355 ;
        RECT 93.675 -113.045 94.005 -112.715 ;
        RECT 93.675 -114.405 94.005 -114.075 ;
        RECT 93.675 -115.765 94.005 -115.435 ;
        RECT 93.675 -117.125 94.005 -116.795 ;
        RECT 93.675 -118.485 94.005 -118.155 ;
        RECT 93.675 -119.845 94.005 -119.515 ;
        RECT 93.675 -121.205 94.005 -120.875 ;
        RECT 93.675 -122.565 94.005 -122.235 ;
        RECT 93.675 -123.925 94.005 -123.595 ;
        RECT 93.675 -125.285 94.005 -124.955 ;
        RECT 93.675 -126.645 94.005 -126.315 ;
        RECT 93.675 -128.005 94.005 -127.675 ;
        RECT 93.675 -129.365 94.005 -129.035 ;
        RECT 93.675 -130.725 94.005 -130.395 ;
        RECT 93.675 -132.085 94.005 -131.755 ;
        RECT 93.675 -133.445 94.005 -133.115 ;
        RECT 93.675 -134.805 94.005 -134.475 ;
        RECT 93.675 -136.165 94.005 -135.835 ;
        RECT 93.675 -137.525 94.005 -137.195 ;
        RECT 93.675 -138.885 94.005 -138.555 ;
        RECT 93.675 -140.245 94.005 -139.915 ;
        RECT 93.675 -141.605 94.005 -141.275 ;
        RECT 93.675 -142.965 94.005 -142.635 ;
        RECT 93.675 -144.325 94.005 -143.995 ;
        RECT 93.675 -145.685 94.005 -145.355 ;
        RECT 93.675 -147.045 94.005 -146.715 ;
        RECT 93.675 -148.405 94.005 -148.075 ;
        RECT 93.675 -149.765 94.005 -149.435 ;
        RECT 93.675 -151.125 94.005 -150.795 ;
        RECT 93.675 -152.485 94.005 -152.155 ;
        RECT 93.675 -153.845 94.005 -153.515 ;
        RECT 93.675 -155.205 94.005 -154.875 ;
        RECT 93.675 -156.565 94.005 -156.235 ;
        RECT 93.675 -157.925 94.005 -157.595 ;
        RECT 93.675 -159.285 94.005 -158.955 ;
        RECT 93.675 -160.645 94.005 -160.315 ;
        RECT 93.675 -162.005 94.005 -161.675 ;
        RECT 93.675 -163.365 94.005 -163.035 ;
        RECT 93.675 -164.725 94.005 -164.395 ;
        RECT 93.675 -166.085 94.005 -165.755 ;
        RECT 93.675 -167.445 94.005 -167.115 ;
        RECT 93.675 -168.805 94.005 -168.475 ;
        RECT 93.675 -170.165 94.005 -169.835 ;
        RECT 93.675 -171.525 94.005 -171.195 ;
        RECT 93.675 -172.885 94.005 -172.555 ;
        RECT 93.675 -174.245 94.005 -173.915 ;
        RECT 93.675 -175.605 94.005 -175.275 ;
        RECT 93.675 -176.965 94.005 -176.635 ;
        RECT 93.675 -178.325 94.005 -177.995 ;
        RECT 93.675 -180.57 94.005 -179.44 ;
        RECT 93.68 -180.685 94 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 94.81 -94.075 95.14 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 95.035 241.32 95.365 242.45 ;
        RECT 95.035 239.195 95.365 239.525 ;
        RECT 95.035 237.835 95.365 238.165 ;
        RECT 95.04 237.16 95.36 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 96.395 241.32 96.725 242.45 ;
        RECT 96.395 239.195 96.725 239.525 ;
        RECT 96.395 237.835 96.725 238.165 ;
        RECT 96.4 237.16 96.72 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 96.395 -1.525 96.725 -1.195 ;
        RECT 96.395 -2.885 96.725 -2.555 ;
        RECT 96.4 -3.56 96.72 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 96.395 -91.285 96.725 -90.955 ;
        RECT 96.395 -92.645 96.725 -92.315 ;
        RECT 96.395 -94.005 96.725 -93.675 ;
        RECT 96.395 -95.365 96.725 -95.035 ;
        RECT 96.395 -96.725 96.725 -96.395 ;
        RECT 96.395 -98.085 96.725 -97.755 ;
        RECT 96.395 -99.445 96.725 -99.115 ;
        RECT 96.395 -100.805 96.725 -100.475 ;
        RECT 96.395 -102.165 96.725 -101.835 ;
        RECT 96.395 -103.525 96.725 -103.195 ;
        RECT 96.395 -104.885 96.725 -104.555 ;
        RECT 96.395 -106.245 96.725 -105.915 ;
        RECT 96.395 -107.605 96.725 -107.275 ;
        RECT 96.395 -108.965 96.725 -108.635 ;
        RECT 96.395 -110.325 96.725 -109.995 ;
        RECT 96.395 -111.685 96.725 -111.355 ;
        RECT 96.395 -113.045 96.725 -112.715 ;
        RECT 96.395 -114.405 96.725 -114.075 ;
        RECT 96.395 -115.765 96.725 -115.435 ;
        RECT 96.395 -117.125 96.725 -116.795 ;
        RECT 96.395 -118.485 96.725 -118.155 ;
        RECT 96.395 -119.845 96.725 -119.515 ;
        RECT 96.395 -121.205 96.725 -120.875 ;
        RECT 96.395 -122.565 96.725 -122.235 ;
        RECT 96.395 -123.925 96.725 -123.595 ;
        RECT 96.395 -125.285 96.725 -124.955 ;
        RECT 96.395 -126.645 96.725 -126.315 ;
        RECT 96.395 -128.005 96.725 -127.675 ;
        RECT 96.395 -129.365 96.725 -129.035 ;
        RECT 96.395 -130.725 96.725 -130.395 ;
        RECT 96.395 -132.085 96.725 -131.755 ;
        RECT 96.395 -133.445 96.725 -133.115 ;
        RECT 96.395 -134.805 96.725 -134.475 ;
        RECT 96.395 -136.165 96.725 -135.835 ;
        RECT 96.395 -137.525 96.725 -137.195 ;
        RECT 96.395 -138.885 96.725 -138.555 ;
        RECT 96.395 -140.245 96.725 -139.915 ;
        RECT 96.395 -141.605 96.725 -141.275 ;
        RECT 96.395 -142.965 96.725 -142.635 ;
        RECT 96.395 -144.325 96.725 -143.995 ;
        RECT 96.395 -145.685 96.725 -145.355 ;
        RECT 96.395 -147.045 96.725 -146.715 ;
        RECT 96.395 -148.405 96.725 -148.075 ;
        RECT 96.395 -149.765 96.725 -149.435 ;
        RECT 96.395 -151.125 96.725 -150.795 ;
        RECT 96.395 -152.485 96.725 -152.155 ;
        RECT 96.395 -153.845 96.725 -153.515 ;
        RECT 96.395 -155.205 96.725 -154.875 ;
        RECT 96.395 -156.565 96.725 -156.235 ;
        RECT 96.395 -157.925 96.725 -157.595 ;
        RECT 96.395 -159.285 96.725 -158.955 ;
        RECT 96.395 -160.645 96.725 -160.315 ;
        RECT 96.395 -162.005 96.725 -161.675 ;
        RECT 96.395 -163.365 96.725 -163.035 ;
        RECT 96.395 -164.725 96.725 -164.395 ;
        RECT 96.395 -166.085 96.725 -165.755 ;
        RECT 96.395 -167.445 96.725 -167.115 ;
        RECT 96.395 -168.805 96.725 -168.475 ;
        RECT 96.395 -170.165 96.725 -169.835 ;
        RECT 96.395 -171.525 96.725 -171.195 ;
        RECT 96.395 -172.885 96.725 -172.555 ;
        RECT 96.395 -174.245 96.725 -173.915 ;
        RECT 96.395 -175.605 96.725 -175.275 ;
        RECT 96.395 -176.965 96.725 -176.635 ;
        RECT 96.395 -178.325 96.725 -177.995 ;
        RECT 96.395 -180.57 96.725 -179.44 ;
        RECT 96.4 -180.685 96.72 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 97.755 241.32 98.085 242.45 ;
        RECT 97.755 239.195 98.085 239.525 ;
        RECT 97.755 237.835 98.085 238.165 ;
        RECT 97.76 237.16 98.08 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 97.755 -1.525 98.085 -1.195 ;
        RECT 97.755 -2.885 98.085 -2.555 ;
        RECT 97.76 -3.56 98.08 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 99.115 241.32 99.445 242.45 ;
        RECT 99.115 239.195 99.445 239.525 ;
        RECT 99.115 237.835 99.445 238.165 ;
        RECT 99.12 237.16 99.44 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 99.115 -1.525 99.445 -1.195 ;
        RECT 99.115 -2.885 99.445 -2.555 ;
        RECT 99.12 -3.56 99.44 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 99.115 -123.925 99.445 -123.595 ;
        RECT 99.115 -125.285 99.445 -124.955 ;
        RECT 99.115 -126.645 99.445 -126.315 ;
        RECT 99.115 -128.005 99.445 -127.675 ;
        RECT 99.115 -129.365 99.445 -129.035 ;
        RECT 99.115 -130.725 99.445 -130.395 ;
        RECT 99.115 -132.085 99.445 -131.755 ;
        RECT 99.115 -133.445 99.445 -133.115 ;
        RECT 99.115 -134.805 99.445 -134.475 ;
        RECT 99.115 -136.165 99.445 -135.835 ;
        RECT 99.115 -137.525 99.445 -137.195 ;
        RECT 99.115 -138.885 99.445 -138.555 ;
        RECT 99.115 -140.245 99.445 -139.915 ;
        RECT 99.115 -141.605 99.445 -141.275 ;
        RECT 99.115 -142.965 99.445 -142.635 ;
        RECT 99.115 -144.325 99.445 -143.995 ;
        RECT 99.115 -145.685 99.445 -145.355 ;
        RECT 99.115 -147.045 99.445 -146.715 ;
        RECT 99.115 -148.405 99.445 -148.075 ;
        RECT 99.115 -149.765 99.445 -149.435 ;
        RECT 99.115 -151.125 99.445 -150.795 ;
        RECT 99.115 -152.485 99.445 -152.155 ;
        RECT 99.115 -153.845 99.445 -153.515 ;
        RECT 99.115 -155.205 99.445 -154.875 ;
        RECT 99.115 -156.565 99.445 -156.235 ;
        RECT 99.115 -157.925 99.445 -157.595 ;
        RECT 99.115 -159.285 99.445 -158.955 ;
        RECT 99.115 -160.645 99.445 -160.315 ;
        RECT 99.115 -162.005 99.445 -161.675 ;
        RECT 99.115 -163.365 99.445 -163.035 ;
        RECT 99.115 -164.725 99.445 -164.395 ;
        RECT 99.115 -166.085 99.445 -165.755 ;
        RECT 99.115 -167.445 99.445 -167.115 ;
        RECT 99.115 -168.805 99.445 -168.475 ;
        RECT 99.115 -170.165 99.445 -169.835 ;
        RECT 99.115 -171.525 99.445 -171.195 ;
        RECT 99.115 -172.885 99.445 -172.555 ;
        RECT 99.115 -174.245 99.445 -173.915 ;
        RECT 99.115 -175.605 99.445 -175.275 ;
        RECT 99.115 -176.965 99.445 -176.635 ;
        RECT 99.115 -178.325 99.445 -177.995 ;
        RECT 99.115 -180.57 99.445 -179.44 ;
        RECT 99.12 -180.685 99.44 -90.955 ;
        RECT 99.115 -91.285 99.445 -90.955 ;
        RECT 99.115 -92.645 99.445 -92.315 ;
        RECT 99.115 -94.005 99.445 -93.675 ;
        RECT 99.115 -95.365 99.445 -95.035 ;
        RECT 99.115 -96.725 99.445 -96.395 ;
        RECT 99.115 -98.085 99.445 -97.755 ;
        RECT 99.115 -99.445 99.445 -99.115 ;
        RECT 99.115 -100.805 99.445 -100.475 ;
        RECT 99.115 -102.165 99.445 -101.835 ;
        RECT 99.115 -103.525 99.445 -103.195 ;
        RECT 99.115 -104.885 99.445 -104.555 ;
        RECT 99.115 -106.245 99.445 -105.915 ;
        RECT 99.115 -107.605 99.445 -107.275 ;
        RECT 99.115 -108.965 99.445 -108.635 ;
        RECT 99.115 -110.325 99.445 -109.995 ;
        RECT 99.115 -111.685 99.445 -111.355 ;
        RECT 99.115 -113.045 99.445 -112.715 ;
        RECT 99.115 -114.405 99.445 -114.075 ;
        RECT 99.115 -115.765 99.445 -115.435 ;
        RECT 99.115 -117.125 99.445 -116.795 ;
        RECT 99.115 -118.485 99.445 -118.155 ;
        RECT 99.115 -119.845 99.445 -119.515 ;
        RECT 99.115 -121.205 99.445 -120.875 ;
        RECT 99.115 -122.565 99.445 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT 32.475 241.32 32.805 242.45 ;
        RECT 32.475 239.195 32.805 239.525 ;
        RECT 32.475 237.835 32.805 238.165 ;
        RECT 32.48 237.16 32.8 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 32.475 -1.525 32.805 -1.195 ;
        RECT 32.475 -2.885 32.805 -2.555 ;
        RECT 32.48 -3.56 32.8 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 32.475 -91.285 32.805 -90.955 ;
        RECT 32.475 -92.645 32.805 -92.315 ;
        RECT 32.475 -94.005 32.805 -93.675 ;
        RECT 32.475 -95.365 32.805 -95.035 ;
        RECT 32.475 -96.725 32.805 -96.395 ;
        RECT 32.475 -98.085 32.805 -97.755 ;
        RECT 32.475 -99.445 32.805 -99.115 ;
        RECT 32.475 -100.805 32.805 -100.475 ;
        RECT 32.475 -102.165 32.805 -101.835 ;
        RECT 32.475 -103.525 32.805 -103.195 ;
        RECT 32.475 -104.885 32.805 -104.555 ;
        RECT 32.475 -106.245 32.805 -105.915 ;
        RECT 32.475 -107.605 32.805 -107.275 ;
        RECT 32.475 -108.965 32.805 -108.635 ;
        RECT 32.475 -110.325 32.805 -109.995 ;
        RECT 32.475 -111.685 32.805 -111.355 ;
        RECT 32.475 -113.045 32.805 -112.715 ;
        RECT 32.475 -114.405 32.805 -114.075 ;
        RECT 32.475 -115.765 32.805 -115.435 ;
        RECT 32.475 -117.125 32.805 -116.795 ;
        RECT 32.475 -118.485 32.805 -118.155 ;
        RECT 32.475 -119.845 32.805 -119.515 ;
        RECT 32.475 -121.205 32.805 -120.875 ;
        RECT 32.475 -122.565 32.805 -122.235 ;
        RECT 32.475 -123.925 32.805 -123.595 ;
        RECT 32.475 -125.285 32.805 -124.955 ;
        RECT 32.475 -126.645 32.805 -126.315 ;
        RECT 32.475 -128.005 32.805 -127.675 ;
        RECT 32.475 -129.365 32.805 -129.035 ;
        RECT 32.475 -130.725 32.805 -130.395 ;
        RECT 32.475 -132.085 32.805 -131.755 ;
        RECT 32.475 -133.445 32.805 -133.115 ;
        RECT 32.475 -134.805 32.805 -134.475 ;
        RECT 32.475 -136.165 32.805 -135.835 ;
        RECT 32.475 -137.525 32.805 -137.195 ;
        RECT 32.475 -138.885 32.805 -138.555 ;
        RECT 32.475 -140.245 32.805 -139.915 ;
        RECT 32.475 -141.605 32.805 -141.275 ;
        RECT 32.475 -142.965 32.805 -142.635 ;
        RECT 32.475 -144.325 32.805 -143.995 ;
        RECT 32.475 -145.685 32.805 -145.355 ;
        RECT 32.475 -147.045 32.805 -146.715 ;
        RECT 32.475 -148.405 32.805 -148.075 ;
        RECT 32.475 -149.765 32.805 -149.435 ;
        RECT 32.475 -151.125 32.805 -150.795 ;
        RECT 32.475 -152.485 32.805 -152.155 ;
        RECT 32.475 -153.845 32.805 -153.515 ;
        RECT 32.475 -155.205 32.805 -154.875 ;
        RECT 32.475 -156.565 32.805 -156.235 ;
        RECT 32.475 -157.925 32.805 -157.595 ;
        RECT 32.475 -159.285 32.805 -158.955 ;
        RECT 32.475 -160.645 32.805 -160.315 ;
        RECT 32.475 -162.005 32.805 -161.675 ;
        RECT 32.475 -163.365 32.805 -163.035 ;
        RECT 32.475 -164.725 32.805 -164.395 ;
        RECT 32.475 -166.085 32.805 -165.755 ;
        RECT 32.475 -167.445 32.805 -167.115 ;
        RECT 32.475 -168.805 32.805 -168.475 ;
        RECT 32.475 -170.165 32.805 -169.835 ;
        RECT 32.475 -171.525 32.805 -171.195 ;
        RECT 32.475 -172.885 32.805 -172.555 ;
        RECT 32.475 -174.245 32.805 -173.915 ;
        RECT 32.475 -175.605 32.805 -175.275 ;
        RECT 32.475 -176.965 32.805 -176.635 ;
        RECT 32.475 -178.325 32.805 -177.995 ;
        RECT 32.475 -180.57 32.805 -179.44 ;
        RECT 32.48 -180.685 32.8 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.81 -94.075 34.14 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.835 241.32 34.165 242.45 ;
        RECT 33.835 239.195 34.165 239.525 ;
        RECT 33.835 237.835 34.165 238.165 ;
        RECT 33.84 237.16 34.16 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.195 241.32 35.525 242.45 ;
        RECT 35.195 239.195 35.525 239.525 ;
        RECT 35.195 237.835 35.525 238.165 ;
        RECT 35.2 237.16 35.52 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.195 -1.525 35.525 -1.195 ;
        RECT 35.195 -2.885 35.525 -2.555 ;
        RECT 35.2 -3.56 35.52 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 36.555 241.32 36.885 242.45 ;
        RECT 36.555 239.195 36.885 239.525 ;
        RECT 36.555 237.835 36.885 238.165 ;
        RECT 36.56 237.16 36.88 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 36.555 -1.525 36.885 -1.195 ;
        RECT 36.555 -2.885 36.885 -2.555 ;
        RECT 36.56 -3.56 36.88 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.915 241.32 38.245 242.45 ;
        RECT 37.915 239.195 38.245 239.525 ;
        RECT 37.915 237.835 38.245 238.165 ;
        RECT 37.92 237.16 38.24 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.915 -1.525 38.245 -1.195 ;
        RECT 37.915 -2.885 38.245 -2.555 ;
        RECT 37.92 -3.56 38.24 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.915 -91.285 38.245 -90.955 ;
        RECT 37.915 -92.645 38.245 -92.315 ;
        RECT 37.915 -94.005 38.245 -93.675 ;
        RECT 37.915 -95.365 38.245 -95.035 ;
        RECT 37.915 -96.725 38.245 -96.395 ;
        RECT 37.915 -98.085 38.245 -97.755 ;
        RECT 37.915 -99.445 38.245 -99.115 ;
        RECT 37.915 -100.805 38.245 -100.475 ;
        RECT 37.915 -102.165 38.245 -101.835 ;
        RECT 37.915 -103.525 38.245 -103.195 ;
        RECT 37.915 -104.885 38.245 -104.555 ;
        RECT 37.915 -106.245 38.245 -105.915 ;
        RECT 37.915 -107.605 38.245 -107.275 ;
        RECT 37.915 -108.965 38.245 -108.635 ;
        RECT 37.915 -110.325 38.245 -109.995 ;
        RECT 37.915 -111.685 38.245 -111.355 ;
        RECT 37.915 -113.045 38.245 -112.715 ;
        RECT 37.915 -114.405 38.245 -114.075 ;
        RECT 37.915 -115.765 38.245 -115.435 ;
        RECT 37.915 -117.125 38.245 -116.795 ;
        RECT 37.915 -118.485 38.245 -118.155 ;
        RECT 37.915 -119.845 38.245 -119.515 ;
        RECT 37.915 -121.205 38.245 -120.875 ;
        RECT 37.915 -122.565 38.245 -122.235 ;
        RECT 37.915 -123.925 38.245 -123.595 ;
        RECT 37.915 -125.285 38.245 -124.955 ;
        RECT 37.915 -126.645 38.245 -126.315 ;
        RECT 37.915 -128.005 38.245 -127.675 ;
        RECT 37.915 -129.365 38.245 -129.035 ;
        RECT 37.915 -130.725 38.245 -130.395 ;
        RECT 37.915 -132.085 38.245 -131.755 ;
        RECT 37.915 -133.445 38.245 -133.115 ;
        RECT 37.915 -134.805 38.245 -134.475 ;
        RECT 37.915 -136.165 38.245 -135.835 ;
        RECT 37.915 -137.525 38.245 -137.195 ;
        RECT 37.915 -138.885 38.245 -138.555 ;
        RECT 37.915 -140.245 38.245 -139.915 ;
        RECT 37.915 -141.605 38.245 -141.275 ;
        RECT 37.915 -142.965 38.245 -142.635 ;
        RECT 37.915 -144.325 38.245 -143.995 ;
        RECT 37.915 -145.685 38.245 -145.355 ;
        RECT 37.915 -147.045 38.245 -146.715 ;
        RECT 37.915 -148.405 38.245 -148.075 ;
        RECT 37.915 -149.765 38.245 -149.435 ;
        RECT 37.915 -151.125 38.245 -150.795 ;
        RECT 37.915 -152.485 38.245 -152.155 ;
        RECT 37.915 -153.845 38.245 -153.515 ;
        RECT 37.915 -155.205 38.245 -154.875 ;
        RECT 37.915 -156.565 38.245 -156.235 ;
        RECT 37.915 -157.925 38.245 -157.595 ;
        RECT 37.915 -159.285 38.245 -158.955 ;
        RECT 37.915 -160.645 38.245 -160.315 ;
        RECT 37.915 -162.005 38.245 -161.675 ;
        RECT 37.915 -163.365 38.245 -163.035 ;
        RECT 37.915 -164.725 38.245 -164.395 ;
        RECT 37.915 -166.085 38.245 -165.755 ;
        RECT 37.915 -167.445 38.245 -167.115 ;
        RECT 37.915 -168.805 38.245 -168.475 ;
        RECT 37.915 -170.165 38.245 -169.835 ;
        RECT 37.915 -171.525 38.245 -171.195 ;
        RECT 37.915 -172.885 38.245 -172.555 ;
        RECT 37.915 -174.245 38.245 -173.915 ;
        RECT 37.915 -175.605 38.245 -175.275 ;
        RECT 37.915 -176.965 38.245 -176.635 ;
        RECT 37.915 -178.325 38.245 -177.995 ;
        RECT 37.915 -180.57 38.245 -179.44 ;
        RECT 37.92 -180.685 38.24 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.275 241.32 39.605 242.45 ;
        RECT 39.275 239.195 39.605 239.525 ;
        RECT 39.275 237.835 39.605 238.165 ;
        RECT 39.28 237.16 39.6 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.275 -95.365 39.605 -95.035 ;
        RECT 39.275 -96.725 39.605 -96.395 ;
        RECT 39.275 -98.085 39.605 -97.755 ;
        RECT 39.275 -99.445 39.605 -99.115 ;
        RECT 39.275 -100.805 39.605 -100.475 ;
        RECT 39.275 -102.165 39.605 -101.835 ;
        RECT 39.275 -103.525 39.605 -103.195 ;
        RECT 39.275 -104.885 39.605 -104.555 ;
        RECT 39.275 -106.245 39.605 -105.915 ;
        RECT 39.275 -107.605 39.605 -107.275 ;
        RECT 39.275 -108.965 39.605 -108.635 ;
        RECT 39.275 -110.325 39.605 -109.995 ;
        RECT 39.275 -111.685 39.605 -111.355 ;
        RECT 39.275 -113.045 39.605 -112.715 ;
        RECT 39.275 -114.405 39.605 -114.075 ;
        RECT 39.275 -115.765 39.605 -115.435 ;
        RECT 39.275 -117.125 39.605 -116.795 ;
        RECT 39.275 -118.485 39.605 -118.155 ;
        RECT 39.275 -119.845 39.605 -119.515 ;
        RECT 39.275 -121.205 39.605 -120.875 ;
        RECT 39.275 -122.565 39.605 -122.235 ;
        RECT 39.275 -123.925 39.605 -123.595 ;
        RECT 39.275 -125.285 39.605 -124.955 ;
        RECT 39.275 -126.645 39.605 -126.315 ;
        RECT 39.275 -128.005 39.605 -127.675 ;
        RECT 39.275 -129.365 39.605 -129.035 ;
        RECT 39.275 -130.725 39.605 -130.395 ;
        RECT 39.275 -132.085 39.605 -131.755 ;
        RECT 39.275 -133.445 39.605 -133.115 ;
        RECT 39.275 -134.805 39.605 -134.475 ;
        RECT 39.275 -136.165 39.605 -135.835 ;
        RECT 39.275 -137.525 39.605 -137.195 ;
        RECT 39.275 -138.885 39.605 -138.555 ;
        RECT 39.275 -140.245 39.605 -139.915 ;
        RECT 39.275 -141.605 39.605 -141.275 ;
        RECT 39.275 -142.965 39.605 -142.635 ;
        RECT 39.275 -144.325 39.605 -143.995 ;
        RECT 39.275 -145.685 39.605 -145.355 ;
        RECT 39.275 -147.045 39.605 -146.715 ;
        RECT 39.275 -148.405 39.605 -148.075 ;
        RECT 39.275 -149.765 39.605 -149.435 ;
        RECT 39.275 -151.125 39.605 -150.795 ;
        RECT 39.275 -152.485 39.605 -152.155 ;
        RECT 39.275 -153.845 39.605 -153.515 ;
        RECT 39.275 -155.205 39.605 -154.875 ;
        RECT 39.275 -156.565 39.605 -156.235 ;
        RECT 39.275 -157.925 39.605 -157.595 ;
        RECT 39.275 -159.285 39.605 -158.955 ;
        RECT 39.275 -160.645 39.605 -160.315 ;
        RECT 39.275 -162.005 39.605 -161.675 ;
        RECT 39.275 -163.365 39.605 -163.035 ;
        RECT 39.275 -164.725 39.605 -164.395 ;
        RECT 39.275 -166.085 39.605 -165.755 ;
        RECT 39.275 -167.445 39.605 -167.115 ;
        RECT 39.275 -168.805 39.605 -168.475 ;
        RECT 39.275 -170.165 39.605 -169.835 ;
        RECT 39.275 -171.525 39.605 -171.195 ;
        RECT 39.275 -172.885 39.605 -172.555 ;
        RECT 39.275 -174.245 39.605 -173.915 ;
        RECT 39.275 -175.605 39.605 -175.275 ;
        RECT 39.275 -176.965 39.605 -176.635 ;
        RECT 39.275 -178.325 39.605 -177.995 ;
        RECT 39.275 -180.57 39.605 -179.44 ;
        RECT 39.28 -180.685 39.6 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.91 -94.075 40.24 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.635 241.32 40.965 242.45 ;
        RECT 40.635 239.195 40.965 239.525 ;
        RECT 40.635 237.835 40.965 238.165 ;
        RECT 40.64 237.16 40.96 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.635 -1.525 40.965 -1.195 ;
        RECT 40.635 -2.885 40.965 -2.555 ;
        RECT 40.64 -3.56 40.96 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.995 241.32 42.325 242.45 ;
        RECT 41.995 239.195 42.325 239.525 ;
        RECT 41.995 237.835 42.325 238.165 ;
        RECT 42 237.16 42.32 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.995 -1.525 42.325 -1.195 ;
        RECT 41.995 -2.885 42.325 -2.555 ;
        RECT 42 -3.56 42.32 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 43.355 241.32 43.685 242.45 ;
        RECT 43.355 239.195 43.685 239.525 ;
        RECT 43.355 237.835 43.685 238.165 ;
        RECT 43.36 237.16 43.68 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 43.355 -1.525 43.685 -1.195 ;
        RECT 43.355 -2.885 43.685 -2.555 ;
        RECT 43.36 -3.56 43.68 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 43.355 -91.285 43.685 -90.955 ;
        RECT 43.355 -92.645 43.685 -92.315 ;
        RECT 43.355 -94.005 43.685 -93.675 ;
        RECT 43.355 -95.365 43.685 -95.035 ;
        RECT 43.355 -96.725 43.685 -96.395 ;
        RECT 43.355 -98.085 43.685 -97.755 ;
        RECT 43.355 -99.445 43.685 -99.115 ;
        RECT 43.355 -100.805 43.685 -100.475 ;
        RECT 43.355 -102.165 43.685 -101.835 ;
        RECT 43.355 -103.525 43.685 -103.195 ;
        RECT 43.355 -104.885 43.685 -104.555 ;
        RECT 43.355 -106.245 43.685 -105.915 ;
        RECT 43.355 -107.605 43.685 -107.275 ;
        RECT 43.355 -108.965 43.685 -108.635 ;
        RECT 43.355 -110.325 43.685 -109.995 ;
        RECT 43.355 -111.685 43.685 -111.355 ;
        RECT 43.355 -113.045 43.685 -112.715 ;
        RECT 43.355 -114.405 43.685 -114.075 ;
        RECT 43.355 -115.765 43.685 -115.435 ;
        RECT 43.355 -117.125 43.685 -116.795 ;
        RECT 43.355 -118.485 43.685 -118.155 ;
        RECT 43.355 -119.845 43.685 -119.515 ;
        RECT 43.355 -121.205 43.685 -120.875 ;
        RECT 43.355 -122.565 43.685 -122.235 ;
        RECT 43.355 -123.925 43.685 -123.595 ;
        RECT 43.355 -125.285 43.685 -124.955 ;
        RECT 43.355 -126.645 43.685 -126.315 ;
        RECT 43.355 -128.005 43.685 -127.675 ;
        RECT 43.355 -129.365 43.685 -129.035 ;
        RECT 43.355 -130.725 43.685 -130.395 ;
        RECT 43.355 -132.085 43.685 -131.755 ;
        RECT 43.355 -133.445 43.685 -133.115 ;
        RECT 43.355 -134.805 43.685 -134.475 ;
        RECT 43.355 -136.165 43.685 -135.835 ;
        RECT 43.355 -137.525 43.685 -137.195 ;
        RECT 43.355 -138.885 43.685 -138.555 ;
        RECT 43.355 -140.245 43.685 -139.915 ;
        RECT 43.355 -141.605 43.685 -141.275 ;
        RECT 43.355 -142.965 43.685 -142.635 ;
        RECT 43.355 -144.325 43.685 -143.995 ;
        RECT 43.355 -145.685 43.685 -145.355 ;
        RECT 43.355 -147.045 43.685 -146.715 ;
        RECT 43.355 -148.405 43.685 -148.075 ;
        RECT 43.355 -149.765 43.685 -149.435 ;
        RECT 43.355 -151.125 43.685 -150.795 ;
        RECT 43.355 -152.485 43.685 -152.155 ;
        RECT 43.355 -153.845 43.685 -153.515 ;
        RECT 43.355 -155.205 43.685 -154.875 ;
        RECT 43.355 -156.565 43.685 -156.235 ;
        RECT 43.355 -157.925 43.685 -157.595 ;
        RECT 43.355 -159.285 43.685 -158.955 ;
        RECT 43.355 -160.645 43.685 -160.315 ;
        RECT 43.355 -162.005 43.685 -161.675 ;
        RECT 43.355 -163.365 43.685 -163.035 ;
        RECT 43.355 -164.725 43.685 -164.395 ;
        RECT 43.355 -166.085 43.685 -165.755 ;
        RECT 43.355 -167.445 43.685 -167.115 ;
        RECT 43.355 -168.805 43.685 -168.475 ;
        RECT 43.355 -170.165 43.685 -169.835 ;
        RECT 43.355 -171.525 43.685 -171.195 ;
        RECT 43.355 -172.885 43.685 -172.555 ;
        RECT 43.355 -174.245 43.685 -173.915 ;
        RECT 43.355 -175.605 43.685 -175.275 ;
        RECT 43.355 -176.965 43.685 -176.635 ;
        RECT 43.355 -178.325 43.685 -177.995 ;
        RECT 43.355 -180.57 43.685 -179.44 ;
        RECT 43.36 -180.685 43.68 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.715 241.32 45.045 242.45 ;
        RECT 44.715 239.195 45.045 239.525 ;
        RECT 44.715 237.835 45.045 238.165 ;
        RECT 44.72 237.16 45.04 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.715 -95.365 45.045 -95.035 ;
        RECT 44.715 -96.725 45.045 -96.395 ;
        RECT 44.715 -98.085 45.045 -97.755 ;
        RECT 44.715 -99.445 45.045 -99.115 ;
        RECT 44.715 -100.805 45.045 -100.475 ;
        RECT 44.715 -102.165 45.045 -101.835 ;
        RECT 44.715 -103.525 45.045 -103.195 ;
        RECT 44.715 -104.885 45.045 -104.555 ;
        RECT 44.715 -106.245 45.045 -105.915 ;
        RECT 44.715 -107.605 45.045 -107.275 ;
        RECT 44.715 -108.965 45.045 -108.635 ;
        RECT 44.715 -110.325 45.045 -109.995 ;
        RECT 44.715 -111.685 45.045 -111.355 ;
        RECT 44.715 -113.045 45.045 -112.715 ;
        RECT 44.715 -114.405 45.045 -114.075 ;
        RECT 44.715 -115.765 45.045 -115.435 ;
        RECT 44.715 -117.125 45.045 -116.795 ;
        RECT 44.715 -118.485 45.045 -118.155 ;
        RECT 44.715 -119.845 45.045 -119.515 ;
        RECT 44.715 -121.205 45.045 -120.875 ;
        RECT 44.715 -122.565 45.045 -122.235 ;
        RECT 44.715 -123.925 45.045 -123.595 ;
        RECT 44.715 -125.285 45.045 -124.955 ;
        RECT 44.715 -126.645 45.045 -126.315 ;
        RECT 44.715 -128.005 45.045 -127.675 ;
        RECT 44.715 -129.365 45.045 -129.035 ;
        RECT 44.715 -130.725 45.045 -130.395 ;
        RECT 44.715 -132.085 45.045 -131.755 ;
        RECT 44.715 -133.445 45.045 -133.115 ;
        RECT 44.715 -134.805 45.045 -134.475 ;
        RECT 44.715 -136.165 45.045 -135.835 ;
        RECT 44.715 -137.525 45.045 -137.195 ;
        RECT 44.715 -138.885 45.045 -138.555 ;
        RECT 44.715 -140.245 45.045 -139.915 ;
        RECT 44.715 -141.605 45.045 -141.275 ;
        RECT 44.715 -142.965 45.045 -142.635 ;
        RECT 44.715 -144.325 45.045 -143.995 ;
        RECT 44.715 -145.685 45.045 -145.355 ;
        RECT 44.715 -147.045 45.045 -146.715 ;
        RECT 44.715 -148.405 45.045 -148.075 ;
        RECT 44.715 -149.765 45.045 -149.435 ;
        RECT 44.715 -151.125 45.045 -150.795 ;
        RECT 44.715 -152.485 45.045 -152.155 ;
        RECT 44.715 -153.845 45.045 -153.515 ;
        RECT 44.715 -155.205 45.045 -154.875 ;
        RECT 44.715 -156.565 45.045 -156.235 ;
        RECT 44.715 -157.925 45.045 -157.595 ;
        RECT 44.715 -159.285 45.045 -158.955 ;
        RECT 44.715 -160.645 45.045 -160.315 ;
        RECT 44.715 -162.005 45.045 -161.675 ;
        RECT 44.715 -163.365 45.045 -163.035 ;
        RECT 44.715 -164.725 45.045 -164.395 ;
        RECT 44.715 -166.085 45.045 -165.755 ;
        RECT 44.715 -167.445 45.045 -167.115 ;
        RECT 44.715 -168.805 45.045 -168.475 ;
        RECT 44.715 -170.165 45.045 -169.835 ;
        RECT 44.715 -171.525 45.045 -171.195 ;
        RECT 44.715 -172.885 45.045 -172.555 ;
        RECT 44.715 -174.245 45.045 -173.915 ;
        RECT 44.715 -175.605 45.045 -175.275 ;
        RECT 44.715 -176.965 45.045 -176.635 ;
        RECT 44.715 -178.325 45.045 -177.995 ;
        RECT 44.715 -180.57 45.045 -179.44 ;
        RECT 44.72 -180.685 45.04 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.01 -94.075 46.34 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.075 241.32 46.405 242.45 ;
        RECT 46.075 239.195 46.405 239.525 ;
        RECT 46.075 237.835 46.405 238.165 ;
        RECT 46.08 237.16 46.4 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.435 241.32 47.765 242.45 ;
        RECT 47.435 239.195 47.765 239.525 ;
        RECT 47.435 237.835 47.765 238.165 ;
        RECT 47.44 237.16 47.76 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.435 -1.525 47.765 -1.195 ;
        RECT 47.435 -2.885 47.765 -2.555 ;
        RECT 47.44 -3.56 47.76 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.795 241.32 49.125 242.45 ;
        RECT 48.795 239.195 49.125 239.525 ;
        RECT 48.795 237.835 49.125 238.165 ;
        RECT 48.8 237.16 49.12 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.795 -1.525 49.125 -1.195 ;
        RECT 48.795 -2.885 49.125 -2.555 ;
        RECT 48.8 -3.56 49.12 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.155 241.32 50.485 242.45 ;
        RECT 50.155 239.195 50.485 239.525 ;
        RECT 50.155 237.835 50.485 238.165 ;
        RECT 50.16 237.16 50.48 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.155 -1.525 50.485 -1.195 ;
        RECT 50.155 -2.885 50.485 -2.555 ;
        RECT 50.16 -3.56 50.48 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.155 -91.285 50.485 -90.955 ;
        RECT 50.155 -92.645 50.485 -92.315 ;
        RECT 50.155 -94.005 50.485 -93.675 ;
        RECT 50.155 -95.365 50.485 -95.035 ;
        RECT 50.155 -96.725 50.485 -96.395 ;
        RECT 50.155 -98.085 50.485 -97.755 ;
        RECT 50.155 -99.445 50.485 -99.115 ;
        RECT 50.155 -100.805 50.485 -100.475 ;
        RECT 50.155 -102.165 50.485 -101.835 ;
        RECT 50.155 -103.525 50.485 -103.195 ;
        RECT 50.155 -104.885 50.485 -104.555 ;
        RECT 50.155 -106.245 50.485 -105.915 ;
        RECT 50.155 -107.605 50.485 -107.275 ;
        RECT 50.155 -108.965 50.485 -108.635 ;
        RECT 50.155 -110.325 50.485 -109.995 ;
        RECT 50.155 -111.685 50.485 -111.355 ;
        RECT 50.155 -113.045 50.485 -112.715 ;
        RECT 50.155 -114.405 50.485 -114.075 ;
        RECT 50.155 -115.765 50.485 -115.435 ;
        RECT 50.155 -117.125 50.485 -116.795 ;
        RECT 50.155 -118.485 50.485 -118.155 ;
        RECT 50.155 -119.845 50.485 -119.515 ;
        RECT 50.155 -121.205 50.485 -120.875 ;
        RECT 50.155 -122.565 50.485 -122.235 ;
        RECT 50.155 -123.925 50.485 -123.595 ;
        RECT 50.155 -125.285 50.485 -124.955 ;
        RECT 50.155 -126.645 50.485 -126.315 ;
        RECT 50.155 -128.005 50.485 -127.675 ;
        RECT 50.155 -129.365 50.485 -129.035 ;
        RECT 50.155 -130.725 50.485 -130.395 ;
        RECT 50.155 -132.085 50.485 -131.755 ;
        RECT 50.155 -133.445 50.485 -133.115 ;
        RECT 50.155 -134.805 50.485 -134.475 ;
        RECT 50.155 -136.165 50.485 -135.835 ;
        RECT 50.155 -137.525 50.485 -137.195 ;
        RECT 50.155 -138.885 50.485 -138.555 ;
        RECT 50.155 -140.245 50.485 -139.915 ;
        RECT 50.155 -141.605 50.485 -141.275 ;
        RECT 50.155 -142.965 50.485 -142.635 ;
        RECT 50.155 -144.325 50.485 -143.995 ;
        RECT 50.155 -145.685 50.485 -145.355 ;
        RECT 50.155 -147.045 50.485 -146.715 ;
        RECT 50.155 -148.405 50.485 -148.075 ;
        RECT 50.155 -149.765 50.485 -149.435 ;
        RECT 50.155 -151.125 50.485 -150.795 ;
        RECT 50.155 -152.485 50.485 -152.155 ;
        RECT 50.155 -153.845 50.485 -153.515 ;
        RECT 50.155 -155.205 50.485 -154.875 ;
        RECT 50.155 -156.565 50.485 -156.235 ;
        RECT 50.155 -157.925 50.485 -157.595 ;
        RECT 50.155 -159.285 50.485 -158.955 ;
        RECT 50.155 -160.645 50.485 -160.315 ;
        RECT 50.155 -162.005 50.485 -161.675 ;
        RECT 50.155 -163.365 50.485 -163.035 ;
        RECT 50.155 -164.725 50.485 -164.395 ;
        RECT 50.155 -166.085 50.485 -165.755 ;
        RECT 50.155 -167.445 50.485 -167.115 ;
        RECT 50.155 -168.805 50.485 -168.475 ;
        RECT 50.155 -170.165 50.485 -169.835 ;
        RECT 50.155 -171.525 50.485 -171.195 ;
        RECT 50.155 -172.885 50.485 -172.555 ;
        RECT 50.155 -174.245 50.485 -173.915 ;
        RECT 50.155 -175.605 50.485 -175.275 ;
        RECT 50.155 -176.965 50.485 -176.635 ;
        RECT 50.155 -178.325 50.485 -177.995 ;
        RECT 50.155 -180.57 50.485 -179.44 ;
        RECT 50.16 -180.685 50.48 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.515 241.32 51.845 242.45 ;
        RECT 51.515 239.195 51.845 239.525 ;
        RECT 51.515 237.835 51.845 238.165 ;
        RECT 51.52 237.16 51.84 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.515 -95.365 51.845 -95.035 ;
        RECT 51.515 -96.725 51.845 -96.395 ;
        RECT 51.515 -98.085 51.845 -97.755 ;
        RECT 51.515 -99.445 51.845 -99.115 ;
        RECT 51.515 -100.805 51.845 -100.475 ;
        RECT 51.515 -102.165 51.845 -101.835 ;
        RECT 51.515 -103.525 51.845 -103.195 ;
        RECT 51.515 -104.885 51.845 -104.555 ;
        RECT 51.515 -106.245 51.845 -105.915 ;
        RECT 51.515 -107.605 51.845 -107.275 ;
        RECT 51.515 -108.965 51.845 -108.635 ;
        RECT 51.515 -110.325 51.845 -109.995 ;
        RECT 51.515 -111.685 51.845 -111.355 ;
        RECT 51.515 -113.045 51.845 -112.715 ;
        RECT 51.515 -114.405 51.845 -114.075 ;
        RECT 51.515 -115.765 51.845 -115.435 ;
        RECT 51.515 -117.125 51.845 -116.795 ;
        RECT 51.515 -118.485 51.845 -118.155 ;
        RECT 51.515 -119.845 51.845 -119.515 ;
        RECT 51.515 -121.205 51.845 -120.875 ;
        RECT 51.515 -122.565 51.845 -122.235 ;
        RECT 51.515 -123.925 51.845 -123.595 ;
        RECT 51.515 -125.285 51.845 -124.955 ;
        RECT 51.515 -126.645 51.845 -126.315 ;
        RECT 51.515 -128.005 51.845 -127.675 ;
        RECT 51.515 -129.365 51.845 -129.035 ;
        RECT 51.515 -130.725 51.845 -130.395 ;
        RECT 51.515 -132.085 51.845 -131.755 ;
        RECT 51.515 -133.445 51.845 -133.115 ;
        RECT 51.515 -134.805 51.845 -134.475 ;
        RECT 51.515 -136.165 51.845 -135.835 ;
        RECT 51.515 -137.525 51.845 -137.195 ;
        RECT 51.515 -138.885 51.845 -138.555 ;
        RECT 51.515 -140.245 51.845 -139.915 ;
        RECT 51.515 -141.605 51.845 -141.275 ;
        RECT 51.515 -142.965 51.845 -142.635 ;
        RECT 51.515 -144.325 51.845 -143.995 ;
        RECT 51.515 -145.685 51.845 -145.355 ;
        RECT 51.515 -147.045 51.845 -146.715 ;
        RECT 51.515 -148.405 51.845 -148.075 ;
        RECT 51.515 -149.765 51.845 -149.435 ;
        RECT 51.515 -151.125 51.845 -150.795 ;
        RECT 51.515 -152.485 51.845 -152.155 ;
        RECT 51.515 -153.845 51.845 -153.515 ;
        RECT 51.515 -155.205 51.845 -154.875 ;
        RECT 51.515 -156.565 51.845 -156.235 ;
        RECT 51.515 -157.925 51.845 -157.595 ;
        RECT 51.515 -159.285 51.845 -158.955 ;
        RECT 51.515 -160.645 51.845 -160.315 ;
        RECT 51.515 -162.005 51.845 -161.675 ;
        RECT 51.515 -163.365 51.845 -163.035 ;
        RECT 51.515 -164.725 51.845 -164.395 ;
        RECT 51.515 -166.085 51.845 -165.755 ;
        RECT 51.515 -167.445 51.845 -167.115 ;
        RECT 51.515 -168.805 51.845 -168.475 ;
        RECT 51.515 -170.165 51.845 -169.835 ;
        RECT 51.515 -171.525 51.845 -171.195 ;
        RECT 51.515 -172.885 51.845 -172.555 ;
        RECT 51.515 -174.245 51.845 -173.915 ;
        RECT 51.515 -175.605 51.845 -175.275 ;
        RECT 51.515 -176.965 51.845 -176.635 ;
        RECT 51.515 -178.325 51.845 -177.995 ;
        RECT 51.515 -180.57 51.845 -179.44 ;
        RECT 51.52 -180.685 51.84 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.11 -94.075 52.44 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.875 241.32 53.205 242.45 ;
        RECT 52.875 239.195 53.205 239.525 ;
        RECT 52.875 237.835 53.205 238.165 ;
        RECT 52.88 237.16 53.2 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.875 -1.525 53.205 -1.195 ;
        RECT 52.875 -2.885 53.205 -2.555 ;
        RECT 52.88 -3.56 53.2 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.235 241.32 54.565 242.45 ;
        RECT 54.235 239.195 54.565 239.525 ;
        RECT 54.235 237.835 54.565 238.165 ;
        RECT 54.24 237.16 54.56 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.235 -1.525 54.565 -1.195 ;
        RECT 54.235 -2.885 54.565 -2.555 ;
        RECT 54.24 -3.56 54.56 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.595 241.32 55.925 242.45 ;
        RECT 55.595 239.195 55.925 239.525 ;
        RECT 55.595 237.835 55.925 238.165 ;
        RECT 55.6 237.16 55.92 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.595 -1.525 55.925 -1.195 ;
        RECT 55.595 -2.885 55.925 -2.555 ;
        RECT 55.6 -3.56 55.92 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.955 241.32 57.285 242.45 ;
        RECT 56.955 239.195 57.285 239.525 ;
        RECT 56.955 237.835 57.285 238.165 ;
        RECT 56.96 237.16 57.28 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.955 -95.365 57.285 -95.035 ;
        RECT 56.955 -96.725 57.285 -96.395 ;
        RECT 56.955 -98.085 57.285 -97.755 ;
        RECT 56.955 -99.445 57.285 -99.115 ;
        RECT 56.955 -100.805 57.285 -100.475 ;
        RECT 56.955 -102.165 57.285 -101.835 ;
        RECT 56.955 -103.525 57.285 -103.195 ;
        RECT 56.955 -104.885 57.285 -104.555 ;
        RECT 56.955 -106.245 57.285 -105.915 ;
        RECT 56.955 -107.605 57.285 -107.275 ;
        RECT 56.955 -108.965 57.285 -108.635 ;
        RECT 56.955 -110.325 57.285 -109.995 ;
        RECT 56.955 -111.685 57.285 -111.355 ;
        RECT 56.955 -113.045 57.285 -112.715 ;
        RECT 56.955 -114.405 57.285 -114.075 ;
        RECT 56.955 -115.765 57.285 -115.435 ;
        RECT 56.955 -117.125 57.285 -116.795 ;
        RECT 56.955 -118.485 57.285 -118.155 ;
        RECT 56.955 -119.845 57.285 -119.515 ;
        RECT 56.955 -121.205 57.285 -120.875 ;
        RECT 56.955 -122.565 57.285 -122.235 ;
        RECT 56.955 -123.925 57.285 -123.595 ;
        RECT 56.955 -125.285 57.285 -124.955 ;
        RECT 56.955 -126.645 57.285 -126.315 ;
        RECT 56.955 -128.005 57.285 -127.675 ;
        RECT 56.955 -129.365 57.285 -129.035 ;
        RECT 56.955 -130.725 57.285 -130.395 ;
        RECT 56.955 -132.085 57.285 -131.755 ;
        RECT 56.955 -133.445 57.285 -133.115 ;
        RECT 56.955 -134.805 57.285 -134.475 ;
        RECT 56.955 -136.165 57.285 -135.835 ;
        RECT 56.955 -137.525 57.285 -137.195 ;
        RECT 56.955 -138.885 57.285 -138.555 ;
        RECT 56.955 -140.245 57.285 -139.915 ;
        RECT 56.955 -141.605 57.285 -141.275 ;
        RECT 56.955 -142.965 57.285 -142.635 ;
        RECT 56.955 -144.325 57.285 -143.995 ;
        RECT 56.955 -145.685 57.285 -145.355 ;
        RECT 56.955 -147.045 57.285 -146.715 ;
        RECT 56.955 -148.405 57.285 -148.075 ;
        RECT 56.955 -149.765 57.285 -149.435 ;
        RECT 56.955 -151.125 57.285 -150.795 ;
        RECT 56.955 -152.485 57.285 -152.155 ;
        RECT 56.955 -153.845 57.285 -153.515 ;
        RECT 56.955 -155.205 57.285 -154.875 ;
        RECT 56.955 -156.565 57.285 -156.235 ;
        RECT 56.955 -157.925 57.285 -157.595 ;
        RECT 56.955 -159.285 57.285 -158.955 ;
        RECT 56.955 -160.645 57.285 -160.315 ;
        RECT 56.955 -162.005 57.285 -161.675 ;
        RECT 56.955 -163.365 57.285 -163.035 ;
        RECT 56.955 -164.725 57.285 -164.395 ;
        RECT 56.955 -166.085 57.285 -165.755 ;
        RECT 56.955 -167.445 57.285 -167.115 ;
        RECT 56.955 -168.805 57.285 -168.475 ;
        RECT 56.955 -170.165 57.285 -169.835 ;
        RECT 56.955 -171.525 57.285 -171.195 ;
        RECT 56.955 -172.885 57.285 -172.555 ;
        RECT 56.955 -174.245 57.285 -173.915 ;
        RECT 56.955 -175.605 57.285 -175.275 ;
        RECT 56.955 -176.965 57.285 -176.635 ;
        RECT 56.955 -178.325 57.285 -177.995 ;
        RECT 56.955 -180.57 57.285 -179.44 ;
        RECT 56.96 -180.685 57.28 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.21 -94.075 58.54 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.315 241.32 58.645 242.45 ;
        RECT 58.315 239.195 58.645 239.525 ;
        RECT 58.315 237.835 58.645 238.165 ;
        RECT 58.32 237.16 58.64 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.675 241.32 60.005 242.45 ;
        RECT 59.675 239.195 60.005 239.525 ;
        RECT 59.675 237.835 60.005 238.165 ;
        RECT 59.68 237.16 60 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.675 -1.525 60.005 -1.195 ;
        RECT 59.675 -2.885 60.005 -2.555 ;
        RECT 59.68 -3.56 60 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.675 -91.285 60.005 -90.955 ;
        RECT 59.675 -92.645 60.005 -92.315 ;
        RECT 59.675 -94.005 60.005 -93.675 ;
        RECT 59.675 -95.365 60.005 -95.035 ;
        RECT 59.675 -96.725 60.005 -96.395 ;
        RECT 59.675 -98.085 60.005 -97.755 ;
        RECT 59.675 -99.445 60.005 -99.115 ;
        RECT 59.675 -100.805 60.005 -100.475 ;
        RECT 59.675 -102.165 60.005 -101.835 ;
        RECT 59.675 -103.525 60.005 -103.195 ;
        RECT 59.675 -104.885 60.005 -104.555 ;
        RECT 59.675 -106.245 60.005 -105.915 ;
        RECT 59.675 -107.605 60.005 -107.275 ;
        RECT 59.675 -108.965 60.005 -108.635 ;
        RECT 59.675 -110.325 60.005 -109.995 ;
        RECT 59.675 -111.685 60.005 -111.355 ;
        RECT 59.675 -113.045 60.005 -112.715 ;
        RECT 59.675 -114.405 60.005 -114.075 ;
        RECT 59.675 -115.765 60.005 -115.435 ;
        RECT 59.675 -117.125 60.005 -116.795 ;
        RECT 59.675 -118.485 60.005 -118.155 ;
        RECT 59.675 -119.845 60.005 -119.515 ;
        RECT 59.675 -121.205 60.005 -120.875 ;
        RECT 59.675 -122.565 60.005 -122.235 ;
        RECT 59.675 -123.925 60.005 -123.595 ;
        RECT 59.675 -125.285 60.005 -124.955 ;
        RECT 59.675 -126.645 60.005 -126.315 ;
        RECT 59.675 -128.005 60.005 -127.675 ;
        RECT 59.675 -129.365 60.005 -129.035 ;
        RECT 59.675 -130.725 60.005 -130.395 ;
        RECT 59.675 -132.085 60.005 -131.755 ;
        RECT 59.675 -133.445 60.005 -133.115 ;
        RECT 59.675 -134.805 60.005 -134.475 ;
        RECT 59.675 -136.165 60.005 -135.835 ;
        RECT 59.675 -137.525 60.005 -137.195 ;
        RECT 59.675 -138.885 60.005 -138.555 ;
        RECT 59.675 -140.245 60.005 -139.915 ;
        RECT 59.675 -141.605 60.005 -141.275 ;
        RECT 59.675 -142.965 60.005 -142.635 ;
        RECT 59.675 -144.325 60.005 -143.995 ;
        RECT 59.675 -145.685 60.005 -145.355 ;
        RECT 59.675 -147.045 60.005 -146.715 ;
        RECT 59.675 -148.405 60.005 -148.075 ;
        RECT 59.675 -149.765 60.005 -149.435 ;
        RECT 59.675 -151.125 60.005 -150.795 ;
        RECT 59.675 -152.485 60.005 -152.155 ;
        RECT 59.675 -153.845 60.005 -153.515 ;
        RECT 59.675 -155.205 60.005 -154.875 ;
        RECT 59.675 -156.565 60.005 -156.235 ;
        RECT 59.675 -157.925 60.005 -157.595 ;
        RECT 59.675 -159.285 60.005 -158.955 ;
        RECT 59.675 -160.645 60.005 -160.315 ;
        RECT 59.675 -162.005 60.005 -161.675 ;
        RECT 59.675 -163.365 60.005 -163.035 ;
        RECT 59.675 -164.725 60.005 -164.395 ;
        RECT 59.675 -166.085 60.005 -165.755 ;
        RECT 59.675 -167.445 60.005 -167.115 ;
        RECT 59.675 -168.805 60.005 -168.475 ;
        RECT 59.675 -170.165 60.005 -169.835 ;
        RECT 59.675 -171.525 60.005 -171.195 ;
        RECT 59.675 -172.885 60.005 -172.555 ;
        RECT 59.675 -174.245 60.005 -173.915 ;
        RECT 59.675 -175.605 60.005 -175.275 ;
        RECT 59.675 -176.965 60.005 -176.635 ;
        RECT 59.675 -178.325 60.005 -177.995 ;
        RECT 59.675 -180.57 60.005 -179.44 ;
        RECT 59.68 -180.685 60 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.035 241.32 61.365 242.45 ;
        RECT 61.035 239.195 61.365 239.525 ;
        RECT 61.035 237.835 61.365 238.165 ;
        RECT 61.04 237.16 61.36 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.035 -1.525 61.365 -1.195 ;
        RECT 61.035 -2.885 61.365 -2.555 ;
        RECT 61.04 -3.56 61.36 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.395 241.32 62.725 242.45 ;
        RECT 62.395 239.195 62.725 239.525 ;
        RECT 62.395 237.835 62.725 238.165 ;
        RECT 62.4 237.16 62.72 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.395 -1.525 62.725 -1.195 ;
        RECT 62.395 -2.885 62.725 -2.555 ;
        RECT 62.4 -3.56 62.72 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.395 -91.285 62.725 -90.955 ;
        RECT 62.395 -92.645 62.725 -92.315 ;
        RECT 62.395 -94.005 62.725 -93.675 ;
        RECT 62.395 -95.365 62.725 -95.035 ;
        RECT 62.395 -96.725 62.725 -96.395 ;
        RECT 62.395 -98.085 62.725 -97.755 ;
        RECT 62.395 -99.445 62.725 -99.115 ;
        RECT 62.395 -100.805 62.725 -100.475 ;
        RECT 62.395 -102.165 62.725 -101.835 ;
        RECT 62.395 -103.525 62.725 -103.195 ;
        RECT 62.395 -104.885 62.725 -104.555 ;
        RECT 62.395 -106.245 62.725 -105.915 ;
        RECT 62.395 -107.605 62.725 -107.275 ;
        RECT 62.395 -108.965 62.725 -108.635 ;
        RECT 62.395 -110.325 62.725 -109.995 ;
        RECT 62.395 -111.685 62.725 -111.355 ;
        RECT 62.395 -113.045 62.725 -112.715 ;
        RECT 62.395 -114.405 62.725 -114.075 ;
        RECT 62.395 -115.765 62.725 -115.435 ;
        RECT 62.395 -117.125 62.725 -116.795 ;
        RECT 62.395 -118.485 62.725 -118.155 ;
        RECT 62.395 -119.845 62.725 -119.515 ;
        RECT 62.395 -121.205 62.725 -120.875 ;
        RECT 62.395 -122.565 62.725 -122.235 ;
        RECT 62.395 -123.925 62.725 -123.595 ;
        RECT 62.395 -125.285 62.725 -124.955 ;
        RECT 62.395 -126.645 62.725 -126.315 ;
        RECT 62.395 -128.005 62.725 -127.675 ;
        RECT 62.395 -129.365 62.725 -129.035 ;
        RECT 62.395 -130.725 62.725 -130.395 ;
        RECT 62.395 -132.085 62.725 -131.755 ;
        RECT 62.395 -133.445 62.725 -133.115 ;
        RECT 62.395 -134.805 62.725 -134.475 ;
        RECT 62.395 -136.165 62.725 -135.835 ;
        RECT 62.395 -137.525 62.725 -137.195 ;
        RECT 62.395 -138.885 62.725 -138.555 ;
        RECT 62.395 -140.245 62.725 -139.915 ;
        RECT 62.395 -141.605 62.725 -141.275 ;
        RECT 62.395 -142.965 62.725 -142.635 ;
        RECT 62.395 -144.325 62.725 -143.995 ;
        RECT 62.395 -145.685 62.725 -145.355 ;
        RECT 62.395 -147.045 62.725 -146.715 ;
        RECT 62.395 -148.405 62.725 -148.075 ;
        RECT 62.395 -149.765 62.725 -149.435 ;
        RECT 62.395 -151.125 62.725 -150.795 ;
        RECT 62.395 -152.485 62.725 -152.155 ;
        RECT 62.395 -153.845 62.725 -153.515 ;
        RECT 62.395 -155.205 62.725 -154.875 ;
        RECT 62.395 -156.565 62.725 -156.235 ;
        RECT 62.395 -157.925 62.725 -157.595 ;
        RECT 62.395 -159.285 62.725 -158.955 ;
        RECT 62.395 -160.645 62.725 -160.315 ;
        RECT 62.395 -162.005 62.725 -161.675 ;
        RECT 62.395 -163.365 62.725 -163.035 ;
        RECT 62.395 -164.725 62.725 -164.395 ;
        RECT 62.395 -166.085 62.725 -165.755 ;
        RECT 62.395 -167.445 62.725 -167.115 ;
        RECT 62.395 -168.805 62.725 -168.475 ;
        RECT 62.395 -170.165 62.725 -169.835 ;
        RECT 62.395 -171.525 62.725 -171.195 ;
        RECT 62.395 -172.885 62.725 -172.555 ;
        RECT 62.395 -174.245 62.725 -173.915 ;
        RECT 62.395 -175.605 62.725 -175.275 ;
        RECT 62.395 -176.965 62.725 -176.635 ;
        RECT 62.395 -178.325 62.725 -177.995 ;
        RECT 62.395 -180.57 62.725 -179.44 ;
        RECT 62.4 -180.685 62.72 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.755 241.32 64.085 242.45 ;
        RECT 63.755 239.195 64.085 239.525 ;
        RECT 63.755 237.835 64.085 238.165 ;
        RECT 63.76 237.16 64.08 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.755 -95.365 64.085 -95.035 ;
        RECT 63.755 -96.725 64.085 -96.395 ;
        RECT 63.755 -98.085 64.085 -97.755 ;
        RECT 63.755 -99.445 64.085 -99.115 ;
        RECT 63.755 -100.805 64.085 -100.475 ;
        RECT 63.755 -102.165 64.085 -101.835 ;
        RECT 63.755 -103.525 64.085 -103.195 ;
        RECT 63.755 -104.885 64.085 -104.555 ;
        RECT 63.755 -106.245 64.085 -105.915 ;
        RECT 63.755 -107.605 64.085 -107.275 ;
        RECT 63.755 -108.965 64.085 -108.635 ;
        RECT 63.755 -110.325 64.085 -109.995 ;
        RECT 63.755 -111.685 64.085 -111.355 ;
        RECT 63.755 -113.045 64.085 -112.715 ;
        RECT 63.755 -114.405 64.085 -114.075 ;
        RECT 63.755 -115.765 64.085 -115.435 ;
        RECT 63.755 -117.125 64.085 -116.795 ;
        RECT 63.755 -118.485 64.085 -118.155 ;
        RECT 63.755 -119.845 64.085 -119.515 ;
        RECT 63.755 -121.205 64.085 -120.875 ;
        RECT 63.755 -122.565 64.085 -122.235 ;
        RECT 63.755 -123.925 64.085 -123.595 ;
        RECT 63.755 -125.285 64.085 -124.955 ;
        RECT 63.755 -126.645 64.085 -126.315 ;
        RECT 63.755 -128.005 64.085 -127.675 ;
        RECT 63.755 -129.365 64.085 -129.035 ;
        RECT 63.755 -130.725 64.085 -130.395 ;
        RECT 63.755 -132.085 64.085 -131.755 ;
        RECT 63.755 -133.445 64.085 -133.115 ;
        RECT 63.755 -134.805 64.085 -134.475 ;
        RECT 63.755 -136.165 64.085 -135.835 ;
        RECT 63.755 -137.525 64.085 -137.195 ;
        RECT 63.755 -138.885 64.085 -138.555 ;
        RECT 63.755 -140.245 64.085 -139.915 ;
        RECT 63.755 -141.605 64.085 -141.275 ;
        RECT 63.755 -142.965 64.085 -142.635 ;
        RECT 63.755 -144.325 64.085 -143.995 ;
        RECT 63.755 -145.685 64.085 -145.355 ;
        RECT 63.755 -147.045 64.085 -146.715 ;
        RECT 63.755 -148.405 64.085 -148.075 ;
        RECT 63.755 -149.765 64.085 -149.435 ;
        RECT 63.755 -151.125 64.085 -150.795 ;
        RECT 63.755 -152.485 64.085 -152.155 ;
        RECT 63.755 -153.845 64.085 -153.515 ;
        RECT 63.755 -155.205 64.085 -154.875 ;
        RECT 63.755 -156.565 64.085 -156.235 ;
        RECT 63.755 -157.925 64.085 -157.595 ;
        RECT 63.755 -159.285 64.085 -158.955 ;
        RECT 63.755 -160.645 64.085 -160.315 ;
        RECT 63.755 -162.005 64.085 -161.675 ;
        RECT 63.755 -163.365 64.085 -163.035 ;
        RECT 63.755 -164.725 64.085 -164.395 ;
        RECT 63.755 -166.085 64.085 -165.755 ;
        RECT 63.755 -167.445 64.085 -167.115 ;
        RECT 63.755 -168.805 64.085 -168.475 ;
        RECT 63.755 -170.165 64.085 -169.835 ;
        RECT 63.755 -171.525 64.085 -171.195 ;
        RECT 63.755 -172.885 64.085 -172.555 ;
        RECT 63.755 -174.245 64.085 -173.915 ;
        RECT 63.755 -175.605 64.085 -175.275 ;
        RECT 63.755 -176.965 64.085 -176.635 ;
        RECT 63.755 -178.325 64.085 -177.995 ;
        RECT 63.755 -180.57 64.085 -179.44 ;
        RECT 63.76 -180.685 64.08 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.31 -94.075 64.64 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.115 241.32 65.445 242.45 ;
        RECT 65.115 239.195 65.445 239.525 ;
        RECT 65.115 237.835 65.445 238.165 ;
        RECT 65.12 237.16 65.44 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.115 -1.525 65.445 -1.195 ;
        RECT 65.115 -2.885 65.445 -2.555 ;
        RECT 65.12 -3.56 65.44 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.475 241.32 66.805 242.45 ;
        RECT 66.475 239.195 66.805 239.525 ;
        RECT 66.475 237.835 66.805 238.165 ;
        RECT 66.48 237.16 66.8 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.475 -1.525 66.805 -1.195 ;
        RECT 66.475 -2.885 66.805 -2.555 ;
        RECT 66.48 -3.56 66.8 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.835 241.32 68.165 242.45 ;
        RECT 67.835 239.195 68.165 239.525 ;
        RECT 67.835 237.835 68.165 238.165 ;
        RECT 67.84 237.16 68.16 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.835 -1.525 68.165 -1.195 ;
        RECT 67.835 -2.885 68.165 -2.555 ;
        RECT 67.84 -3.56 68.16 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.835 -126.645 68.165 -126.315 ;
        RECT 67.835 -128.005 68.165 -127.675 ;
        RECT 67.835 -129.365 68.165 -129.035 ;
        RECT 67.835 -130.725 68.165 -130.395 ;
        RECT 67.835 -132.085 68.165 -131.755 ;
        RECT 67.835 -133.445 68.165 -133.115 ;
        RECT 67.835 -134.805 68.165 -134.475 ;
        RECT 67.835 -136.165 68.165 -135.835 ;
        RECT 67.835 -137.525 68.165 -137.195 ;
        RECT 67.835 -138.885 68.165 -138.555 ;
        RECT 67.835 -140.245 68.165 -139.915 ;
        RECT 67.835 -141.605 68.165 -141.275 ;
        RECT 67.835 -142.965 68.165 -142.635 ;
        RECT 67.835 -144.325 68.165 -143.995 ;
        RECT 67.835 -145.685 68.165 -145.355 ;
        RECT 67.835 -147.045 68.165 -146.715 ;
        RECT 67.835 -148.405 68.165 -148.075 ;
        RECT 67.835 -149.765 68.165 -149.435 ;
        RECT 67.835 -151.125 68.165 -150.795 ;
        RECT 67.835 -152.485 68.165 -152.155 ;
        RECT 67.835 -153.845 68.165 -153.515 ;
        RECT 67.835 -155.205 68.165 -154.875 ;
        RECT 67.835 -156.565 68.165 -156.235 ;
        RECT 67.835 -157.925 68.165 -157.595 ;
        RECT 67.835 -159.285 68.165 -158.955 ;
        RECT 67.835 -160.645 68.165 -160.315 ;
        RECT 67.835 -162.005 68.165 -161.675 ;
        RECT 67.835 -163.365 68.165 -163.035 ;
        RECT 67.835 -164.725 68.165 -164.395 ;
        RECT 67.835 -166.085 68.165 -165.755 ;
        RECT 67.835 -167.445 68.165 -167.115 ;
        RECT 67.835 -168.805 68.165 -168.475 ;
        RECT 67.835 -170.165 68.165 -169.835 ;
        RECT 67.835 -171.525 68.165 -171.195 ;
        RECT 67.835 -172.885 68.165 -172.555 ;
        RECT 67.835 -174.245 68.165 -173.915 ;
        RECT 67.835 -175.605 68.165 -175.275 ;
        RECT 67.835 -176.965 68.165 -176.635 ;
        RECT 67.835 -178.325 68.165 -177.995 ;
        RECT 67.835 -180.57 68.165 -179.44 ;
        RECT 67.84 -180.685 68.16 -90.955 ;
        RECT 67.835 -91.285 68.165 -90.955 ;
        RECT 67.835 -92.645 68.165 -92.315 ;
        RECT 67.835 -94.005 68.165 -93.675 ;
        RECT 67.835 -95.365 68.165 -95.035 ;
        RECT 67.835 -96.725 68.165 -96.395 ;
        RECT 67.835 -98.085 68.165 -97.755 ;
        RECT 67.835 -99.445 68.165 -99.115 ;
        RECT 67.835 -100.805 68.165 -100.475 ;
        RECT 67.835 -102.165 68.165 -101.835 ;
        RECT 67.835 -103.525 68.165 -103.195 ;
        RECT 67.835 -104.885 68.165 -104.555 ;
        RECT 67.835 -106.245 68.165 -105.915 ;
        RECT 67.835 -107.605 68.165 -107.275 ;
        RECT 67.835 -108.965 68.165 -108.635 ;
        RECT 67.835 -110.325 68.165 -109.995 ;
        RECT 67.835 -111.685 68.165 -111.355 ;
        RECT 67.835 -113.045 68.165 -112.715 ;
        RECT 67.835 -114.405 68.165 -114.075 ;
        RECT 67.835 -115.765 68.165 -115.435 ;
        RECT 67.835 -117.125 68.165 -116.795 ;
        RECT 67.835 -118.485 68.165 -118.155 ;
        RECT 67.835 -119.845 68.165 -119.515 ;
        RECT 67.835 -121.205 68.165 -120.875 ;
        RECT 67.835 -122.565 68.165 -122.235 ;
        RECT 67.835 -123.925 68.165 -123.595 ;
        RECT 67.835 -125.285 68.165 -124.955 ;
    END
    PORT
      LAYER met3 ;
        RECT -0.165 241.32 0.165 242.45 ;
        RECT -0.165 239.195 0.165 239.525 ;
        RECT -0.165 237.835 0.165 238.165 ;
        RECT -0.16 237.16 0.16 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -0.165 -1.525 0.165 -1.195 ;
        RECT -0.165 -2.885 0.165 -2.555 ;
        RECT -0.16 -3.56 0.16 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT -0.165 -91.285 0.165 -90.955 ;
        RECT -0.165 -92.645 0.165 -92.315 ;
        RECT -0.165 -94.005 0.165 -93.675 ;
        RECT -0.165 -95.365 0.165 -95.035 ;
        RECT -0.165 -96.725 0.165 -96.395 ;
        RECT -0.165 -98.085 0.165 -97.755 ;
        RECT -0.165 -99.445 0.165 -99.115 ;
        RECT -0.165 -100.805 0.165 -100.475 ;
        RECT -0.165 -102.165 0.165 -101.835 ;
        RECT -0.165 -103.525 0.165 -103.195 ;
        RECT -0.165 -104.885 0.165 -104.555 ;
        RECT -0.165 -106.245 0.165 -105.915 ;
        RECT -0.165 -107.605 0.165 -107.275 ;
        RECT -0.165 -108.965 0.165 -108.635 ;
        RECT -0.165 -110.325 0.165 -109.995 ;
        RECT -0.165 -111.685 0.165 -111.355 ;
        RECT -0.165 -113.045 0.165 -112.715 ;
        RECT -0.165 -114.405 0.165 -114.075 ;
        RECT -0.165 -115.765 0.165 -115.435 ;
        RECT -0.165 -117.125 0.165 -116.795 ;
        RECT -0.165 -119.845 0.165 -119.515 ;
        RECT -0.165 -121.205 0.165 -120.875 ;
        RECT -0.165 -122.565 0.165 -122.235 ;
        RECT -0.165 -123.925 0.165 -123.595 ;
        RECT -0.165 -125.285 0.165 -124.955 ;
        RECT -0.165 -126.645 0.165 -126.315 ;
        RECT -0.165 -128.005 0.165 -127.675 ;
        RECT -0.165 -129.365 0.165 -129.035 ;
        RECT -0.165 -130.725 0.165 -130.395 ;
        RECT -0.165 -132.085 0.165 -131.755 ;
        RECT -0.165 -133.445 0.165 -133.115 ;
        RECT -0.165 -134.805 0.165 -134.475 ;
        RECT -0.165 -136.165 0.165 -135.835 ;
        RECT -0.165 -137.525 0.165 -137.195 ;
        RECT -0.165 -138.885 0.165 -138.555 ;
        RECT -0.165 -140.245 0.165 -139.915 ;
        RECT -0.165 -141.605 0.165 -141.275 ;
        RECT -0.165 -142.965 0.165 -142.635 ;
        RECT -0.165 -144.325 0.165 -143.995 ;
        RECT -0.165 -145.685 0.165 -145.355 ;
        RECT -0.165 -147.045 0.165 -146.715 ;
        RECT -0.165 -148.405 0.165 -148.075 ;
        RECT -0.165 -149.765 0.165 -149.435 ;
        RECT -0.165 -151.125 0.165 -150.795 ;
        RECT -0.165 -152.485 0.165 -152.155 ;
        RECT -0.165 -153.845 0.165 -153.515 ;
        RECT -0.165 -155.205 0.165 -154.875 ;
        RECT -0.165 -156.565 0.165 -156.235 ;
        RECT -0.165 -157.925 0.165 -157.595 ;
        RECT -0.165 -159.285 0.165 -158.955 ;
        RECT -0.165 -160.645 0.165 -160.315 ;
        RECT -0.165 -162.005 0.165 -161.675 ;
        RECT -0.165 -163.365 0.165 -163.035 ;
        RECT -0.165 -164.725 0.165 -164.395 ;
        RECT -0.165 -166.085 0.165 -165.755 ;
        RECT -0.165 -167.445 0.165 -167.115 ;
        RECT -0.165 -168.805 0.165 -168.475 ;
        RECT -0.165 -170.165 0.165 -169.835 ;
        RECT -0.165 -171.525 0.165 -171.195 ;
        RECT -0.165 -172.885 0.165 -172.555 ;
        RECT -0.165 -174.245 0.165 -173.915 ;
        RECT -0.165 -175.605 0.165 -175.275 ;
        RECT -0.165 -176.965 0.165 -176.635 ;
        RECT -0.165 -178.325 0.165 -177.995 ;
        RECT -0.165 -180.57 0.165 -179.44 ;
        RECT -0.16 -180.685 0.16 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.195 241.32 1.525 242.45 ;
        RECT 1.195 239.195 1.525 239.525 ;
        RECT 1.195 237.835 1.525 238.165 ;
        RECT 1.2 237.16 1.52 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.195 -1.525 1.525 -1.195 ;
        RECT 1.195 -2.885 1.525 -2.555 ;
        RECT 1.2 -3.56 1.52 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.195 -91.285 1.525 -90.955 ;
        RECT 1.195 -92.645 1.525 -92.315 ;
        RECT 1.195 -94.005 1.525 -93.675 ;
        RECT 1.195 -95.365 1.525 -95.035 ;
        RECT 1.195 -96.725 1.525 -96.395 ;
        RECT 1.195 -98.085 1.525 -97.755 ;
        RECT 1.195 -99.445 1.525 -99.115 ;
        RECT 1.195 -100.805 1.525 -100.475 ;
        RECT 1.195 -102.165 1.525 -101.835 ;
        RECT 1.195 -103.525 1.525 -103.195 ;
        RECT 1.195 -104.885 1.525 -104.555 ;
        RECT 1.195 -106.245 1.525 -105.915 ;
        RECT 1.195 -107.605 1.525 -107.275 ;
        RECT 1.195 -108.965 1.525 -108.635 ;
        RECT 1.195 -110.325 1.525 -109.995 ;
        RECT 1.195 -111.685 1.525 -111.355 ;
        RECT 1.195 -113.045 1.525 -112.715 ;
        RECT 1.195 -114.405 1.525 -114.075 ;
        RECT 1.195 -115.765 1.525 -115.435 ;
        RECT 1.195 -117.125 1.525 -116.795 ;
        RECT 1.195 -118.485 1.525 -118.155 ;
        RECT 1.195 -119.845 1.525 -119.515 ;
        RECT 1.195 -121.205 1.525 -120.875 ;
        RECT 1.195 -122.565 1.525 -122.235 ;
        RECT 1.195 -123.925 1.525 -123.595 ;
        RECT 1.195 -125.285 1.525 -124.955 ;
        RECT 1.195 -126.645 1.525 -126.315 ;
        RECT 1.195 -128.005 1.525 -127.675 ;
        RECT 1.195 -129.365 1.525 -129.035 ;
        RECT 1.195 -130.725 1.525 -130.395 ;
        RECT 1.195 -132.085 1.525 -131.755 ;
        RECT 1.195 -133.445 1.525 -133.115 ;
        RECT 1.195 -134.805 1.525 -134.475 ;
        RECT 1.195 -136.165 1.525 -135.835 ;
        RECT 1.195 -137.525 1.525 -137.195 ;
        RECT 1.195 -138.885 1.525 -138.555 ;
        RECT 1.195 -140.245 1.525 -139.915 ;
        RECT 1.195 -141.605 1.525 -141.275 ;
        RECT 1.195 -142.965 1.525 -142.635 ;
        RECT 1.195 -144.325 1.525 -143.995 ;
        RECT 1.195 -145.685 1.525 -145.355 ;
        RECT 1.195 -147.045 1.525 -146.715 ;
        RECT 1.195 -148.405 1.525 -148.075 ;
        RECT 1.195 -149.765 1.525 -149.435 ;
        RECT 1.195 -151.125 1.525 -150.795 ;
        RECT 1.195 -152.485 1.525 -152.155 ;
        RECT 1.195 -153.845 1.525 -153.515 ;
        RECT 1.195 -155.205 1.525 -154.875 ;
        RECT 1.195 -156.565 1.525 -156.235 ;
        RECT 1.195 -157.925 1.525 -157.595 ;
        RECT 1.195 -159.285 1.525 -158.955 ;
        RECT 1.195 -160.645 1.525 -160.315 ;
        RECT 1.195 -162.005 1.525 -161.675 ;
        RECT 1.195 -163.365 1.525 -163.035 ;
        RECT 1.195 -164.725 1.525 -164.395 ;
        RECT 1.195 -166.085 1.525 -165.755 ;
        RECT 1.195 -167.445 1.525 -167.115 ;
        RECT 1.195 -168.805 1.525 -168.475 ;
        RECT 1.195 -170.165 1.525 -169.835 ;
        RECT 1.195 -171.525 1.525 -171.195 ;
        RECT 1.195 -172.885 1.525 -172.555 ;
        RECT 1.195 -174.245 1.525 -173.915 ;
        RECT 1.195 -175.605 1.525 -175.275 ;
        RECT 1.195 -176.965 1.525 -176.635 ;
        RECT 1.195 -178.325 1.525 -177.995 ;
        RECT 1.195 -180.57 1.525 -179.44 ;
        RECT 1.2 -180.685 1.52 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 241.32 2.885 242.45 ;
        RECT 2.555 239.195 2.885 239.525 ;
        RECT 2.555 237.835 2.885 238.165 ;
        RECT 2.56 237.16 2.88 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 -95.365 2.885 -95.035 ;
        RECT 2.555 -96.725 2.885 -96.395 ;
        RECT 2.555 -98.085 2.885 -97.755 ;
        RECT 2.555 -99.445 2.885 -99.115 ;
        RECT 2.555 -100.805 2.885 -100.475 ;
        RECT 2.555 -102.165 2.885 -101.835 ;
        RECT 2.555 -103.525 2.885 -103.195 ;
        RECT 2.555 -104.885 2.885 -104.555 ;
        RECT 2.555 -106.245 2.885 -105.915 ;
        RECT 2.555 -107.605 2.885 -107.275 ;
        RECT 2.555 -108.965 2.885 -108.635 ;
        RECT 2.555 -110.325 2.885 -109.995 ;
        RECT 2.555 -111.685 2.885 -111.355 ;
        RECT 2.555 -113.045 2.885 -112.715 ;
        RECT 2.555 -114.405 2.885 -114.075 ;
        RECT 2.555 -115.765 2.885 -115.435 ;
        RECT 2.555 -117.125 2.885 -116.795 ;
        RECT 2.555 -118.485 2.885 -118.155 ;
        RECT 2.555 -119.845 2.885 -119.515 ;
        RECT 2.555 -121.205 2.885 -120.875 ;
        RECT 2.555 -122.565 2.885 -122.235 ;
        RECT 2.555 -123.925 2.885 -123.595 ;
        RECT 2.555 -125.285 2.885 -124.955 ;
        RECT 2.555 -126.645 2.885 -126.315 ;
        RECT 2.555 -128.005 2.885 -127.675 ;
        RECT 2.555 -129.365 2.885 -129.035 ;
        RECT 2.555 -130.725 2.885 -130.395 ;
        RECT 2.555 -132.085 2.885 -131.755 ;
        RECT 2.555 -133.445 2.885 -133.115 ;
        RECT 2.555 -134.805 2.885 -134.475 ;
        RECT 2.555 -136.165 2.885 -135.835 ;
        RECT 2.555 -137.525 2.885 -137.195 ;
        RECT 2.555 -138.885 2.885 -138.555 ;
        RECT 2.555 -140.245 2.885 -139.915 ;
        RECT 2.555 -141.605 2.885 -141.275 ;
        RECT 2.555 -142.965 2.885 -142.635 ;
        RECT 2.555 -144.325 2.885 -143.995 ;
        RECT 2.555 -145.685 2.885 -145.355 ;
        RECT 2.555 -147.045 2.885 -146.715 ;
        RECT 2.555 -148.405 2.885 -148.075 ;
        RECT 2.555 -149.765 2.885 -149.435 ;
        RECT 2.555 -151.125 2.885 -150.795 ;
        RECT 2.555 -152.485 2.885 -152.155 ;
        RECT 2.555 -153.845 2.885 -153.515 ;
        RECT 2.555 -155.205 2.885 -154.875 ;
        RECT 2.555 -156.565 2.885 -156.235 ;
        RECT 2.555 -157.925 2.885 -157.595 ;
        RECT 2.555 -159.285 2.885 -158.955 ;
        RECT 2.555 -160.645 2.885 -160.315 ;
        RECT 2.555 -162.005 2.885 -161.675 ;
        RECT 2.555 -163.365 2.885 -163.035 ;
        RECT 2.555 -164.725 2.885 -164.395 ;
        RECT 2.555 -166.085 2.885 -165.755 ;
        RECT 2.555 -167.445 2.885 -167.115 ;
        RECT 2.555 -168.805 2.885 -168.475 ;
        RECT 2.555 -170.165 2.885 -169.835 ;
        RECT 2.555 -171.525 2.885 -171.195 ;
        RECT 2.555 -172.885 2.885 -172.555 ;
        RECT 2.555 -174.245 2.885 -173.915 ;
        RECT 2.555 -175.605 2.885 -175.275 ;
        RECT 2.555 -176.965 2.885 -176.635 ;
        RECT 2.555 -178.325 2.885 -177.995 ;
        RECT 2.555 -180.57 2.885 -179.44 ;
        RECT 2.56 -180.685 2.88 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.31 -94.075 3.64 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.915 241.32 4.245 242.45 ;
        RECT 3.915 239.195 4.245 239.525 ;
        RECT 3.915 237.835 4.245 238.165 ;
        RECT 3.92 237.16 4.24 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.275 241.32 5.605 242.45 ;
        RECT 5.275 239.195 5.605 239.525 ;
        RECT 5.275 237.835 5.605 238.165 ;
        RECT 5.28 237.16 5.6 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.275 -1.525 5.605 -1.195 ;
        RECT 5.275 -2.885 5.605 -2.555 ;
        RECT 5.28 -3.56 5.6 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635 241.32 6.965 242.45 ;
        RECT 6.635 239.195 6.965 239.525 ;
        RECT 6.635 237.835 6.965 238.165 ;
        RECT 6.64 237.16 6.96 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635 -1.525 6.965 -1.195 ;
        RECT 6.635 -2.885 6.965 -2.555 ;
        RECT 6.64 -3.56 6.96 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.995 241.32 8.325 242.45 ;
        RECT 7.995 239.195 8.325 239.525 ;
        RECT 7.995 237.835 8.325 238.165 ;
        RECT 8 237.16 8.32 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.995 -1.525 8.325 -1.195 ;
        RECT 7.995 -2.885 8.325 -2.555 ;
        RECT 8 -3.56 8.32 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.995 -91.285 8.325 -90.955 ;
        RECT 7.995 -92.645 8.325 -92.315 ;
        RECT 7.995 -94.005 8.325 -93.675 ;
        RECT 7.995 -95.365 8.325 -95.035 ;
        RECT 7.995 -96.725 8.325 -96.395 ;
        RECT 7.995 -98.085 8.325 -97.755 ;
        RECT 7.995 -99.445 8.325 -99.115 ;
        RECT 7.995 -100.805 8.325 -100.475 ;
        RECT 7.995 -102.165 8.325 -101.835 ;
        RECT 7.995 -103.525 8.325 -103.195 ;
        RECT 7.995 -104.885 8.325 -104.555 ;
        RECT 7.995 -106.245 8.325 -105.915 ;
        RECT 7.995 -107.605 8.325 -107.275 ;
        RECT 7.995 -108.965 8.325 -108.635 ;
        RECT 7.995 -110.325 8.325 -109.995 ;
        RECT 7.995 -111.685 8.325 -111.355 ;
        RECT 7.995 -113.045 8.325 -112.715 ;
        RECT 7.995 -114.405 8.325 -114.075 ;
        RECT 7.995 -115.765 8.325 -115.435 ;
        RECT 7.995 -117.125 8.325 -116.795 ;
        RECT 7.995 -118.485 8.325 -118.155 ;
        RECT 7.995 -119.845 8.325 -119.515 ;
        RECT 7.995 -121.205 8.325 -120.875 ;
        RECT 7.995 -122.565 8.325 -122.235 ;
        RECT 7.995 -123.925 8.325 -123.595 ;
        RECT 7.995 -125.285 8.325 -124.955 ;
        RECT 7.995 -126.645 8.325 -126.315 ;
        RECT 7.995 -128.005 8.325 -127.675 ;
        RECT 7.995 -129.365 8.325 -129.035 ;
        RECT 7.995 -130.725 8.325 -130.395 ;
        RECT 7.995 -132.085 8.325 -131.755 ;
        RECT 7.995 -133.445 8.325 -133.115 ;
        RECT 7.995 -134.805 8.325 -134.475 ;
        RECT 7.995 -136.165 8.325 -135.835 ;
        RECT 7.995 -137.525 8.325 -137.195 ;
        RECT 7.995 -138.885 8.325 -138.555 ;
        RECT 7.995 -140.245 8.325 -139.915 ;
        RECT 7.995 -141.605 8.325 -141.275 ;
        RECT 7.995 -142.965 8.325 -142.635 ;
        RECT 7.995 -144.325 8.325 -143.995 ;
        RECT 7.995 -145.685 8.325 -145.355 ;
        RECT 7.995 -147.045 8.325 -146.715 ;
        RECT 7.995 -148.405 8.325 -148.075 ;
        RECT 7.995 -149.765 8.325 -149.435 ;
        RECT 7.995 -151.125 8.325 -150.795 ;
        RECT 7.995 -152.485 8.325 -152.155 ;
        RECT 7.995 -153.845 8.325 -153.515 ;
        RECT 7.995 -155.205 8.325 -154.875 ;
        RECT 7.995 -156.565 8.325 -156.235 ;
        RECT 7.995 -157.925 8.325 -157.595 ;
        RECT 7.995 -159.285 8.325 -158.955 ;
        RECT 7.995 -160.645 8.325 -160.315 ;
        RECT 7.995 -162.005 8.325 -161.675 ;
        RECT 7.995 -163.365 8.325 -163.035 ;
        RECT 7.995 -164.725 8.325 -164.395 ;
        RECT 7.995 -166.085 8.325 -165.755 ;
        RECT 7.995 -167.445 8.325 -167.115 ;
        RECT 7.995 -168.805 8.325 -168.475 ;
        RECT 7.995 -170.165 8.325 -169.835 ;
        RECT 7.995 -171.525 8.325 -171.195 ;
        RECT 7.995 -172.885 8.325 -172.555 ;
        RECT 7.995 -174.245 8.325 -173.915 ;
        RECT 7.995 -175.605 8.325 -175.275 ;
        RECT 7.995 -176.965 8.325 -176.635 ;
        RECT 7.995 -178.325 8.325 -177.995 ;
        RECT 7.995 -180.57 8.325 -179.44 ;
        RECT 8 -180.685 8.32 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 241.32 9.685 242.45 ;
        RECT 9.355 239.195 9.685 239.525 ;
        RECT 9.355 237.835 9.685 238.165 ;
        RECT 9.36 237.16 9.68 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 -95.365 9.685 -95.035 ;
        RECT 9.355 -96.725 9.685 -96.395 ;
        RECT 9.355 -98.085 9.685 -97.755 ;
        RECT 9.355 -99.445 9.685 -99.115 ;
        RECT 9.355 -100.805 9.685 -100.475 ;
        RECT 9.355 -102.165 9.685 -101.835 ;
        RECT 9.355 -103.525 9.685 -103.195 ;
        RECT 9.355 -104.885 9.685 -104.555 ;
        RECT 9.355 -106.245 9.685 -105.915 ;
        RECT 9.355 -107.605 9.685 -107.275 ;
        RECT 9.355 -108.965 9.685 -108.635 ;
        RECT 9.355 -110.325 9.685 -109.995 ;
        RECT 9.355 -111.685 9.685 -111.355 ;
        RECT 9.355 -113.045 9.685 -112.715 ;
        RECT 9.355 -114.405 9.685 -114.075 ;
        RECT 9.355 -115.765 9.685 -115.435 ;
        RECT 9.355 -117.125 9.685 -116.795 ;
        RECT 9.355 -118.485 9.685 -118.155 ;
        RECT 9.355 -119.845 9.685 -119.515 ;
        RECT 9.355 -121.205 9.685 -120.875 ;
        RECT 9.355 -122.565 9.685 -122.235 ;
        RECT 9.355 -123.925 9.685 -123.595 ;
        RECT 9.355 -125.285 9.685 -124.955 ;
        RECT 9.355 -126.645 9.685 -126.315 ;
        RECT 9.355 -128.005 9.685 -127.675 ;
        RECT 9.355 -129.365 9.685 -129.035 ;
        RECT 9.355 -130.725 9.685 -130.395 ;
        RECT 9.355 -132.085 9.685 -131.755 ;
        RECT 9.355 -133.445 9.685 -133.115 ;
        RECT 9.355 -134.805 9.685 -134.475 ;
        RECT 9.355 -136.165 9.685 -135.835 ;
        RECT 9.355 -137.525 9.685 -137.195 ;
        RECT 9.355 -138.885 9.685 -138.555 ;
        RECT 9.355 -140.245 9.685 -139.915 ;
        RECT 9.355 -141.605 9.685 -141.275 ;
        RECT 9.355 -142.965 9.685 -142.635 ;
        RECT 9.355 -144.325 9.685 -143.995 ;
        RECT 9.355 -145.685 9.685 -145.355 ;
        RECT 9.355 -147.045 9.685 -146.715 ;
        RECT 9.355 -148.405 9.685 -148.075 ;
        RECT 9.355 -149.765 9.685 -149.435 ;
        RECT 9.355 -151.125 9.685 -150.795 ;
        RECT 9.355 -152.485 9.685 -152.155 ;
        RECT 9.355 -153.845 9.685 -153.515 ;
        RECT 9.355 -155.205 9.685 -154.875 ;
        RECT 9.355 -156.565 9.685 -156.235 ;
        RECT 9.355 -157.925 9.685 -157.595 ;
        RECT 9.355 -159.285 9.685 -158.955 ;
        RECT 9.355 -160.645 9.685 -160.315 ;
        RECT 9.355 -162.005 9.685 -161.675 ;
        RECT 9.355 -163.365 9.685 -163.035 ;
        RECT 9.355 -164.725 9.685 -164.395 ;
        RECT 9.355 -166.085 9.685 -165.755 ;
        RECT 9.355 -167.445 9.685 -167.115 ;
        RECT 9.355 -168.805 9.685 -168.475 ;
        RECT 9.355 -170.165 9.685 -169.835 ;
        RECT 9.355 -171.525 9.685 -171.195 ;
        RECT 9.355 -172.885 9.685 -172.555 ;
        RECT 9.355 -174.245 9.685 -173.915 ;
        RECT 9.355 -175.605 9.685 -175.275 ;
        RECT 9.355 -176.965 9.685 -176.635 ;
        RECT 9.355 -178.325 9.685 -177.995 ;
        RECT 9.355 -180.57 9.685 -179.44 ;
        RECT 9.36 -180.685 9.68 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.41 -94.075 9.74 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.715 241.32 11.045 242.45 ;
        RECT 10.715 239.195 11.045 239.525 ;
        RECT 10.715 237.835 11.045 238.165 ;
        RECT 10.72 237.16 11.04 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.715 -1.525 11.045 -1.195 ;
        RECT 10.715 -2.885 11.045 -2.555 ;
        RECT 10.72 -3.56 11.04 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.075 241.32 12.405 242.45 ;
        RECT 12.075 239.195 12.405 239.525 ;
        RECT 12.075 237.835 12.405 238.165 ;
        RECT 12.08 237.16 12.4 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.075 -1.525 12.405 -1.195 ;
        RECT 12.075 -2.885 12.405 -2.555 ;
        RECT 12.08 -3.56 12.4 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.435 241.32 13.765 242.45 ;
        RECT 13.435 239.195 13.765 239.525 ;
        RECT 13.435 237.835 13.765 238.165 ;
        RECT 13.44 237.16 13.76 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.435 -1.525 13.765 -1.195 ;
        RECT 13.435 -2.885 13.765 -2.555 ;
        RECT 13.44 -3.56 13.76 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.435 -91.285 13.765 -90.955 ;
        RECT 13.435 -92.645 13.765 -92.315 ;
        RECT 13.435 -94.005 13.765 -93.675 ;
        RECT 13.435 -95.365 13.765 -95.035 ;
        RECT 13.435 -96.725 13.765 -96.395 ;
        RECT 13.435 -98.085 13.765 -97.755 ;
        RECT 13.435 -99.445 13.765 -99.115 ;
        RECT 13.435 -100.805 13.765 -100.475 ;
        RECT 13.435 -102.165 13.765 -101.835 ;
        RECT 13.435 -103.525 13.765 -103.195 ;
        RECT 13.435 -104.885 13.765 -104.555 ;
        RECT 13.435 -106.245 13.765 -105.915 ;
        RECT 13.435 -107.605 13.765 -107.275 ;
        RECT 13.435 -108.965 13.765 -108.635 ;
        RECT 13.435 -110.325 13.765 -109.995 ;
        RECT 13.435 -111.685 13.765 -111.355 ;
        RECT 13.435 -113.045 13.765 -112.715 ;
        RECT 13.435 -114.405 13.765 -114.075 ;
        RECT 13.435 -115.765 13.765 -115.435 ;
        RECT 13.435 -117.125 13.765 -116.795 ;
        RECT 13.435 -118.485 13.765 -118.155 ;
        RECT 13.435 -119.845 13.765 -119.515 ;
        RECT 13.435 -121.205 13.765 -120.875 ;
        RECT 13.435 -122.565 13.765 -122.235 ;
        RECT 13.435 -123.925 13.765 -123.595 ;
        RECT 13.435 -125.285 13.765 -124.955 ;
        RECT 13.435 -126.645 13.765 -126.315 ;
        RECT 13.435 -128.005 13.765 -127.675 ;
        RECT 13.435 -129.365 13.765 -129.035 ;
        RECT 13.435 -130.725 13.765 -130.395 ;
        RECT 13.435 -132.085 13.765 -131.755 ;
        RECT 13.435 -133.445 13.765 -133.115 ;
        RECT 13.435 -134.805 13.765 -134.475 ;
        RECT 13.435 -136.165 13.765 -135.835 ;
        RECT 13.435 -137.525 13.765 -137.195 ;
        RECT 13.435 -138.885 13.765 -138.555 ;
        RECT 13.435 -140.245 13.765 -139.915 ;
        RECT 13.435 -141.605 13.765 -141.275 ;
        RECT 13.435 -142.965 13.765 -142.635 ;
        RECT 13.435 -144.325 13.765 -143.995 ;
        RECT 13.435 -145.685 13.765 -145.355 ;
        RECT 13.435 -147.045 13.765 -146.715 ;
        RECT 13.435 -148.405 13.765 -148.075 ;
        RECT 13.435 -149.765 13.765 -149.435 ;
        RECT 13.435 -151.125 13.765 -150.795 ;
        RECT 13.435 -152.485 13.765 -152.155 ;
        RECT 13.435 -153.845 13.765 -153.515 ;
        RECT 13.435 -155.205 13.765 -154.875 ;
        RECT 13.435 -156.565 13.765 -156.235 ;
        RECT 13.435 -157.925 13.765 -157.595 ;
        RECT 13.435 -159.285 13.765 -158.955 ;
        RECT 13.435 -160.645 13.765 -160.315 ;
        RECT 13.435 -162.005 13.765 -161.675 ;
        RECT 13.435 -163.365 13.765 -163.035 ;
        RECT 13.435 -164.725 13.765 -164.395 ;
        RECT 13.435 -166.085 13.765 -165.755 ;
        RECT 13.435 -167.445 13.765 -167.115 ;
        RECT 13.435 -168.805 13.765 -168.475 ;
        RECT 13.435 -170.165 13.765 -169.835 ;
        RECT 13.435 -171.525 13.765 -171.195 ;
        RECT 13.435 -172.885 13.765 -172.555 ;
        RECT 13.435 -174.245 13.765 -173.915 ;
        RECT 13.435 -175.605 13.765 -175.275 ;
        RECT 13.435 -176.965 13.765 -176.635 ;
        RECT 13.435 -178.325 13.765 -177.995 ;
        RECT 13.435 -180.57 13.765 -179.44 ;
        RECT 13.44 -180.685 13.76 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.795 241.32 15.125 242.45 ;
        RECT 14.795 239.195 15.125 239.525 ;
        RECT 14.795 237.835 15.125 238.165 ;
        RECT 14.8 237.16 15.12 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.795 -95.365 15.125 -95.035 ;
        RECT 14.795 -96.725 15.125 -96.395 ;
        RECT 14.795 -98.085 15.125 -97.755 ;
        RECT 14.795 -99.445 15.125 -99.115 ;
        RECT 14.795 -100.805 15.125 -100.475 ;
        RECT 14.795 -102.165 15.125 -101.835 ;
        RECT 14.795 -103.525 15.125 -103.195 ;
        RECT 14.795 -104.885 15.125 -104.555 ;
        RECT 14.795 -106.245 15.125 -105.915 ;
        RECT 14.795 -107.605 15.125 -107.275 ;
        RECT 14.795 -108.965 15.125 -108.635 ;
        RECT 14.795 -110.325 15.125 -109.995 ;
        RECT 14.795 -111.685 15.125 -111.355 ;
        RECT 14.795 -113.045 15.125 -112.715 ;
        RECT 14.795 -114.405 15.125 -114.075 ;
        RECT 14.795 -115.765 15.125 -115.435 ;
        RECT 14.795 -117.125 15.125 -116.795 ;
        RECT 14.795 -118.485 15.125 -118.155 ;
        RECT 14.795 -119.845 15.125 -119.515 ;
        RECT 14.795 -121.205 15.125 -120.875 ;
        RECT 14.795 -122.565 15.125 -122.235 ;
        RECT 14.795 -123.925 15.125 -123.595 ;
        RECT 14.795 -125.285 15.125 -124.955 ;
        RECT 14.795 -126.645 15.125 -126.315 ;
        RECT 14.795 -128.005 15.125 -127.675 ;
        RECT 14.795 -129.365 15.125 -129.035 ;
        RECT 14.795 -130.725 15.125 -130.395 ;
        RECT 14.795 -132.085 15.125 -131.755 ;
        RECT 14.795 -133.445 15.125 -133.115 ;
        RECT 14.795 -134.805 15.125 -134.475 ;
        RECT 14.795 -136.165 15.125 -135.835 ;
        RECT 14.795 -137.525 15.125 -137.195 ;
        RECT 14.795 -138.885 15.125 -138.555 ;
        RECT 14.795 -140.245 15.125 -139.915 ;
        RECT 14.795 -141.605 15.125 -141.275 ;
        RECT 14.795 -142.965 15.125 -142.635 ;
        RECT 14.795 -144.325 15.125 -143.995 ;
        RECT 14.795 -145.685 15.125 -145.355 ;
        RECT 14.795 -147.045 15.125 -146.715 ;
        RECT 14.795 -148.405 15.125 -148.075 ;
        RECT 14.795 -149.765 15.125 -149.435 ;
        RECT 14.795 -151.125 15.125 -150.795 ;
        RECT 14.795 -152.485 15.125 -152.155 ;
        RECT 14.795 -153.845 15.125 -153.515 ;
        RECT 14.795 -155.205 15.125 -154.875 ;
        RECT 14.795 -156.565 15.125 -156.235 ;
        RECT 14.795 -157.925 15.125 -157.595 ;
        RECT 14.795 -159.285 15.125 -158.955 ;
        RECT 14.795 -160.645 15.125 -160.315 ;
        RECT 14.795 -162.005 15.125 -161.675 ;
        RECT 14.795 -163.365 15.125 -163.035 ;
        RECT 14.795 -164.725 15.125 -164.395 ;
        RECT 14.795 -166.085 15.125 -165.755 ;
        RECT 14.795 -167.445 15.125 -167.115 ;
        RECT 14.795 -168.805 15.125 -168.475 ;
        RECT 14.795 -170.165 15.125 -169.835 ;
        RECT 14.795 -171.525 15.125 -171.195 ;
        RECT 14.795 -172.885 15.125 -172.555 ;
        RECT 14.795 -174.245 15.125 -173.915 ;
        RECT 14.795 -175.605 15.125 -175.275 ;
        RECT 14.795 -176.965 15.125 -176.635 ;
        RECT 14.795 -178.325 15.125 -177.995 ;
        RECT 14.795 -180.57 15.125 -179.44 ;
        RECT 14.8 -180.685 15.12 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.51 -94.075 15.84 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.155 241.32 16.485 242.45 ;
        RECT 16.155 239.195 16.485 239.525 ;
        RECT 16.155 237.835 16.485 238.165 ;
        RECT 16.16 237.16 16.48 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.515 241.32 17.845 242.45 ;
        RECT 17.515 239.195 17.845 239.525 ;
        RECT 17.515 237.835 17.845 238.165 ;
        RECT 17.52 237.16 17.84 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.515 -1.525 17.845 -1.195 ;
        RECT 17.515 -2.885 17.845 -2.555 ;
        RECT 17.52 -3.56 17.84 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.875 241.32 19.205 242.45 ;
        RECT 18.875 239.195 19.205 239.525 ;
        RECT 18.875 237.835 19.205 238.165 ;
        RECT 18.88 237.16 19.2 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.875 -1.525 19.205 -1.195 ;
        RECT 18.875 -2.885 19.205 -2.555 ;
        RECT 18.88 -3.56 19.2 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.875 -91.285 19.205 -90.955 ;
        RECT 18.875 -92.645 19.205 -92.315 ;
        RECT 18.875 -94.005 19.205 -93.675 ;
        RECT 18.875 -95.365 19.205 -95.035 ;
        RECT 18.875 -96.725 19.205 -96.395 ;
        RECT 18.875 -98.085 19.205 -97.755 ;
        RECT 18.875 -99.445 19.205 -99.115 ;
        RECT 18.875 -100.805 19.205 -100.475 ;
        RECT 18.875 -102.165 19.205 -101.835 ;
        RECT 18.875 -103.525 19.205 -103.195 ;
        RECT 18.875 -104.885 19.205 -104.555 ;
        RECT 18.875 -106.245 19.205 -105.915 ;
        RECT 18.875 -107.605 19.205 -107.275 ;
        RECT 18.875 -108.965 19.205 -108.635 ;
        RECT 18.875 -110.325 19.205 -109.995 ;
        RECT 18.875 -111.685 19.205 -111.355 ;
        RECT 18.875 -113.045 19.205 -112.715 ;
        RECT 18.875 -114.405 19.205 -114.075 ;
        RECT 18.875 -115.765 19.205 -115.435 ;
        RECT 18.875 -117.125 19.205 -116.795 ;
        RECT 18.875 -118.485 19.205 -118.155 ;
        RECT 18.875 -119.845 19.205 -119.515 ;
        RECT 18.875 -121.205 19.205 -120.875 ;
        RECT 18.875 -122.565 19.205 -122.235 ;
        RECT 18.875 -123.925 19.205 -123.595 ;
        RECT 18.875 -125.285 19.205 -124.955 ;
        RECT 18.875 -126.645 19.205 -126.315 ;
        RECT 18.875 -128.005 19.205 -127.675 ;
        RECT 18.875 -129.365 19.205 -129.035 ;
        RECT 18.875 -130.725 19.205 -130.395 ;
        RECT 18.875 -132.085 19.205 -131.755 ;
        RECT 18.875 -133.445 19.205 -133.115 ;
        RECT 18.875 -134.805 19.205 -134.475 ;
        RECT 18.875 -136.165 19.205 -135.835 ;
        RECT 18.875 -137.525 19.205 -137.195 ;
        RECT 18.875 -138.885 19.205 -138.555 ;
        RECT 18.875 -140.245 19.205 -139.915 ;
        RECT 18.875 -141.605 19.205 -141.275 ;
        RECT 18.875 -142.965 19.205 -142.635 ;
        RECT 18.875 -144.325 19.205 -143.995 ;
        RECT 18.875 -145.685 19.205 -145.355 ;
        RECT 18.875 -147.045 19.205 -146.715 ;
        RECT 18.875 -148.405 19.205 -148.075 ;
        RECT 18.875 -149.765 19.205 -149.435 ;
        RECT 18.875 -151.125 19.205 -150.795 ;
        RECT 18.875 -152.485 19.205 -152.155 ;
        RECT 18.875 -153.845 19.205 -153.515 ;
        RECT 18.875 -155.205 19.205 -154.875 ;
        RECT 18.875 -156.565 19.205 -156.235 ;
        RECT 18.875 -157.925 19.205 -157.595 ;
        RECT 18.875 -159.285 19.205 -158.955 ;
        RECT 18.875 -160.645 19.205 -160.315 ;
        RECT 18.875 -162.005 19.205 -161.675 ;
        RECT 18.875 -163.365 19.205 -163.035 ;
        RECT 18.875 -164.725 19.205 -164.395 ;
        RECT 18.875 -166.085 19.205 -165.755 ;
        RECT 18.875 -167.445 19.205 -167.115 ;
        RECT 18.875 -168.805 19.205 -168.475 ;
        RECT 18.875 -170.165 19.205 -169.835 ;
        RECT 18.875 -171.525 19.205 -171.195 ;
        RECT 18.875 -172.885 19.205 -172.555 ;
        RECT 18.875 -174.245 19.205 -173.915 ;
        RECT 18.875 -175.605 19.205 -175.275 ;
        RECT 18.875 -176.965 19.205 -176.635 ;
        RECT 18.875 -178.325 19.205 -177.995 ;
        RECT 18.875 -180.57 19.205 -179.44 ;
        RECT 18.88 -180.685 19.2 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.235 241.32 20.565 242.45 ;
        RECT 20.235 239.195 20.565 239.525 ;
        RECT 20.235 237.835 20.565 238.165 ;
        RECT 20.24 237.16 20.56 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.235 -1.525 20.565 -1.195 ;
        RECT 20.235 -2.885 20.565 -2.555 ;
        RECT 20.24 -3.56 20.56 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.235 -91.285 20.565 -90.955 ;
        RECT 20.235 -92.645 20.565 -92.315 ;
        RECT 20.235 -94.005 20.565 -93.675 ;
        RECT 20.235 -95.365 20.565 -95.035 ;
        RECT 20.235 -96.725 20.565 -96.395 ;
        RECT 20.235 -98.085 20.565 -97.755 ;
        RECT 20.235 -99.445 20.565 -99.115 ;
        RECT 20.235 -100.805 20.565 -100.475 ;
        RECT 20.235 -102.165 20.565 -101.835 ;
        RECT 20.235 -103.525 20.565 -103.195 ;
        RECT 20.235 -104.885 20.565 -104.555 ;
        RECT 20.235 -106.245 20.565 -105.915 ;
        RECT 20.235 -107.605 20.565 -107.275 ;
        RECT 20.235 -108.965 20.565 -108.635 ;
        RECT 20.235 -110.325 20.565 -109.995 ;
        RECT 20.235 -111.685 20.565 -111.355 ;
        RECT 20.235 -113.045 20.565 -112.715 ;
        RECT 20.235 -114.405 20.565 -114.075 ;
        RECT 20.235 -115.765 20.565 -115.435 ;
        RECT 20.235 -117.125 20.565 -116.795 ;
        RECT 20.235 -118.485 20.565 -118.155 ;
        RECT 20.235 -119.845 20.565 -119.515 ;
        RECT 20.235 -121.205 20.565 -120.875 ;
        RECT 20.235 -122.565 20.565 -122.235 ;
        RECT 20.235 -123.925 20.565 -123.595 ;
        RECT 20.235 -125.285 20.565 -124.955 ;
        RECT 20.235 -126.645 20.565 -126.315 ;
        RECT 20.235 -128.005 20.565 -127.675 ;
        RECT 20.235 -129.365 20.565 -129.035 ;
        RECT 20.235 -130.725 20.565 -130.395 ;
        RECT 20.235 -132.085 20.565 -131.755 ;
        RECT 20.235 -133.445 20.565 -133.115 ;
        RECT 20.235 -134.805 20.565 -134.475 ;
        RECT 20.235 -136.165 20.565 -135.835 ;
        RECT 20.235 -137.525 20.565 -137.195 ;
        RECT 20.235 -138.885 20.565 -138.555 ;
        RECT 20.235 -140.245 20.565 -139.915 ;
        RECT 20.235 -141.605 20.565 -141.275 ;
        RECT 20.235 -142.965 20.565 -142.635 ;
        RECT 20.235 -144.325 20.565 -143.995 ;
        RECT 20.235 -145.685 20.565 -145.355 ;
        RECT 20.235 -147.045 20.565 -146.715 ;
        RECT 20.235 -148.405 20.565 -148.075 ;
        RECT 20.235 -149.765 20.565 -149.435 ;
        RECT 20.235 -151.125 20.565 -150.795 ;
        RECT 20.235 -152.485 20.565 -152.155 ;
        RECT 20.235 -153.845 20.565 -153.515 ;
        RECT 20.235 -155.205 20.565 -154.875 ;
        RECT 20.235 -156.565 20.565 -156.235 ;
        RECT 20.235 -157.925 20.565 -157.595 ;
        RECT 20.235 -159.285 20.565 -158.955 ;
        RECT 20.235 -160.645 20.565 -160.315 ;
        RECT 20.235 -162.005 20.565 -161.675 ;
        RECT 20.235 -163.365 20.565 -163.035 ;
        RECT 20.235 -164.725 20.565 -164.395 ;
        RECT 20.235 -166.085 20.565 -165.755 ;
        RECT 20.235 -167.445 20.565 -167.115 ;
        RECT 20.235 -168.805 20.565 -168.475 ;
        RECT 20.235 -170.165 20.565 -169.835 ;
        RECT 20.235 -171.525 20.565 -171.195 ;
        RECT 20.235 -172.885 20.565 -172.555 ;
        RECT 20.235 -174.245 20.565 -173.915 ;
        RECT 20.235 -175.605 20.565 -175.275 ;
        RECT 20.235 -176.965 20.565 -176.635 ;
        RECT 20.235 -178.325 20.565 -177.995 ;
        RECT 20.235 -180.57 20.565 -179.44 ;
        RECT 20.24 -180.685 20.56 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.595 241.32 21.925 242.45 ;
        RECT 21.595 239.195 21.925 239.525 ;
        RECT 21.595 237.835 21.925 238.165 ;
        RECT 21.6 237.16 21.92 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.595 -95.365 21.925 -95.035 ;
        RECT 21.595 -96.725 21.925 -96.395 ;
        RECT 21.595 -98.085 21.925 -97.755 ;
        RECT 21.595 -99.445 21.925 -99.115 ;
        RECT 21.595 -100.805 21.925 -100.475 ;
        RECT 21.595 -102.165 21.925 -101.835 ;
        RECT 21.595 -103.525 21.925 -103.195 ;
        RECT 21.595 -104.885 21.925 -104.555 ;
        RECT 21.595 -106.245 21.925 -105.915 ;
        RECT 21.595 -107.605 21.925 -107.275 ;
        RECT 21.595 -108.965 21.925 -108.635 ;
        RECT 21.595 -110.325 21.925 -109.995 ;
        RECT 21.595 -111.685 21.925 -111.355 ;
        RECT 21.595 -113.045 21.925 -112.715 ;
        RECT 21.595 -114.405 21.925 -114.075 ;
        RECT 21.595 -115.765 21.925 -115.435 ;
        RECT 21.595 -117.125 21.925 -116.795 ;
        RECT 21.595 -118.485 21.925 -118.155 ;
        RECT 21.595 -119.845 21.925 -119.515 ;
        RECT 21.595 -121.205 21.925 -120.875 ;
        RECT 21.595 -122.565 21.925 -122.235 ;
        RECT 21.595 -123.925 21.925 -123.595 ;
        RECT 21.595 -125.285 21.925 -124.955 ;
        RECT 21.595 -126.645 21.925 -126.315 ;
        RECT 21.595 -128.005 21.925 -127.675 ;
        RECT 21.595 -129.365 21.925 -129.035 ;
        RECT 21.595 -130.725 21.925 -130.395 ;
        RECT 21.595 -132.085 21.925 -131.755 ;
        RECT 21.595 -133.445 21.925 -133.115 ;
        RECT 21.595 -134.805 21.925 -134.475 ;
        RECT 21.595 -136.165 21.925 -135.835 ;
        RECT 21.595 -137.525 21.925 -137.195 ;
        RECT 21.595 -138.885 21.925 -138.555 ;
        RECT 21.595 -140.245 21.925 -139.915 ;
        RECT 21.595 -141.605 21.925 -141.275 ;
        RECT 21.595 -142.965 21.925 -142.635 ;
        RECT 21.595 -144.325 21.925 -143.995 ;
        RECT 21.595 -145.685 21.925 -145.355 ;
        RECT 21.595 -147.045 21.925 -146.715 ;
        RECT 21.595 -148.405 21.925 -148.075 ;
        RECT 21.595 -149.765 21.925 -149.435 ;
        RECT 21.595 -151.125 21.925 -150.795 ;
        RECT 21.595 -152.485 21.925 -152.155 ;
        RECT 21.595 -153.845 21.925 -153.515 ;
        RECT 21.595 -155.205 21.925 -154.875 ;
        RECT 21.595 -156.565 21.925 -156.235 ;
        RECT 21.595 -157.925 21.925 -157.595 ;
        RECT 21.595 -159.285 21.925 -158.955 ;
        RECT 21.595 -160.645 21.925 -160.315 ;
        RECT 21.595 -162.005 21.925 -161.675 ;
        RECT 21.595 -163.365 21.925 -163.035 ;
        RECT 21.595 -164.725 21.925 -164.395 ;
        RECT 21.595 -166.085 21.925 -165.755 ;
        RECT 21.595 -167.445 21.925 -167.115 ;
        RECT 21.595 -168.805 21.925 -168.475 ;
        RECT 21.595 -170.165 21.925 -169.835 ;
        RECT 21.595 -171.525 21.925 -171.195 ;
        RECT 21.595 -172.885 21.925 -172.555 ;
        RECT 21.595 -174.245 21.925 -173.915 ;
        RECT 21.595 -175.605 21.925 -175.275 ;
        RECT 21.595 -176.965 21.925 -176.635 ;
        RECT 21.595 -178.325 21.925 -177.995 ;
        RECT 21.595 -180.57 21.925 -179.44 ;
        RECT 21.6 -180.685 21.92 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.61 -94.075 21.94 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.955 241.32 23.285 242.45 ;
        RECT 22.955 239.195 23.285 239.525 ;
        RECT 22.955 237.835 23.285 238.165 ;
        RECT 22.96 237.16 23.28 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.955 -1.525 23.285 -1.195 ;
        RECT 22.955 -2.885 23.285 -2.555 ;
        RECT 22.96 -3.56 23.28 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.315 241.32 24.645 242.45 ;
        RECT 24.315 239.195 24.645 239.525 ;
        RECT 24.315 237.835 24.645 238.165 ;
        RECT 24.32 237.16 24.64 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.315 -1.525 24.645 -1.195 ;
        RECT 24.315 -2.885 24.645 -2.555 ;
        RECT 24.32 -3.56 24.64 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.675 241.32 26.005 242.45 ;
        RECT 25.675 239.195 26.005 239.525 ;
        RECT 25.675 237.835 26.005 238.165 ;
        RECT 25.68 237.16 26 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.675 -1.525 26.005 -1.195 ;
        RECT 25.675 -2.885 26.005 -2.555 ;
        RECT 25.68 -3.56 26 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.675 -91.285 26.005 -90.955 ;
        RECT 25.675 -92.645 26.005 -92.315 ;
        RECT 25.675 -94.005 26.005 -93.675 ;
        RECT 25.675 -95.365 26.005 -95.035 ;
        RECT 25.675 -96.725 26.005 -96.395 ;
        RECT 25.675 -98.085 26.005 -97.755 ;
        RECT 25.675 -99.445 26.005 -99.115 ;
        RECT 25.675 -100.805 26.005 -100.475 ;
        RECT 25.675 -102.165 26.005 -101.835 ;
        RECT 25.675 -103.525 26.005 -103.195 ;
        RECT 25.675 -104.885 26.005 -104.555 ;
        RECT 25.675 -106.245 26.005 -105.915 ;
        RECT 25.675 -107.605 26.005 -107.275 ;
        RECT 25.675 -108.965 26.005 -108.635 ;
        RECT 25.675 -110.325 26.005 -109.995 ;
        RECT 25.675 -111.685 26.005 -111.355 ;
        RECT 25.675 -113.045 26.005 -112.715 ;
        RECT 25.675 -114.405 26.005 -114.075 ;
        RECT 25.675 -115.765 26.005 -115.435 ;
        RECT 25.675 -117.125 26.005 -116.795 ;
        RECT 25.675 -118.485 26.005 -118.155 ;
        RECT 25.675 -119.845 26.005 -119.515 ;
        RECT 25.675 -121.205 26.005 -120.875 ;
        RECT 25.675 -122.565 26.005 -122.235 ;
        RECT 25.675 -123.925 26.005 -123.595 ;
        RECT 25.675 -125.285 26.005 -124.955 ;
        RECT 25.675 -126.645 26.005 -126.315 ;
        RECT 25.675 -128.005 26.005 -127.675 ;
        RECT 25.675 -129.365 26.005 -129.035 ;
        RECT 25.675 -130.725 26.005 -130.395 ;
        RECT 25.675 -132.085 26.005 -131.755 ;
        RECT 25.675 -133.445 26.005 -133.115 ;
        RECT 25.675 -134.805 26.005 -134.475 ;
        RECT 25.675 -136.165 26.005 -135.835 ;
        RECT 25.675 -137.525 26.005 -137.195 ;
        RECT 25.675 -138.885 26.005 -138.555 ;
        RECT 25.675 -140.245 26.005 -139.915 ;
        RECT 25.675 -141.605 26.005 -141.275 ;
        RECT 25.675 -142.965 26.005 -142.635 ;
        RECT 25.675 -144.325 26.005 -143.995 ;
        RECT 25.675 -145.685 26.005 -145.355 ;
        RECT 25.675 -147.045 26.005 -146.715 ;
        RECT 25.675 -148.405 26.005 -148.075 ;
        RECT 25.675 -149.765 26.005 -149.435 ;
        RECT 25.675 -151.125 26.005 -150.795 ;
        RECT 25.675 -152.485 26.005 -152.155 ;
        RECT 25.675 -153.845 26.005 -153.515 ;
        RECT 25.675 -155.205 26.005 -154.875 ;
        RECT 25.675 -156.565 26.005 -156.235 ;
        RECT 25.675 -157.925 26.005 -157.595 ;
        RECT 25.675 -159.285 26.005 -158.955 ;
        RECT 25.675 -160.645 26.005 -160.315 ;
        RECT 25.675 -162.005 26.005 -161.675 ;
        RECT 25.675 -163.365 26.005 -163.035 ;
        RECT 25.675 -164.725 26.005 -164.395 ;
        RECT 25.675 -166.085 26.005 -165.755 ;
        RECT 25.675 -167.445 26.005 -167.115 ;
        RECT 25.675 -168.805 26.005 -168.475 ;
        RECT 25.675 -170.165 26.005 -169.835 ;
        RECT 25.675 -171.525 26.005 -171.195 ;
        RECT 25.675 -172.885 26.005 -172.555 ;
        RECT 25.675 -174.245 26.005 -173.915 ;
        RECT 25.675 -175.605 26.005 -175.275 ;
        RECT 25.675 -176.965 26.005 -176.635 ;
        RECT 25.675 -178.325 26.005 -177.995 ;
        RECT 25.675 -180.57 26.005 -179.44 ;
        RECT 25.68 -180.685 26 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.035 241.32 27.365 242.45 ;
        RECT 27.035 239.195 27.365 239.525 ;
        RECT 27.035 237.835 27.365 238.165 ;
        RECT 27.04 237.16 27.36 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.035 -95.365 27.365 -95.035 ;
        RECT 27.035 -96.725 27.365 -96.395 ;
        RECT 27.035 -98.085 27.365 -97.755 ;
        RECT 27.035 -99.445 27.365 -99.115 ;
        RECT 27.035 -100.805 27.365 -100.475 ;
        RECT 27.035 -102.165 27.365 -101.835 ;
        RECT 27.035 -103.525 27.365 -103.195 ;
        RECT 27.035 -104.885 27.365 -104.555 ;
        RECT 27.035 -106.245 27.365 -105.915 ;
        RECT 27.035 -107.605 27.365 -107.275 ;
        RECT 27.035 -108.965 27.365 -108.635 ;
        RECT 27.035 -110.325 27.365 -109.995 ;
        RECT 27.035 -111.685 27.365 -111.355 ;
        RECT 27.035 -113.045 27.365 -112.715 ;
        RECT 27.035 -114.405 27.365 -114.075 ;
        RECT 27.035 -115.765 27.365 -115.435 ;
        RECT 27.035 -117.125 27.365 -116.795 ;
        RECT 27.035 -118.485 27.365 -118.155 ;
        RECT 27.035 -119.845 27.365 -119.515 ;
        RECT 27.035 -121.205 27.365 -120.875 ;
        RECT 27.035 -122.565 27.365 -122.235 ;
        RECT 27.035 -123.925 27.365 -123.595 ;
        RECT 27.035 -125.285 27.365 -124.955 ;
        RECT 27.035 -126.645 27.365 -126.315 ;
        RECT 27.035 -128.005 27.365 -127.675 ;
        RECT 27.035 -129.365 27.365 -129.035 ;
        RECT 27.035 -130.725 27.365 -130.395 ;
        RECT 27.035 -132.085 27.365 -131.755 ;
        RECT 27.035 -133.445 27.365 -133.115 ;
        RECT 27.035 -134.805 27.365 -134.475 ;
        RECT 27.035 -136.165 27.365 -135.835 ;
        RECT 27.035 -137.525 27.365 -137.195 ;
        RECT 27.035 -138.885 27.365 -138.555 ;
        RECT 27.035 -140.245 27.365 -139.915 ;
        RECT 27.035 -141.605 27.365 -141.275 ;
        RECT 27.035 -142.965 27.365 -142.635 ;
        RECT 27.035 -144.325 27.365 -143.995 ;
        RECT 27.035 -145.685 27.365 -145.355 ;
        RECT 27.035 -147.045 27.365 -146.715 ;
        RECT 27.035 -148.405 27.365 -148.075 ;
        RECT 27.035 -149.765 27.365 -149.435 ;
        RECT 27.035 -151.125 27.365 -150.795 ;
        RECT 27.035 -152.485 27.365 -152.155 ;
        RECT 27.035 -153.845 27.365 -153.515 ;
        RECT 27.035 -155.205 27.365 -154.875 ;
        RECT 27.035 -156.565 27.365 -156.235 ;
        RECT 27.035 -157.925 27.365 -157.595 ;
        RECT 27.035 -159.285 27.365 -158.955 ;
        RECT 27.035 -160.645 27.365 -160.315 ;
        RECT 27.035 -162.005 27.365 -161.675 ;
        RECT 27.035 -163.365 27.365 -163.035 ;
        RECT 27.035 -164.725 27.365 -164.395 ;
        RECT 27.035 -166.085 27.365 -165.755 ;
        RECT 27.035 -167.445 27.365 -167.115 ;
        RECT 27.035 -168.805 27.365 -168.475 ;
        RECT 27.035 -170.165 27.365 -169.835 ;
        RECT 27.035 -171.525 27.365 -171.195 ;
        RECT 27.035 -172.885 27.365 -172.555 ;
        RECT 27.035 -174.245 27.365 -173.915 ;
        RECT 27.035 -175.605 27.365 -175.275 ;
        RECT 27.035 -176.965 27.365 -176.635 ;
        RECT 27.035 -178.325 27.365 -177.995 ;
        RECT 27.035 -180.57 27.365 -179.44 ;
        RECT 27.04 -180.685 27.36 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.71 -94.075 28.04 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.395 241.32 28.725 242.45 ;
        RECT 28.395 239.195 28.725 239.525 ;
        RECT 28.395 237.835 28.725 238.165 ;
        RECT 28.4 237.16 28.72 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.395 -1.525 28.725 -1.195 ;
        RECT 28.395 -2.885 28.725 -2.555 ;
        RECT 28.4 -3.56 28.72 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.755 241.32 30.085 242.45 ;
        RECT 29.755 239.195 30.085 239.525 ;
        RECT 29.755 237.835 30.085 238.165 ;
        RECT 29.76 237.16 30.08 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.755 -1.525 30.085 -1.195 ;
        RECT 29.755 -2.885 30.085 -2.555 ;
        RECT 29.76 -3.56 30.08 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.115 241.32 31.445 242.45 ;
        RECT 31.115 239.195 31.445 239.525 ;
        RECT 31.115 237.835 31.445 238.165 ;
        RECT 31.12 237.16 31.44 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.115 -1.525 31.445 -1.195 ;
        RECT 31.115 -2.885 31.445 -2.555 ;
        RECT 31.12 -3.56 31.44 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.12 -180.685 31.44 -90.955 ;
        RECT 31.115 -91.285 31.445 -90.955 ;
        RECT 31.115 -92.645 31.445 -92.315 ;
        RECT 31.115 -94.005 31.445 -93.675 ;
        RECT 31.115 -95.365 31.445 -95.035 ;
        RECT 31.115 -96.725 31.445 -96.395 ;
        RECT 31.115 -98.085 31.445 -97.755 ;
        RECT 31.115 -99.445 31.445 -99.115 ;
        RECT 31.115 -100.805 31.445 -100.475 ;
        RECT 31.115 -102.165 31.445 -101.835 ;
        RECT 31.115 -103.525 31.445 -103.195 ;
        RECT 31.115 -104.885 31.445 -104.555 ;
        RECT 31.115 -106.245 31.445 -105.915 ;
        RECT 31.115 -107.605 31.445 -107.275 ;
        RECT 31.115 -108.965 31.445 -108.635 ;
        RECT 31.115 -110.325 31.445 -109.995 ;
        RECT 31.115 -111.685 31.445 -111.355 ;
        RECT 31.115 -113.045 31.445 -112.715 ;
        RECT 31.115 -114.405 31.445 -114.075 ;
        RECT 31.115 -115.765 31.445 -115.435 ;
        RECT 31.115 -117.125 31.445 -116.795 ;
        RECT 31.115 -118.485 31.445 -118.155 ;
        RECT 31.115 -119.845 31.445 -119.515 ;
        RECT 31.115 -121.205 31.445 -120.875 ;
        RECT 31.115 -122.565 31.445 -122.235 ;
        RECT 31.115 -123.925 31.445 -123.595 ;
        RECT 31.115 -125.285 31.445 -124.955 ;
        RECT 31.115 -126.645 31.445 -126.315 ;
        RECT 31.115 -128.005 31.445 -127.675 ;
        RECT 31.115 -129.365 31.445 -129.035 ;
        RECT 31.115 -130.725 31.445 -130.395 ;
        RECT 31.115 -132.085 31.445 -131.755 ;
        RECT 31.115 -133.445 31.445 -133.115 ;
        RECT 31.115 -134.805 31.445 -134.475 ;
        RECT 31.115 -136.165 31.445 -135.835 ;
        RECT 31.115 -137.525 31.445 -137.195 ;
        RECT 31.115 -138.885 31.445 -138.555 ;
        RECT 31.115 -140.245 31.445 -139.915 ;
        RECT 31.115 -141.605 31.445 -141.275 ;
        RECT 31.115 -142.965 31.445 -142.635 ;
        RECT 31.115 -144.325 31.445 -143.995 ;
        RECT 31.115 -145.685 31.445 -145.355 ;
        RECT 31.115 -147.045 31.445 -146.715 ;
        RECT 31.115 -148.405 31.445 -148.075 ;
        RECT 31.115 -149.765 31.445 -149.435 ;
        RECT 31.115 -151.125 31.445 -150.795 ;
        RECT 31.115 -152.485 31.445 -152.155 ;
        RECT 31.115 -153.845 31.445 -153.515 ;
        RECT 31.115 -155.205 31.445 -154.875 ;
        RECT 31.115 -156.565 31.445 -156.235 ;
        RECT 31.115 -157.925 31.445 -157.595 ;
        RECT 31.115 -159.285 31.445 -158.955 ;
        RECT 31.115 -160.645 31.445 -160.315 ;
        RECT 31.115 -162.005 31.445 -161.675 ;
        RECT 31.115 -163.365 31.445 -163.035 ;
        RECT 31.115 -164.725 31.445 -164.395 ;
        RECT 31.115 -166.085 31.445 -165.755 ;
        RECT 31.115 -167.445 31.445 -167.115 ;
        RECT 31.115 -168.805 31.445 -168.475 ;
        RECT 31.115 -170.165 31.445 -169.835 ;
        RECT 31.115 -171.525 31.445 -171.195 ;
        RECT 31.115 -172.885 31.445 -172.555 ;
        RECT 31.115 -174.245 31.445 -173.915 ;
        RECT 31.115 -175.605 31.445 -175.275 ;
        RECT 31.115 -176.965 31.445 -176.635 ;
        RECT 31.115 -178.325 31.445 -177.995 ;
        RECT 31.115 -180.57 31.445 -179.44 ;
    END
    PORT
      LAYER met3 ;
        RECT -4.245 241.32 -3.915 242.45 ;
        RECT -4.245 239.195 -3.915 239.525 ;
        RECT -4.245 237.835 -3.915 238.165 ;
        RECT -4.245 235.975 -3.915 236.305 ;
        RECT -4.245 233.925 -3.915 234.255 ;
        RECT -4.245 231.995 -3.915 232.325 ;
        RECT -4.245 230.155 -3.915 230.485 ;
        RECT -4.245 228.665 -3.915 228.995 ;
        RECT -4.245 226.995 -3.915 227.325 ;
        RECT -4.245 225.505 -3.915 225.835 ;
        RECT -4.245 223.835 -3.915 224.165 ;
        RECT -4.245 222.345 -3.915 222.675 ;
        RECT -4.245 220.675 -3.915 221.005 ;
        RECT -4.245 219.185 -3.915 219.515 ;
        RECT -4.245 217.775 -3.915 218.105 ;
        RECT -4.245 215.935 -3.915 216.265 ;
        RECT -4.245 214.445 -3.915 214.775 ;
        RECT -4.245 212.775 -3.915 213.105 ;
        RECT -4.245 211.285 -3.915 211.615 ;
        RECT -4.245 209.615 -3.915 209.945 ;
        RECT -4.245 208.125 -3.915 208.455 ;
        RECT -4.245 206.455 -3.915 206.785 ;
        RECT -4.245 204.965 -3.915 205.295 ;
        RECT -4.245 203.555 -3.915 203.885 ;
        RECT -4.245 201.715 -3.915 202.045 ;
        RECT -4.245 200.225 -3.915 200.555 ;
        RECT -4.245 198.555 -3.915 198.885 ;
        RECT -4.245 197.065 -3.915 197.395 ;
        RECT -4.245 195.395 -3.915 195.725 ;
        RECT -4.245 193.905 -3.915 194.235 ;
        RECT -4.245 192.235 -3.915 192.565 ;
        RECT -4.245 190.745 -3.915 191.075 ;
        RECT -4.245 189.335 -3.915 189.665 ;
        RECT -4.245 187.495 -3.915 187.825 ;
        RECT -4.245 186.005 -3.915 186.335 ;
        RECT -4.245 184.335 -3.915 184.665 ;
        RECT -4.245 182.845 -3.915 183.175 ;
        RECT -4.245 181.175 -3.915 181.505 ;
        RECT -4.245 179.685 -3.915 180.015 ;
        RECT -4.245 178.015 -3.915 178.345 ;
        RECT -4.245 176.525 -3.915 176.855 ;
        RECT -4.245 175.115 -3.915 175.445 ;
        RECT -4.245 173.275 -3.915 173.605 ;
        RECT -4.245 171.785 -3.915 172.115 ;
        RECT -4.245 170.115 -3.915 170.445 ;
        RECT -4.245 168.625 -3.915 168.955 ;
        RECT -4.245 166.955 -3.915 167.285 ;
        RECT -4.245 165.465 -3.915 165.795 ;
        RECT -4.245 163.795 -3.915 164.125 ;
        RECT -4.245 162.305 -3.915 162.635 ;
        RECT -4.245 160.895 -3.915 161.225 ;
        RECT -4.245 159.055 -3.915 159.385 ;
        RECT -4.245 157.565 -3.915 157.895 ;
        RECT -4.245 155.895 -3.915 156.225 ;
        RECT -4.245 154.405 -3.915 154.735 ;
        RECT -4.245 152.735 -3.915 153.065 ;
        RECT -4.245 151.245 -3.915 151.575 ;
        RECT -4.245 149.575 -3.915 149.905 ;
        RECT -4.245 148.085 -3.915 148.415 ;
        RECT -4.245 146.675 -3.915 147.005 ;
        RECT -4.245 144.835 -3.915 145.165 ;
        RECT -4.245 143.345 -3.915 143.675 ;
        RECT -4.245 141.675 -3.915 142.005 ;
        RECT -4.245 140.185 -3.915 140.515 ;
        RECT -4.245 138.515 -3.915 138.845 ;
        RECT -4.245 137.025 -3.915 137.355 ;
        RECT -4.245 135.355 -3.915 135.685 ;
        RECT -4.245 133.865 -3.915 134.195 ;
        RECT -4.245 132.455 -3.915 132.785 ;
        RECT -4.245 130.615 -3.915 130.945 ;
        RECT -4.245 129.125 -3.915 129.455 ;
        RECT -4.245 127.455 -3.915 127.785 ;
        RECT -4.245 125.965 -3.915 126.295 ;
        RECT -4.245 124.295 -3.915 124.625 ;
        RECT -4.245 122.805 -3.915 123.135 ;
        RECT -4.245 121.135 -3.915 121.465 ;
        RECT -4.245 119.645 -3.915 119.975 ;
        RECT -4.245 118.235 -3.915 118.565 ;
        RECT -4.245 116.395 -3.915 116.725 ;
        RECT -4.245 114.905 -3.915 115.235 ;
        RECT -4.245 113.235 -3.915 113.565 ;
        RECT -4.245 111.745 -3.915 112.075 ;
        RECT -4.245 110.075 -3.915 110.405 ;
        RECT -4.245 108.585 -3.915 108.915 ;
        RECT -4.245 106.915 -3.915 107.245 ;
        RECT -4.245 105.425 -3.915 105.755 ;
        RECT -4.245 104.015 -3.915 104.345 ;
        RECT -4.245 102.175 -3.915 102.505 ;
        RECT -4.245 100.685 -3.915 101.015 ;
        RECT -4.245 99.015 -3.915 99.345 ;
        RECT -4.245 97.525 -3.915 97.855 ;
        RECT -4.245 95.855 -3.915 96.185 ;
        RECT -4.245 94.365 -3.915 94.695 ;
        RECT -4.245 92.695 -3.915 93.025 ;
        RECT -4.245 91.205 -3.915 91.535 ;
        RECT -4.245 89.795 -3.915 90.125 ;
        RECT -4.245 87.955 -3.915 88.285 ;
        RECT -4.245 86.465 -3.915 86.795 ;
        RECT -4.245 84.795 -3.915 85.125 ;
        RECT -4.245 83.305 -3.915 83.635 ;
        RECT -4.245 81.635 -3.915 81.965 ;
        RECT -4.245 80.145 -3.915 80.475 ;
        RECT -4.245 78.475 -3.915 78.805 ;
        RECT -4.245 76.985 -3.915 77.315 ;
        RECT -4.245 75.575 -3.915 75.905 ;
        RECT -4.245 73.735 -3.915 74.065 ;
        RECT -4.245 72.245 -3.915 72.575 ;
        RECT -4.245 70.575 -3.915 70.905 ;
        RECT -4.245 69.085 -3.915 69.415 ;
        RECT -4.245 67.415 -3.915 67.745 ;
        RECT -4.245 65.925 -3.915 66.255 ;
        RECT -4.245 64.255 -3.915 64.585 ;
        RECT -4.245 62.765 -3.915 63.095 ;
        RECT -4.245 61.355 -3.915 61.685 ;
        RECT -4.245 59.515 -3.915 59.845 ;
        RECT -4.245 58.025 -3.915 58.355 ;
        RECT -4.245 56.355 -3.915 56.685 ;
        RECT -4.245 54.865 -3.915 55.195 ;
        RECT -4.245 53.195 -3.915 53.525 ;
        RECT -4.245 51.705 -3.915 52.035 ;
        RECT -4.245 50.035 -3.915 50.365 ;
        RECT -4.245 48.545 -3.915 48.875 ;
        RECT -4.245 47.135 -3.915 47.465 ;
        RECT -4.245 45.295 -3.915 45.625 ;
        RECT -4.245 43.805 -3.915 44.135 ;
        RECT -4.245 42.135 -3.915 42.465 ;
        RECT -4.245 40.645 -3.915 40.975 ;
        RECT -4.245 38.975 -3.915 39.305 ;
        RECT -4.245 37.485 -3.915 37.815 ;
        RECT -4.245 35.815 -3.915 36.145 ;
        RECT -4.245 34.325 -3.915 34.655 ;
        RECT -4.245 32.915 -3.915 33.245 ;
        RECT -4.245 31.075 -3.915 31.405 ;
        RECT -4.245 29.585 -3.915 29.915 ;
        RECT -4.245 27.915 -3.915 28.245 ;
        RECT -4.245 26.425 -3.915 26.755 ;
        RECT -4.245 24.755 -3.915 25.085 ;
        RECT -4.245 23.265 -3.915 23.595 ;
        RECT -4.245 21.595 -3.915 21.925 ;
        RECT -4.245 20.105 -3.915 20.435 ;
        RECT -4.245 18.695 -3.915 19.025 ;
        RECT -4.245 16.855 -3.915 17.185 ;
        RECT -4.245 15.365 -3.915 15.695 ;
        RECT -4.245 13.695 -3.915 14.025 ;
        RECT -4.245 12.205 -3.915 12.535 ;
        RECT -4.245 10.535 -3.915 10.865 ;
        RECT -4.245 9.045 -3.915 9.375 ;
        RECT -4.245 7.375 -3.915 7.705 ;
        RECT -4.245 5.885 -3.915 6.215 ;
        RECT -4.245 4.475 -3.915 4.805 ;
        RECT -4.245 2.115 -3.915 2.445 ;
        RECT -4.245 0.06 -3.915 0.39 ;
        RECT -4.245 -1.525 -3.915 -1.195 ;
        RECT -4.245 -2.885 -3.915 -2.555 ;
        RECT -4.245 -4.245 -3.915 -3.915 ;
        RECT -4.245 -5.605 -3.915 -5.275 ;
        RECT -4.245 -6.965 -3.915 -6.635 ;
        RECT -4.245 -8.325 -3.915 -7.995 ;
        RECT -4.245 -9.685 -3.915 -9.355 ;
        RECT -4.245 -12.405 -3.915 -12.075 ;
        RECT -4.245 -13.765 -3.915 -13.435 ;
        RECT -4.245 -15.125 -3.915 -14.795 ;
        RECT -4.245 -16.485 -3.915 -16.155 ;
        RECT -4.245 -17.845 -3.915 -17.515 ;
        RECT -4.245 -21.925 -3.915 -21.595 ;
        RECT -4.245 -23.285 -3.915 -22.955 ;
        RECT -4.245 -24.645 -3.915 -24.315 ;
        RECT -4.245 -26.005 -3.915 -25.675 ;
        RECT -4.245 -27.365 -3.915 -27.035 ;
        RECT -4.245 -28.725 -3.915 -28.395 ;
        RECT -4.245 -30.085 -3.915 -29.755 ;
        RECT -4.245 -31.445 -3.915 -31.115 ;
        RECT -4.245 -32.805 -3.915 -32.475 ;
        RECT -4.245 -34.165 -3.915 -33.835 ;
        RECT -4.245 -36.885 -3.915 -36.555 ;
        RECT -4.245 -38.245 -3.915 -37.915 ;
        RECT -4.245 -40.965 -3.915 -40.635 ;
        RECT -4.245 -42.325 -3.915 -41.995 ;
        RECT -4.245 -43.685 -3.915 -43.355 ;
        RECT -4.245 -45.045 -3.915 -44.715 ;
        RECT -4.245 -46.405 -3.915 -46.075 ;
        RECT -4.245 -47.765 -3.915 -47.435 ;
        RECT -4.245 -49.125 -3.915 -48.795 ;
        RECT -4.245 -51.845 -3.915 -51.515 ;
        RECT -4.245 -53.205 -3.915 -52.875 ;
        RECT -4.245 -54.565 -3.915 -54.235 ;
        RECT -4.245 -55.925 -3.915 -55.595 ;
        RECT -4.245 -57.285 -3.915 -56.955 ;
        RECT -4.245 -58.645 -3.915 -58.315 ;
        RECT -4.245 -60.005 -3.915 -59.675 ;
        RECT -4.245 -61.365 -3.915 -61.035 ;
        RECT -4.245 -62.725 -3.915 -62.395 ;
        RECT -4.245 -64.085 -3.915 -63.755 ;
        RECT -4.245 -65.445 -3.915 -65.115 ;
        RECT -4.245 -66.805 -3.915 -66.475 ;
        RECT -4.245 -68.165 -3.915 -67.835 ;
        RECT -4.245 -69.525 -3.915 -69.195 ;
        RECT -4.245 -70.885 -3.915 -70.555 ;
        RECT -4.245 -72.245 -3.915 -71.915 ;
        RECT -4.245 -73.605 -3.915 -73.275 ;
        RECT -4.245 -74.965 -3.915 -74.635 ;
        RECT -4.245 -76.325 -3.915 -75.995 ;
        RECT -4.245 -77.685 -3.915 -77.355 ;
        RECT -4.245 -79.045 -3.915 -78.715 ;
        RECT -4.245 -80.405 -3.915 -80.075 ;
        RECT -4.245 -81.765 -3.915 -81.435 ;
        RECT -4.245 -83.125 -3.915 -82.795 ;
        RECT -4.245 -84.485 -3.915 -84.155 ;
        RECT -4.245 -85.845 -3.915 -85.515 ;
        RECT -4.245 -87.205 -3.915 -86.875 ;
        RECT -4.245 -88.565 -3.915 -88.235 ;
        RECT -4.245 -89.925 -3.915 -89.595 ;
        RECT -4.245 -91.285 -3.915 -90.955 ;
        RECT -4.245 -92.645 -3.915 -92.315 ;
        RECT -4.245 -94.005 -3.915 -93.675 ;
        RECT -4.245 -95.365 -3.915 -95.035 ;
        RECT -4.245 -96.725 -3.915 -96.395 ;
        RECT -4.245 -98.085 -3.915 -97.755 ;
        RECT -4.245 -99.445 -3.915 -99.115 ;
        RECT -4.245 -100.805 -3.915 -100.475 ;
        RECT -4.245 -102.165 -3.915 -101.835 ;
        RECT -4.245 -103.525 -3.915 -103.195 ;
        RECT -4.245 -104.885 -3.915 -104.555 ;
        RECT -4.245 -106.245 -3.915 -105.915 ;
        RECT -4.245 -107.605 -3.915 -107.275 ;
        RECT -4.245 -108.965 -3.915 -108.635 ;
        RECT -4.245 -110.325 -3.915 -109.995 ;
        RECT -4.245 -111.685 -3.915 -111.355 ;
        RECT -4.245 -113.045 -3.915 -112.715 ;
        RECT -4.245 -114.405 -3.915 -114.075 ;
        RECT -4.245 -115.765 -3.915 -115.435 ;
        RECT -4.245 -117.125 -3.915 -116.795 ;
        RECT -4.245 -119.845 -3.915 -119.515 ;
        RECT -4.245 -121.205 -3.915 -120.875 ;
        RECT -4.245 -122.565 -3.915 -122.235 ;
        RECT -4.245 -123.925 -3.915 -123.595 ;
        RECT -4.245 -125.285 -3.915 -124.955 ;
        RECT -4.245 -126.645 -3.915 -126.315 ;
        RECT -4.245 -128.005 -3.915 -127.675 ;
        RECT -4.245 -129.365 -3.915 -129.035 ;
        RECT -4.245 -130.725 -3.915 -130.395 ;
        RECT -4.245 -132.085 -3.915 -131.755 ;
        RECT -4.245 -133.445 -3.915 -133.115 ;
        RECT -4.245 -134.805 -3.915 -134.475 ;
        RECT -4.245 -136.165 -3.915 -135.835 ;
        RECT -4.245 -137.525 -3.915 -137.195 ;
        RECT -4.245 -138.885 -3.915 -138.555 ;
        RECT -4.245 -140.245 -3.915 -139.915 ;
        RECT -4.245 -141.605 -3.915 -141.275 ;
        RECT -4.245 -142.965 -3.915 -142.635 ;
        RECT -4.245 -144.325 -3.915 -143.995 ;
        RECT -4.245 -145.685 -3.915 -145.355 ;
        RECT -4.245 -147.045 -3.915 -146.715 ;
        RECT -4.245 -148.405 -3.915 -148.075 ;
        RECT -4.245 -149.765 -3.915 -149.435 ;
        RECT -4.245 -151.125 -3.915 -150.795 ;
        RECT -4.245 -152.485 -3.915 -152.155 ;
        RECT -4.245 -153.845 -3.915 -153.515 ;
        RECT -4.245 -155.205 -3.915 -154.875 ;
        RECT -4.245 -156.565 -3.915 -156.235 ;
        RECT -4.245 -157.925 -3.915 -157.595 ;
        RECT -4.245 -159.285 -3.915 -158.955 ;
        RECT -4.245 -160.645 -3.915 -160.315 ;
        RECT -4.245 -162.005 -3.915 -161.675 ;
        RECT -4.245 -163.365 -3.915 -163.035 ;
        RECT -4.245 -164.725 -3.915 -164.395 ;
        RECT -4.245 -166.085 -3.915 -165.755 ;
        RECT -4.245 -167.445 -3.915 -167.115 ;
        RECT -4.245 -168.805 -3.915 -168.475 ;
        RECT -4.245 -170.165 -3.915 -169.835 ;
        RECT -4.245 -171.525 -3.915 -171.195 ;
        RECT -4.245 -172.885 -3.915 -172.555 ;
        RECT -4.245 -174.245 -3.915 -173.915 ;
        RECT -4.245 -175.605 -3.915 -175.275 ;
        RECT -4.245 -176.965 -3.915 -176.635 ;
        RECT -4.245 -178.325 -3.915 -177.995 ;
        RECT -4.245 -180.57 -3.915 -179.44 ;
        RECT -4.24 -180.685 -3.92 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -2.885 241.32 -2.555 242.45 ;
        RECT -2.885 239.195 -2.555 239.525 ;
        RECT -2.885 237.835 -2.555 238.165 ;
        RECT -2.885 235.975 -2.555 236.305 ;
        RECT -2.885 233.925 -2.555 234.255 ;
        RECT -2.885 231.995 -2.555 232.325 ;
        RECT -2.885 230.155 -2.555 230.485 ;
        RECT -2.885 228.665 -2.555 228.995 ;
        RECT -2.885 226.995 -2.555 227.325 ;
        RECT -2.885 225.505 -2.555 225.835 ;
        RECT -2.885 223.835 -2.555 224.165 ;
        RECT -2.885 222.345 -2.555 222.675 ;
        RECT -2.885 220.675 -2.555 221.005 ;
        RECT -2.885 219.185 -2.555 219.515 ;
        RECT -2.885 217.775 -2.555 218.105 ;
        RECT -2.885 215.935 -2.555 216.265 ;
        RECT -2.885 214.445 -2.555 214.775 ;
        RECT -2.885 212.775 -2.555 213.105 ;
        RECT -2.885 211.285 -2.555 211.615 ;
        RECT -2.885 209.615 -2.555 209.945 ;
        RECT -2.885 208.125 -2.555 208.455 ;
        RECT -2.885 206.455 -2.555 206.785 ;
        RECT -2.885 204.965 -2.555 205.295 ;
        RECT -2.885 203.555 -2.555 203.885 ;
        RECT -2.885 201.715 -2.555 202.045 ;
        RECT -2.885 200.225 -2.555 200.555 ;
        RECT -2.885 198.555 -2.555 198.885 ;
        RECT -2.885 197.065 -2.555 197.395 ;
        RECT -2.885 195.395 -2.555 195.725 ;
        RECT -2.885 193.905 -2.555 194.235 ;
        RECT -2.885 192.235 -2.555 192.565 ;
        RECT -2.885 190.745 -2.555 191.075 ;
        RECT -2.885 189.335 -2.555 189.665 ;
        RECT -2.885 187.495 -2.555 187.825 ;
        RECT -2.885 186.005 -2.555 186.335 ;
        RECT -2.885 184.335 -2.555 184.665 ;
        RECT -2.885 182.845 -2.555 183.175 ;
        RECT -2.885 181.175 -2.555 181.505 ;
        RECT -2.885 179.685 -2.555 180.015 ;
        RECT -2.885 178.015 -2.555 178.345 ;
        RECT -2.885 176.525 -2.555 176.855 ;
        RECT -2.885 175.115 -2.555 175.445 ;
        RECT -2.885 173.275 -2.555 173.605 ;
        RECT -2.885 171.785 -2.555 172.115 ;
        RECT -2.885 170.115 -2.555 170.445 ;
        RECT -2.885 168.625 -2.555 168.955 ;
        RECT -2.885 166.955 -2.555 167.285 ;
        RECT -2.885 165.465 -2.555 165.795 ;
        RECT -2.885 163.795 -2.555 164.125 ;
        RECT -2.885 162.305 -2.555 162.635 ;
        RECT -2.885 160.895 -2.555 161.225 ;
        RECT -2.885 159.055 -2.555 159.385 ;
        RECT -2.885 157.565 -2.555 157.895 ;
        RECT -2.885 155.895 -2.555 156.225 ;
        RECT -2.885 154.405 -2.555 154.735 ;
        RECT -2.885 152.735 -2.555 153.065 ;
        RECT -2.885 151.245 -2.555 151.575 ;
        RECT -2.885 149.575 -2.555 149.905 ;
        RECT -2.885 148.085 -2.555 148.415 ;
        RECT -2.885 146.675 -2.555 147.005 ;
        RECT -2.885 144.835 -2.555 145.165 ;
        RECT -2.885 143.345 -2.555 143.675 ;
        RECT -2.885 141.675 -2.555 142.005 ;
        RECT -2.885 140.185 -2.555 140.515 ;
        RECT -2.885 138.515 -2.555 138.845 ;
        RECT -2.885 137.025 -2.555 137.355 ;
        RECT -2.885 135.355 -2.555 135.685 ;
        RECT -2.885 133.865 -2.555 134.195 ;
        RECT -2.885 132.455 -2.555 132.785 ;
        RECT -2.885 130.615 -2.555 130.945 ;
        RECT -2.885 129.125 -2.555 129.455 ;
        RECT -2.885 127.455 -2.555 127.785 ;
        RECT -2.885 125.965 -2.555 126.295 ;
        RECT -2.885 124.295 -2.555 124.625 ;
        RECT -2.885 122.805 -2.555 123.135 ;
        RECT -2.885 121.135 -2.555 121.465 ;
        RECT -2.885 119.645 -2.555 119.975 ;
        RECT -2.885 118.235 -2.555 118.565 ;
        RECT -2.885 116.395 -2.555 116.725 ;
        RECT -2.885 114.905 -2.555 115.235 ;
        RECT -2.885 113.235 -2.555 113.565 ;
        RECT -2.885 111.745 -2.555 112.075 ;
        RECT -2.885 110.075 -2.555 110.405 ;
        RECT -2.885 108.585 -2.555 108.915 ;
        RECT -2.885 106.915 -2.555 107.245 ;
        RECT -2.885 105.425 -2.555 105.755 ;
        RECT -2.885 104.015 -2.555 104.345 ;
        RECT -2.885 102.175 -2.555 102.505 ;
        RECT -2.885 100.685 -2.555 101.015 ;
        RECT -2.885 99.015 -2.555 99.345 ;
        RECT -2.885 97.525 -2.555 97.855 ;
        RECT -2.885 95.855 -2.555 96.185 ;
        RECT -2.885 94.365 -2.555 94.695 ;
        RECT -2.885 92.695 -2.555 93.025 ;
        RECT -2.885 91.205 -2.555 91.535 ;
        RECT -2.885 89.795 -2.555 90.125 ;
        RECT -2.885 87.955 -2.555 88.285 ;
        RECT -2.885 86.465 -2.555 86.795 ;
        RECT -2.885 84.795 -2.555 85.125 ;
        RECT -2.885 83.305 -2.555 83.635 ;
        RECT -2.885 81.635 -2.555 81.965 ;
        RECT -2.885 80.145 -2.555 80.475 ;
        RECT -2.885 78.475 -2.555 78.805 ;
        RECT -2.885 76.985 -2.555 77.315 ;
        RECT -2.885 75.575 -2.555 75.905 ;
        RECT -2.885 73.735 -2.555 74.065 ;
        RECT -2.885 72.245 -2.555 72.575 ;
        RECT -2.885 70.575 -2.555 70.905 ;
        RECT -2.885 69.085 -2.555 69.415 ;
        RECT -2.885 67.415 -2.555 67.745 ;
        RECT -2.885 65.925 -2.555 66.255 ;
        RECT -2.885 64.255 -2.555 64.585 ;
        RECT -2.885 62.765 -2.555 63.095 ;
        RECT -2.885 61.355 -2.555 61.685 ;
        RECT -2.885 59.515 -2.555 59.845 ;
        RECT -2.885 58.025 -2.555 58.355 ;
        RECT -2.885 56.355 -2.555 56.685 ;
        RECT -2.885 54.865 -2.555 55.195 ;
        RECT -2.885 53.195 -2.555 53.525 ;
        RECT -2.885 51.705 -2.555 52.035 ;
        RECT -2.885 50.035 -2.555 50.365 ;
        RECT -2.885 48.545 -2.555 48.875 ;
        RECT -2.885 47.135 -2.555 47.465 ;
        RECT -2.885 45.295 -2.555 45.625 ;
        RECT -2.885 43.805 -2.555 44.135 ;
        RECT -2.885 42.135 -2.555 42.465 ;
        RECT -2.885 40.645 -2.555 40.975 ;
        RECT -2.885 38.975 -2.555 39.305 ;
        RECT -2.885 37.485 -2.555 37.815 ;
        RECT -2.885 35.815 -2.555 36.145 ;
        RECT -2.885 34.325 -2.555 34.655 ;
        RECT -2.885 32.915 -2.555 33.245 ;
        RECT -2.885 31.075 -2.555 31.405 ;
        RECT -2.885 29.585 -2.555 29.915 ;
        RECT -2.885 27.915 -2.555 28.245 ;
        RECT -2.885 26.425 -2.555 26.755 ;
        RECT -2.885 24.755 -2.555 25.085 ;
        RECT -2.885 23.265 -2.555 23.595 ;
        RECT -2.885 21.595 -2.555 21.925 ;
        RECT -2.885 20.105 -2.555 20.435 ;
        RECT -2.885 18.695 -2.555 19.025 ;
        RECT -2.885 16.855 -2.555 17.185 ;
        RECT -2.885 15.365 -2.555 15.695 ;
        RECT -2.885 13.695 -2.555 14.025 ;
        RECT -2.885 12.205 -2.555 12.535 ;
        RECT -2.885 10.535 -2.555 10.865 ;
        RECT -2.885 9.045 -2.555 9.375 ;
        RECT -2.885 7.375 -2.555 7.705 ;
        RECT -2.885 5.885 -2.555 6.215 ;
        RECT -2.885 4.475 -2.555 4.805 ;
        RECT -2.885 2.115 -2.555 2.445 ;
        RECT -2.885 0.06 -2.555 0.39 ;
        RECT -2.885 -1.525 -2.555 -1.195 ;
        RECT -2.885 -2.885 -2.555 -2.555 ;
        RECT -2.885 -4.245 -2.555 -3.915 ;
        RECT -2.885 -5.605 -2.555 -5.275 ;
        RECT -2.885 -6.965 -2.555 -6.635 ;
        RECT -2.885 -8.325 -2.555 -7.995 ;
        RECT -2.885 -9.685 -2.555 -9.355 ;
        RECT -2.885 -12.405 -2.555 -12.075 ;
        RECT -2.885 -13.765 -2.555 -13.435 ;
        RECT -2.885 -15.125 -2.555 -14.795 ;
        RECT -2.885 -16.485 -2.555 -16.155 ;
        RECT -2.885 -17.845 -2.555 -17.515 ;
        RECT -2.885 -21.925 -2.555 -21.595 ;
        RECT -2.885 -23.285 -2.555 -22.955 ;
        RECT -2.885 -24.645 -2.555 -24.315 ;
        RECT -2.885 -26.005 -2.555 -25.675 ;
        RECT -2.885 -27.365 -2.555 -27.035 ;
        RECT -2.885 -28.725 -2.555 -28.395 ;
        RECT -2.885 -30.085 -2.555 -29.755 ;
        RECT -2.885 -31.445 -2.555 -31.115 ;
        RECT -2.885 -32.805 -2.555 -32.475 ;
        RECT -2.885 -34.165 -2.555 -33.835 ;
        RECT -2.885 -36.885 -2.555 -36.555 ;
        RECT -2.885 -38.245 -2.555 -37.915 ;
        RECT -2.885 -40.965 -2.555 -40.635 ;
        RECT -2.885 -42.325 -2.555 -41.995 ;
        RECT -2.885 -43.685 -2.555 -43.355 ;
        RECT -2.885 -45.045 -2.555 -44.715 ;
        RECT -2.885 -46.405 -2.555 -46.075 ;
        RECT -2.885 -47.765 -2.555 -47.435 ;
        RECT -2.885 -49.125 -2.555 -48.795 ;
        RECT -2.885 -51.845 -2.555 -51.515 ;
        RECT -2.885 -53.205 -2.555 -52.875 ;
        RECT -2.885 -54.565 -2.555 -54.235 ;
        RECT -2.885 -55.925 -2.555 -55.595 ;
        RECT -2.885 -57.285 -2.555 -56.955 ;
        RECT -2.885 -58.645 -2.555 -58.315 ;
        RECT -2.885 -60.005 -2.555 -59.675 ;
        RECT -2.885 -61.365 -2.555 -61.035 ;
        RECT -2.885 -62.725 -2.555 -62.395 ;
        RECT -2.885 -64.085 -2.555 -63.755 ;
        RECT -2.885 -65.445 -2.555 -65.115 ;
        RECT -2.885 -66.805 -2.555 -66.475 ;
        RECT -2.885 -68.165 -2.555 -67.835 ;
        RECT -2.885 -69.525 -2.555 -69.195 ;
        RECT -2.885 -70.885 -2.555 -70.555 ;
        RECT -2.885 -72.245 -2.555 -71.915 ;
        RECT -2.885 -73.605 -2.555 -73.275 ;
        RECT -2.885 -74.965 -2.555 -74.635 ;
        RECT -2.885 -76.325 -2.555 -75.995 ;
        RECT -2.885 -77.685 -2.555 -77.355 ;
        RECT -2.885 -79.045 -2.555 -78.715 ;
        RECT -2.885 -80.405 -2.555 -80.075 ;
        RECT -2.885 -81.765 -2.555 -81.435 ;
        RECT -2.885 -83.125 -2.555 -82.795 ;
        RECT -2.885 -84.485 -2.555 -84.155 ;
        RECT -2.885 -85.845 -2.555 -85.515 ;
        RECT -2.885 -87.205 -2.555 -86.875 ;
        RECT -2.885 -88.565 -2.555 -88.235 ;
        RECT -2.885 -89.925 -2.555 -89.595 ;
        RECT -2.885 -91.285 -2.555 -90.955 ;
        RECT -2.885 -92.645 -2.555 -92.315 ;
        RECT -2.885 -94.005 -2.555 -93.675 ;
        RECT -2.885 -95.365 -2.555 -95.035 ;
        RECT -2.885 -96.725 -2.555 -96.395 ;
        RECT -2.885 -98.085 -2.555 -97.755 ;
        RECT -2.885 -99.445 -2.555 -99.115 ;
        RECT -2.885 -100.805 -2.555 -100.475 ;
        RECT -2.885 -102.165 -2.555 -101.835 ;
        RECT -2.885 -103.525 -2.555 -103.195 ;
        RECT -2.885 -104.885 -2.555 -104.555 ;
        RECT -2.885 -106.245 -2.555 -105.915 ;
        RECT -2.885 -107.605 -2.555 -107.275 ;
        RECT -2.885 -108.965 -2.555 -108.635 ;
        RECT -2.885 -110.325 -2.555 -109.995 ;
        RECT -2.885 -111.685 -2.555 -111.355 ;
        RECT -2.885 -113.045 -2.555 -112.715 ;
        RECT -2.885 -114.405 -2.555 -114.075 ;
        RECT -2.885 -115.765 -2.555 -115.435 ;
        RECT -2.885 -117.125 -2.555 -116.795 ;
        RECT -2.885 -119.845 -2.555 -119.515 ;
        RECT -2.885 -121.205 -2.555 -120.875 ;
        RECT -2.885 -122.565 -2.555 -122.235 ;
        RECT -2.885 -123.925 -2.555 -123.595 ;
        RECT -2.885 -125.285 -2.555 -124.955 ;
        RECT -2.885 -126.645 -2.555 -126.315 ;
        RECT -2.885 -128.005 -2.555 -127.675 ;
        RECT -2.885 -129.365 -2.555 -129.035 ;
        RECT -2.885 -130.725 -2.555 -130.395 ;
        RECT -2.885 -132.085 -2.555 -131.755 ;
        RECT -2.885 -133.445 -2.555 -133.115 ;
        RECT -2.885 -134.805 -2.555 -134.475 ;
        RECT -2.885 -136.165 -2.555 -135.835 ;
        RECT -2.885 -137.525 -2.555 -137.195 ;
        RECT -2.885 -138.885 -2.555 -138.555 ;
        RECT -2.885 -140.245 -2.555 -139.915 ;
        RECT -2.885 -141.605 -2.555 -141.275 ;
        RECT -2.885 -142.965 -2.555 -142.635 ;
        RECT -2.885 -144.325 -2.555 -143.995 ;
        RECT -2.885 -145.685 -2.555 -145.355 ;
        RECT -2.885 -147.045 -2.555 -146.715 ;
        RECT -2.885 -148.405 -2.555 -148.075 ;
        RECT -2.885 -149.765 -2.555 -149.435 ;
        RECT -2.885 -151.125 -2.555 -150.795 ;
        RECT -2.885 -152.485 -2.555 -152.155 ;
        RECT -2.885 -153.845 -2.555 -153.515 ;
        RECT -2.885 -155.205 -2.555 -154.875 ;
        RECT -2.885 -156.565 -2.555 -156.235 ;
        RECT -2.885 -157.925 -2.555 -157.595 ;
        RECT -2.885 -159.285 -2.555 -158.955 ;
        RECT -2.885 -160.645 -2.555 -160.315 ;
        RECT -2.885 -162.005 -2.555 -161.675 ;
        RECT -2.885 -163.365 -2.555 -163.035 ;
        RECT -2.885 -164.725 -2.555 -164.395 ;
        RECT -2.885 -166.085 -2.555 -165.755 ;
        RECT -2.885 -167.445 -2.555 -167.115 ;
        RECT -2.885 -168.805 -2.555 -168.475 ;
        RECT -2.885 -170.165 -2.555 -169.835 ;
        RECT -2.885 -171.525 -2.555 -171.195 ;
        RECT -2.885 -172.885 -2.555 -172.555 ;
        RECT -2.885 -174.245 -2.555 -173.915 ;
        RECT -2.885 -175.605 -2.555 -175.275 ;
        RECT -2.885 -176.965 -2.555 -176.635 ;
        RECT -2.885 -178.325 -2.555 -177.995 ;
        RECT -2.885 -180.57 -2.555 -179.44 ;
        RECT -2.88 -180.685 -2.56 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -1.525 146.675 -1.195 147.005 ;
        RECT -1.525 144.835 -1.195 145.165 ;
        RECT -1.525 143.345 -1.195 143.675 ;
        RECT -1.525 141.675 -1.195 142.005 ;
        RECT -1.525 140.185 -1.195 140.515 ;
        RECT -1.525 138.515 -1.195 138.845 ;
        RECT -1.525 137.025 -1.195 137.355 ;
        RECT -1.525 135.355 -1.195 135.685 ;
        RECT -1.525 133.865 -1.195 134.195 ;
        RECT -1.525 132.455 -1.195 132.785 ;
        RECT -1.525 130.615 -1.195 130.945 ;
        RECT -1.525 129.125 -1.195 129.455 ;
        RECT -1.525 127.455 -1.195 127.785 ;
        RECT -1.525 125.965 -1.195 126.295 ;
        RECT -1.525 124.295 -1.195 124.625 ;
        RECT -1.525 122.805 -1.195 123.135 ;
        RECT -1.525 121.135 -1.195 121.465 ;
        RECT -1.525 119.645 -1.195 119.975 ;
        RECT -1.525 118.235 -1.195 118.565 ;
        RECT -1.525 116.395 -1.195 116.725 ;
        RECT -1.525 114.905 -1.195 115.235 ;
        RECT -1.525 113.235 -1.195 113.565 ;
        RECT -1.525 111.745 -1.195 112.075 ;
        RECT -1.525 110.075 -1.195 110.405 ;
        RECT -1.525 108.585 -1.195 108.915 ;
        RECT -1.525 106.915 -1.195 107.245 ;
        RECT -1.525 105.425 -1.195 105.755 ;
        RECT -1.525 104.015 -1.195 104.345 ;
        RECT -1.525 102.175 -1.195 102.505 ;
        RECT -1.525 100.685 -1.195 101.015 ;
        RECT -1.525 99.015 -1.195 99.345 ;
        RECT -1.525 97.525 -1.195 97.855 ;
        RECT -1.525 95.855 -1.195 96.185 ;
        RECT -1.525 94.365 -1.195 94.695 ;
        RECT -1.525 92.695 -1.195 93.025 ;
        RECT -1.525 91.205 -1.195 91.535 ;
        RECT -1.525 89.795 -1.195 90.125 ;
        RECT -1.525 87.955 -1.195 88.285 ;
        RECT -1.525 86.465 -1.195 86.795 ;
        RECT -1.525 84.795 -1.195 85.125 ;
        RECT -1.525 83.305 -1.195 83.635 ;
        RECT -1.525 81.635 -1.195 81.965 ;
        RECT -1.525 80.145 -1.195 80.475 ;
        RECT -1.525 78.475 -1.195 78.805 ;
        RECT -1.525 76.985 -1.195 77.315 ;
        RECT -1.525 75.575 -1.195 75.905 ;
        RECT -1.525 73.735 -1.195 74.065 ;
        RECT -1.525 72.245 -1.195 72.575 ;
        RECT -1.525 70.575 -1.195 70.905 ;
        RECT -1.525 69.085 -1.195 69.415 ;
        RECT -1.525 67.415 -1.195 67.745 ;
        RECT -1.525 65.925 -1.195 66.255 ;
        RECT -1.525 64.255 -1.195 64.585 ;
        RECT -1.525 62.765 -1.195 63.095 ;
        RECT -1.525 61.355 -1.195 61.685 ;
        RECT -1.525 59.515 -1.195 59.845 ;
        RECT -1.525 58.025 -1.195 58.355 ;
        RECT -1.525 56.355 -1.195 56.685 ;
        RECT -1.525 54.865 -1.195 55.195 ;
        RECT -1.525 53.195 -1.195 53.525 ;
        RECT -1.525 51.705 -1.195 52.035 ;
        RECT -1.525 50.035 -1.195 50.365 ;
        RECT -1.525 48.545 -1.195 48.875 ;
        RECT -1.525 47.135 -1.195 47.465 ;
        RECT -1.525 45.295 -1.195 45.625 ;
        RECT -1.525 43.805 -1.195 44.135 ;
        RECT -1.525 42.135 -1.195 42.465 ;
        RECT -1.525 40.645 -1.195 40.975 ;
        RECT -1.525 38.975 -1.195 39.305 ;
        RECT -1.525 37.485 -1.195 37.815 ;
        RECT -1.525 35.815 -1.195 36.145 ;
        RECT -1.525 34.325 -1.195 34.655 ;
        RECT -1.525 32.915 -1.195 33.245 ;
        RECT -1.525 31.075 -1.195 31.405 ;
        RECT -1.525 29.585 -1.195 29.915 ;
        RECT -1.525 27.915 -1.195 28.245 ;
        RECT -1.525 26.425 -1.195 26.755 ;
        RECT -1.525 24.755 -1.195 25.085 ;
        RECT -1.525 23.265 -1.195 23.595 ;
        RECT -1.525 21.595 -1.195 21.925 ;
        RECT -1.525 20.105 -1.195 20.435 ;
        RECT -1.525 18.695 -1.195 19.025 ;
        RECT -1.525 16.855 -1.195 17.185 ;
        RECT -1.525 15.365 -1.195 15.695 ;
        RECT -1.525 13.695 -1.195 14.025 ;
        RECT -1.525 12.205 -1.195 12.535 ;
        RECT -1.525 10.535 -1.195 10.865 ;
        RECT -1.525 9.045 -1.195 9.375 ;
        RECT -1.525 7.375 -1.195 7.705 ;
        RECT -1.525 5.885 -1.195 6.215 ;
        RECT -1.525 4.475 -1.195 4.805 ;
        RECT -1.525 2.115 -1.195 2.445 ;
        RECT -1.525 0.06 -1.195 0.39 ;
        RECT -1.525 -1.525 -1.195 -1.195 ;
        RECT -1.525 -2.885 -1.195 -2.555 ;
        RECT -1.525 -4.245 -1.195 -3.915 ;
        RECT -1.525 -5.605 -1.195 -5.275 ;
        RECT -1.525 -6.965 -1.195 -6.635 ;
        RECT -1.525 -8.325 -1.195 -7.995 ;
        RECT -1.525 -9.685 -1.195 -9.355 ;
        RECT -1.525 -12.405 -1.195 -12.075 ;
        RECT -1.525 -13.765 -1.195 -13.435 ;
        RECT -1.525 -15.125 -1.195 -14.795 ;
        RECT -1.525 -16.485 -1.195 -16.155 ;
        RECT -1.525 -17.845 -1.195 -17.515 ;
        RECT -1.525 -21.925 -1.195 -21.595 ;
        RECT -1.525 -23.285 -1.195 -22.955 ;
        RECT -1.525 -24.645 -1.195 -24.315 ;
        RECT -1.525 -26.005 -1.195 -25.675 ;
        RECT -1.525 -27.365 -1.195 -27.035 ;
        RECT -1.525 -28.725 -1.195 -28.395 ;
        RECT -1.525 -30.085 -1.195 -29.755 ;
        RECT -1.525 -31.445 -1.195 -31.115 ;
        RECT -1.525 -32.805 -1.195 -32.475 ;
        RECT -1.525 -34.165 -1.195 -33.835 ;
        RECT -1.525 -36.885 -1.195 -36.555 ;
        RECT -1.525 -38.245 -1.195 -37.915 ;
        RECT -1.525 -40.965 -1.195 -40.635 ;
        RECT -1.525 -42.325 -1.195 -41.995 ;
        RECT -1.525 -43.685 -1.195 -43.355 ;
        RECT -1.525 -45.045 -1.195 -44.715 ;
        RECT -1.525 -46.405 -1.195 -46.075 ;
        RECT -1.525 -47.765 -1.195 -47.435 ;
        RECT -1.525 -49.125 -1.195 -48.795 ;
        RECT -1.525 -51.845 -1.195 -51.515 ;
        RECT -1.525 -53.205 -1.195 -52.875 ;
        RECT -1.525 -54.565 -1.195 -54.235 ;
        RECT -1.525 -55.925 -1.195 -55.595 ;
        RECT -1.525 -57.285 -1.195 -56.955 ;
        RECT -1.525 -58.645 -1.195 -58.315 ;
        RECT -1.525 -60.005 -1.195 -59.675 ;
        RECT -1.525 -61.365 -1.195 -61.035 ;
        RECT -1.525 -62.725 -1.195 -62.395 ;
        RECT -1.525 -64.085 -1.195 -63.755 ;
        RECT -1.525 -65.445 -1.195 -65.115 ;
        RECT -1.525 -66.805 -1.195 -66.475 ;
        RECT -1.525 -68.165 -1.195 -67.835 ;
        RECT -1.525 -69.525 -1.195 -69.195 ;
        RECT -1.525 -70.885 -1.195 -70.555 ;
        RECT -1.525 -72.245 -1.195 -71.915 ;
        RECT -1.525 -73.605 -1.195 -73.275 ;
        RECT -1.525 -74.965 -1.195 -74.635 ;
        RECT -1.525 -76.325 -1.195 -75.995 ;
        RECT -1.525 -77.685 -1.195 -77.355 ;
        RECT -1.525 -79.045 -1.195 -78.715 ;
        RECT -1.525 -80.405 -1.195 -80.075 ;
        RECT -1.525 -81.765 -1.195 -81.435 ;
        RECT -1.525 -83.125 -1.195 -82.795 ;
        RECT -1.525 -84.485 -1.195 -84.155 ;
        RECT -1.525 -85.845 -1.195 -85.515 ;
        RECT -1.525 -87.205 -1.195 -86.875 ;
        RECT -1.525 -88.565 -1.195 -88.235 ;
        RECT -1.525 -89.925 -1.195 -89.595 ;
        RECT -1.525 -91.285 -1.195 -90.955 ;
        RECT -1.525 -92.645 -1.195 -92.315 ;
        RECT -1.525 -94.005 -1.195 -93.675 ;
        RECT -1.525 -95.365 -1.195 -95.035 ;
        RECT -1.525 -96.725 -1.195 -96.395 ;
        RECT -1.525 -98.085 -1.195 -97.755 ;
        RECT -1.525 -99.445 -1.195 -99.115 ;
        RECT -1.525 -100.805 -1.195 -100.475 ;
        RECT -1.525 -102.165 -1.195 -101.835 ;
        RECT -1.525 -103.525 -1.195 -103.195 ;
        RECT -1.525 -104.885 -1.195 -104.555 ;
        RECT -1.525 -106.245 -1.195 -105.915 ;
        RECT -1.525 -107.605 -1.195 -107.275 ;
        RECT -1.525 -108.965 -1.195 -108.635 ;
        RECT -1.525 -110.325 -1.195 -109.995 ;
        RECT -1.525 -111.685 -1.195 -111.355 ;
        RECT -1.525 -113.045 -1.195 -112.715 ;
        RECT -1.525 -114.405 -1.195 -114.075 ;
        RECT -1.525 -115.765 -1.195 -115.435 ;
        RECT -1.525 -117.125 -1.195 -116.795 ;
        RECT -1.525 -119.845 -1.195 -119.515 ;
        RECT -1.525 -121.205 -1.195 -120.875 ;
        RECT -1.525 -122.565 -1.195 -122.235 ;
        RECT -1.525 -123.925 -1.195 -123.595 ;
        RECT -1.525 -125.285 -1.195 -124.955 ;
        RECT -1.525 -126.645 -1.195 -126.315 ;
        RECT -1.525 -128.005 -1.195 -127.675 ;
        RECT -1.525 -129.365 -1.195 -129.035 ;
        RECT -1.525 -130.725 -1.195 -130.395 ;
        RECT -1.525 -132.085 -1.195 -131.755 ;
        RECT -1.525 -133.445 -1.195 -133.115 ;
        RECT -1.525 -134.805 -1.195 -134.475 ;
        RECT -1.525 -136.165 -1.195 -135.835 ;
        RECT -1.525 -137.525 -1.195 -137.195 ;
        RECT -1.525 -138.885 -1.195 -138.555 ;
        RECT -1.525 -140.245 -1.195 -139.915 ;
        RECT -1.525 -141.605 -1.195 -141.275 ;
        RECT -1.525 -142.965 -1.195 -142.635 ;
        RECT -1.525 -144.325 -1.195 -143.995 ;
        RECT -1.525 -145.685 -1.195 -145.355 ;
        RECT -1.525 -147.045 -1.195 -146.715 ;
        RECT -1.525 -148.405 -1.195 -148.075 ;
        RECT -1.525 -149.765 -1.195 -149.435 ;
        RECT -1.525 -151.125 -1.195 -150.795 ;
        RECT -1.525 -152.485 -1.195 -152.155 ;
        RECT -1.525 -153.845 -1.195 -153.515 ;
        RECT -1.525 -155.205 -1.195 -154.875 ;
        RECT -1.525 -156.565 -1.195 -156.235 ;
        RECT -1.525 -157.925 -1.195 -157.595 ;
        RECT -1.525 -159.285 -1.195 -158.955 ;
        RECT -1.525 -160.645 -1.195 -160.315 ;
        RECT -1.525 -162.005 -1.195 -161.675 ;
        RECT -1.525 -163.365 -1.195 -163.035 ;
        RECT -1.525 -164.725 -1.195 -164.395 ;
        RECT -1.525 -166.085 -1.195 -165.755 ;
        RECT -1.525 -167.445 -1.195 -167.115 ;
        RECT -1.525 -168.805 -1.195 -168.475 ;
        RECT -1.525 -170.165 -1.195 -169.835 ;
        RECT -1.525 -171.525 -1.195 -171.195 ;
        RECT -1.525 -172.885 -1.195 -172.555 ;
        RECT -1.525 -174.245 -1.195 -173.915 ;
        RECT -1.525 -175.605 -1.195 -175.275 ;
        RECT -1.525 -176.965 -1.195 -176.635 ;
        RECT -1.525 -178.325 -1.195 -177.995 ;
        RECT -1.525 -180.57 -1.195 -179.44 ;
        RECT -1.52 -180.685 -1.2 242.565 ;
        RECT -1.525 241.32 -1.195 242.45 ;
        RECT -1.525 239.195 -1.195 239.525 ;
        RECT -1.525 237.835 -1.195 238.165 ;
        RECT -1.525 235.975 -1.195 236.305 ;
        RECT -1.525 233.925 -1.195 234.255 ;
        RECT -1.525 231.995 -1.195 232.325 ;
        RECT -1.525 230.155 -1.195 230.485 ;
        RECT -1.525 228.665 -1.195 228.995 ;
        RECT -1.525 226.995 -1.195 227.325 ;
        RECT -1.525 225.505 -1.195 225.835 ;
        RECT -1.525 223.835 -1.195 224.165 ;
        RECT -1.525 222.345 -1.195 222.675 ;
        RECT -1.525 220.675 -1.195 221.005 ;
        RECT -1.525 219.185 -1.195 219.515 ;
        RECT -1.525 217.775 -1.195 218.105 ;
        RECT -1.525 215.935 -1.195 216.265 ;
        RECT -1.525 214.445 -1.195 214.775 ;
        RECT -1.525 212.775 -1.195 213.105 ;
        RECT -1.525 211.285 -1.195 211.615 ;
        RECT -1.525 209.615 -1.195 209.945 ;
        RECT -1.525 208.125 -1.195 208.455 ;
        RECT -1.525 206.455 -1.195 206.785 ;
        RECT -1.525 204.965 -1.195 205.295 ;
        RECT -1.525 203.555 -1.195 203.885 ;
        RECT -1.525 201.715 -1.195 202.045 ;
        RECT -1.525 200.225 -1.195 200.555 ;
        RECT -1.525 198.555 -1.195 198.885 ;
        RECT -1.525 197.065 -1.195 197.395 ;
        RECT -1.525 195.395 -1.195 195.725 ;
        RECT -1.525 193.905 -1.195 194.235 ;
        RECT -1.525 192.235 -1.195 192.565 ;
        RECT -1.525 190.745 -1.195 191.075 ;
        RECT -1.525 189.335 -1.195 189.665 ;
        RECT -1.525 187.495 -1.195 187.825 ;
        RECT -1.525 186.005 -1.195 186.335 ;
        RECT -1.525 184.335 -1.195 184.665 ;
        RECT -1.525 182.845 -1.195 183.175 ;
        RECT -1.525 181.175 -1.195 181.505 ;
        RECT -1.525 179.685 -1.195 180.015 ;
        RECT -1.525 178.015 -1.195 178.345 ;
        RECT -1.525 176.525 -1.195 176.855 ;
        RECT -1.525 175.115 -1.195 175.445 ;
        RECT -1.525 173.275 -1.195 173.605 ;
        RECT -1.525 171.785 -1.195 172.115 ;
        RECT -1.525 170.115 -1.195 170.445 ;
        RECT -1.525 168.625 -1.195 168.955 ;
        RECT -1.525 166.955 -1.195 167.285 ;
        RECT -1.525 165.465 -1.195 165.795 ;
        RECT -1.525 163.795 -1.195 164.125 ;
        RECT -1.525 162.305 -1.195 162.635 ;
        RECT -1.525 160.895 -1.195 161.225 ;
        RECT -1.525 159.055 -1.195 159.385 ;
        RECT -1.525 157.565 -1.195 157.895 ;
        RECT -1.525 155.895 -1.195 156.225 ;
        RECT -1.525 154.405 -1.195 154.735 ;
        RECT -1.525 152.735 -1.195 153.065 ;
        RECT -1.525 151.245 -1.195 151.575 ;
        RECT -1.525 149.575 -1.195 149.905 ;
        RECT -1.525 148.085 -1.195 148.415 ;
    END
    PORT
      LAYER met3 ;
        RECT -12.405 241.32 -12.075 242.45 ;
        RECT -12.405 239.195 -12.075 239.525 ;
        RECT -12.405 237.835 -12.075 238.165 ;
        RECT -12.405 236.475 -12.075 236.805 ;
        RECT -12.405 235.115 -12.075 235.445 ;
        RECT -12.405 233.755 -12.075 234.085 ;
        RECT -12.405 232.395 -12.075 232.725 ;
        RECT -12.405 231.035 -12.075 231.365 ;
        RECT -12.405 229.675 -12.075 230.005 ;
        RECT -12.405 228.315 -12.075 228.645 ;
        RECT -12.405 226.955 -12.075 227.285 ;
        RECT -12.405 225.595 -12.075 225.925 ;
        RECT -12.405 224.235 -12.075 224.565 ;
        RECT -12.405 222.875 -12.075 223.205 ;
        RECT -12.405 221.515 -12.075 221.845 ;
        RECT -12.405 220.155 -12.075 220.485 ;
        RECT -12.405 218.795 -12.075 219.125 ;
        RECT -12.405 217.435 -12.075 217.765 ;
        RECT -12.405 216.075 -12.075 216.405 ;
        RECT -12.405 214.715 -12.075 215.045 ;
        RECT -12.405 213.355 -12.075 213.685 ;
        RECT -12.405 211.995 -12.075 212.325 ;
        RECT -12.405 210.635 -12.075 210.965 ;
        RECT -12.405 209.275 -12.075 209.605 ;
        RECT -12.405 207.915 -12.075 208.245 ;
        RECT -12.405 206.555 -12.075 206.885 ;
        RECT -12.405 205.195 -12.075 205.525 ;
        RECT -12.405 203.835 -12.075 204.165 ;
        RECT -12.405 202.475 -12.075 202.805 ;
        RECT -12.405 201.115 -12.075 201.445 ;
        RECT -12.405 199.755 -12.075 200.085 ;
        RECT -12.405 198.395 -12.075 198.725 ;
        RECT -12.405 197.035 -12.075 197.365 ;
        RECT -12.405 195.675 -12.075 196.005 ;
        RECT -12.405 194.315 -12.075 194.645 ;
        RECT -12.405 192.955 -12.075 193.285 ;
        RECT -12.405 191.595 -12.075 191.925 ;
        RECT -12.405 190.235 -12.075 190.565 ;
        RECT -12.405 188.875 -12.075 189.205 ;
        RECT -12.405 187.515 -12.075 187.845 ;
        RECT -12.405 186.155 -12.075 186.485 ;
        RECT -12.405 184.795 -12.075 185.125 ;
        RECT -12.405 183.435 -12.075 183.765 ;
        RECT -12.405 182.075 -12.075 182.405 ;
        RECT -12.405 180.715 -12.075 181.045 ;
        RECT -12.405 179.355 -12.075 179.685 ;
        RECT -12.405 177.995 -12.075 178.325 ;
        RECT -12.405 176.635 -12.075 176.965 ;
        RECT -12.405 175.275 -12.075 175.605 ;
        RECT -12.405 173.915 -12.075 174.245 ;
        RECT -12.405 172.555 -12.075 172.885 ;
        RECT -12.405 171.195 -12.075 171.525 ;
        RECT -12.405 169.835 -12.075 170.165 ;
        RECT -12.405 168.475 -12.075 168.805 ;
        RECT -12.405 167.115 -12.075 167.445 ;
        RECT -12.405 165.755 -12.075 166.085 ;
        RECT -12.405 164.395 -12.075 164.725 ;
        RECT -12.405 163.035 -12.075 163.365 ;
        RECT -12.405 161.675 -12.075 162.005 ;
        RECT -12.405 160.315 -12.075 160.645 ;
        RECT -12.405 158.955 -12.075 159.285 ;
        RECT -12.405 157.595 -12.075 157.925 ;
        RECT -12.405 156.235 -12.075 156.565 ;
        RECT -12.405 154.875 -12.075 155.205 ;
        RECT -12.405 153.515 -12.075 153.845 ;
        RECT -12.405 152.155 -12.075 152.485 ;
        RECT -12.405 150.795 -12.075 151.125 ;
        RECT -12.405 149.435 -12.075 149.765 ;
        RECT -12.405 148.075 -12.075 148.405 ;
        RECT -12.405 146.715 -12.075 147.045 ;
        RECT -12.405 145.355 -12.075 145.685 ;
        RECT -12.405 143.995 -12.075 144.325 ;
        RECT -12.405 142.635 -12.075 142.965 ;
        RECT -12.405 141.275 -12.075 141.605 ;
        RECT -12.405 139.915 -12.075 140.245 ;
        RECT -12.405 138.555 -12.075 138.885 ;
        RECT -12.405 137.195 -12.075 137.525 ;
        RECT -12.405 135.835 -12.075 136.165 ;
        RECT -12.405 134.475 -12.075 134.805 ;
        RECT -12.405 133.115 -12.075 133.445 ;
        RECT -12.405 131.755 -12.075 132.085 ;
        RECT -12.405 130.395 -12.075 130.725 ;
        RECT -12.405 129.035 -12.075 129.365 ;
        RECT -12.405 127.675 -12.075 128.005 ;
        RECT -12.405 126.315 -12.075 126.645 ;
        RECT -12.405 124.955 -12.075 125.285 ;
        RECT -12.405 123.595 -12.075 123.925 ;
        RECT -12.405 122.235 -12.075 122.565 ;
        RECT -12.405 120.875 -12.075 121.205 ;
        RECT -12.405 119.515 -12.075 119.845 ;
        RECT -12.405 118.155 -12.075 118.485 ;
        RECT -12.405 116.795 -12.075 117.125 ;
        RECT -12.405 115.435 -12.075 115.765 ;
        RECT -12.405 114.075 -12.075 114.405 ;
        RECT -12.405 112.715 -12.075 113.045 ;
        RECT -12.405 111.355 -12.075 111.685 ;
        RECT -12.405 109.995 -12.075 110.325 ;
        RECT -12.405 108.635 -12.075 108.965 ;
        RECT -12.405 107.275 -12.075 107.605 ;
        RECT -12.405 105.915 -12.075 106.245 ;
        RECT -12.405 104.555 -12.075 104.885 ;
        RECT -12.405 103.195 -12.075 103.525 ;
        RECT -12.405 101.835 -12.075 102.165 ;
        RECT -12.405 100.475 -12.075 100.805 ;
        RECT -12.405 99.115 -12.075 99.445 ;
        RECT -12.405 97.755 -12.075 98.085 ;
        RECT -12.405 96.395 -12.075 96.725 ;
        RECT -12.405 95.035 -12.075 95.365 ;
        RECT -12.405 93.675 -12.075 94.005 ;
        RECT -12.405 92.315 -12.075 92.645 ;
        RECT -12.405 90.955 -12.075 91.285 ;
        RECT -12.405 89.595 -12.075 89.925 ;
        RECT -12.405 88.235 -12.075 88.565 ;
        RECT -12.405 86.875 -12.075 87.205 ;
        RECT -12.405 85.515 -12.075 85.845 ;
        RECT -12.405 84.155 -12.075 84.485 ;
        RECT -12.405 82.795 -12.075 83.125 ;
        RECT -12.405 81.435 -12.075 81.765 ;
        RECT -12.405 80.075 -12.075 80.405 ;
        RECT -12.405 78.715 -12.075 79.045 ;
        RECT -12.405 77.355 -12.075 77.685 ;
        RECT -12.405 75.995 -12.075 76.325 ;
        RECT -12.405 74.635 -12.075 74.965 ;
        RECT -12.405 73.275 -12.075 73.605 ;
        RECT -12.405 71.915 -12.075 72.245 ;
        RECT -12.405 70.555 -12.075 70.885 ;
        RECT -12.405 69.195 -12.075 69.525 ;
        RECT -12.405 67.835 -12.075 68.165 ;
        RECT -12.405 66.475 -12.075 66.805 ;
        RECT -12.405 65.115 -12.075 65.445 ;
        RECT -12.405 63.755 -12.075 64.085 ;
        RECT -12.405 62.395 -12.075 62.725 ;
        RECT -12.405 61.035 -12.075 61.365 ;
        RECT -12.405 59.675 -12.075 60.005 ;
        RECT -12.405 58.315 -12.075 58.645 ;
        RECT -12.405 56.955 -12.075 57.285 ;
        RECT -12.405 55.595 -12.075 55.925 ;
        RECT -12.405 54.235 -12.075 54.565 ;
        RECT -12.405 52.875 -12.075 53.205 ;
        RECT -12.405 51.515 -12.075 51.845 ;
        RECT -12.405 50.155 -12.075 50.485 ;
        RECT -12.405 48.795 -12.075 49.125 ;
        RECT -12.405 47.435 -12.075 47.765 ;
        RECT -12.405 46.075 -12.075 46.405 ;
        RECT -12.405 44.715 -12.075 45.045 ;
        RECT -12.405 43.355 -12.075 43.685 ;
        RECT -12.405 41.995 -12.075 42.325 ;
        RECT -12.405 40.635 -12.075 40.965 ;
        RECT -12.405 39.275 -12.075 39.605 ;
        RECT -12.405 37.915 -12.075 38.245 ;
        RECT -12.405 36.555 -12.075 36.885 ;
        RECT -12.405 35.195 -12.075 35.525 ;
        RECT -12.405 33.835 -12.075 34.165 ;
        RECT -12.405 32.475 -12.075 32.805 ;
        RECT -12.405 31.115 -12.075 31.445 ;
        RECT -12.405 29.755 -12.075 30.085 ;
        RECT -12.405 28.395 -12.075 28.725 ;
        RECT -12.405 27.035 -12.075 27.365 ;
        RECT -12.405 25.675 -12.075 26.005 ;
        RECT -12.405 24.315 -12.075 24.645 ;
        RECT -12.405 22.955 -12.075 23.285 ;
        RECT -12.405 21.595 -12.075 21.925 ;
        RECT -12.405 20.235 -12.075 20.565 ;
        RECT -12.405 18.875 -12.075 19.205 ;
        RECT -12.405 17.515 -12.075 17.845 ;
        RECT -12.405 16.155 -12.075 16.485 ;
        RECT -12.405 14.795 -12.075 15.125 ;
        RECT -12.405 13.435 -12.075 13.765 ;
        RECT -12.405 12.075 -12.075 12.405 ;
        RECT -12.405 10.715 -12.075 11.045 ;
        RECT -12.405 9.355 -12.075 9.685 ;
        RECT -12.405 7.995 -12.075 8.325 ;
        RECT -12.405 6.635 -12.075 6.965 ;
        RECT -12.405 5.275 -12.075 5.605 ;
        RECT -12.405 3.915 -12.075 4.245 ;
        RECT -12.405 2.555 -12.075 2.885 ;
        RECT -12.405 1.195 -12.075 1.525 ;
        RECT -12.405 -0.165 -12.075 0.165 ;
        RECT -12.405 -2.885 -12.075 -2.555 ;
        RECT -12.405 -4.245 -12.075 -3.915 ;
        RECT -12.405 -5.605 -12.075 -5.275 ;
        RECT -12.405 -8.325 -12.075 -7.995 ;
        RECT -12.405 -9.685 -12.075 -9.355 ;
        RECT -12.405 -12.405 -12.075 -12.075 ;
        RECT -12.4 -13.08 -12.08 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -12.405 -27.365 -12.075 -27.035 ;
        RECT -12.405 -28.725 -12.075 -28.395 ;
        RECT -12.405 -30.085 -12.075 -29.755 ;
        RECT -12.405 -31.445 -12.075 -31.115 ;
        RECT -12.405 -32.805 -12.075 -32.475 ;
        RECT -12.405 -36.885 -12.075 -36.555 ;
        RECT -12.405 -37.93 -12.075 -37.6 ;
        RECT -12.405 -40.965 -12.075 -40.635 ;
        RECT -12.405 -42.77 -12.075 -42.44 ;
        RECT -12.405 -43.685 -12.075 -43.355 ;
        RECT -12.405 -51.845 -12.075 -51.515 ;
        RECT -12.405 -53.205 -12.075 -52.875 ;
        RECT -12.405 -54.565 -12.075 -54.235 ;
        RECT -12.405 -55.925 -12.075 -55.595 ;
        RECT -12.405 -57.285 -12.075 -56.955 ;
        RECT -12.405 -58.645 -12.075 -58.315 ;
        RECT -12.405 -60.005 -12.075 -59.675 ;
        RECT -12.405 -61.365 -12.075 -61.035 ;
        RECT -12.405 -62.725 -12.075 -62.395 ;
        RECT -12.405 -64.085 -12.075 -63.755 ;
        RECT -12.405 -65.445 -12.075 -65.115 ;
        RECT -12.405 -66.805 -12.075 -66.475 ;
        RECT -12.405 -68.165 -12.075 -67.835 ;
        RECT -12.405 -69.525 -12.075 -69.195 ;
        RECT -12.405 -70.885 -12.075 -70.555 ;
        RECT -12.405 -72.245 -12.075 -71.915 ;
        RECT -12.405 -74.965 -12.075 -74.635 ;
        RECT -12.405 -76.71 -12.075 -76.38 ;
        RECT -12.405 -77.685 -12.075 -77.355 ;
        RECT -12.405 -79.045 -12.075 -78.715 ;
        RECT -12.405 -81.765 -12.075 -81.435 ;
        RECT -12.405 -83.125 -12.075 -82.795 ;
        RECT -12.405 -84.485 -12.075 -84.155 ;
        RECT -12.405 -85.25 -12.075 -84.92 ;
        RECT -12.405 -87.205 -12.075 -86.875 ;
        RECT -12.405 -89.925 -12.075 -89.595 ;
        RECT -12.405 -91.285 -12.075 -90.955 ;
        RECT -12.405 -92.645 -12.075 -92.315 ;
        RECT -12.405 -94.005 -12.075 -93.675 ;
        RECT -12.405 -96.725 -12.075 -96.395 ;
        RECT -12.405 -98.085 -12.075 -97.755 ;
        RECT -12.405 -98.89 -12.075 -98.56 ;
        RECT -12.405 -100.805 -12.075 -100.475 ;
        RECT -12.405 -102.165 -12.075 -101.835 ;
        RECT -12.405 -104.885 -12.075 -104.555 ;
        RECT -12.405 -106.245 -12.075 -105.915 ;
        RECT -12.405 -107.43 -12.075 -107.1 ;
        RECT -12.405 -113.045 -12.075 -112.715 ;
        RECT -12.405 -114.405 -12.075 -114.075 ;
        RECT -12.405 -115.765 -12.075 -115.435 ;
        RECT -12.405 -117.125 -12.075 -116.795 ;
        RECT -12.405 -119.845 -12.075 -119.515 ;
        RECT -12.405 -125.285 -12.075 -124.955 ;
        RECT -12.405 -129.365 -12.075 -129.035 ;
        RECT -12.405 -133.445 -12.075 -133.115 ;
        RECT -12.405 -136.165 -12.075 -135.835 ;
        RECT -12.405 -137.525 -12.075 -137.195 ;
        RECT -12.405 -138.885 -12.075 -138.555 ;
        RECT -12.405 -140.245 -12.075 -139.915 ;
        RECT -12.405 -141.605 -12.075 -141.275 ;
        RECT -12.405 -145.685 -12.075 -145.355 ;
        RECT -12.405 -147.045 -12.075 -146.715 ;
        RECT -12.405 -148.405 -12.075 -148.075 ;
        RECT -12.405 -149.765 -12.075 -149.435 ;
        RECT -12.405 -152.485 -12.075 -152.155 ;
        RECT -12.405 -153.845 -12.075 -153.515 ;
        RECT -12.405 -155.205 -12.075 -154.875 ;
        RECT -12.405 -156.565 -12.075 -156.235 ;
        RECT -12.405 -159.285 -12.075 -158.955 ;
        RECT -12.405 -160.645 -12.075 -160.315 ;
        RECT -12.405 -162.005 -12.075 -161.675 ;
        RECT -12.405 -163.365 -12.075 -163.035 ;
        RECT -12.405 -164.725 -12.075 -164.395 ;
        RECT -12.405 -166.085 -12.075 -165.755 ;
        RECT -12.405 -170.165 -12.075 -169.835 ;
        RECT -12.405 -172.885 -12.075 -172.555 ;
        RECT -12.405 -174.245 -12.075 -173.915 ;
        RECT -12.405 -175.725 -12.075 -175.395 ;
        RECT -12.405 -176.965 -12.075 -176.635 ;
        RECT -12.405 -178.325 -12.075 -177.995 ;
        RECT -12.405 -180.57 -12.075 -179.44 ;
        RECT -12.4 -180.685 -12.08 -26.36 ;
    END
    PORT
      LAYER met3 ;
        RECT -11.045 241.32 -10.715 242.45 ;
        RECT -11.045 239.195 -10.715 239.525 ;
        RECT -11.045 237.835 -10.715 238.165 ;
        RECT -11.045 236.475 -10.715 236.805 ;
        RECT -11.045 235.115 -10.715 235.445 ;
        RECT -11.045 233.755 -10.715 234.085 ;
        RECT -11.045 232.395 -10.715 232.725 ;
        RECT -11.045 231.035 -10.715 231.365 ;
        RECT -11.045 221.515 -10.715 221.845 ;
        RECT -11.045 217.435 -10.715 217.765 ;
        RECT -11.045 213.355 -10.715 213.685 ;
        RECT -11.045 210.635 -10.715 210.965 ;
        RECT -11.045 203.835 -10.715 204.165 ;
        RECT -11.045 202.475 -10.715 202.805 ;
        RECT -11.045 199.755 -10.715 200.085 ;
        RECT -11.045 192.955 -10.715 193.285 ;
        RECT -11.045 190.235 -10.715 190.565 ;
        RECT -11.045 188.875 -10.715 189.205 ;
        RECT -11.045 184.795 -10.715 185.125 ;
        RECT -11.045 182.075 -10.715 182.405 ;
        RECT -11.045 175.275 -10.715 175.605 ;
        RECT -11.045 173.915 -10.715 174.245 ;
        RECT -11.045 171.195 -10.715 171.525 ;
        RECT -11.045 164.395 -10.715 164.725 ;
        RECT -11.045 161.675 -10.715 162.005 ;
        RECT -11.045 160.315 -10.715 160.645 ;
        RECT -11.045 153.515 -10.715 153.845 ;
        RECT -11.045 150.795 -10.715 151.125 ;
        RECT -11.045 146.715 -10.715 147.045 ;
        RECT -11.045 145.355 -10.715 145.685 ;
        RECT -11.045 142.635 -10.715 142.965 ;
        RECT -11.045 135.835 -10.715 136.165 ;
        RECT -11.045 133.115 -10.715 133.445 ;
        RECT -11.045 131.755 -10.715 132.085 ;
        RECT -11.045 124.955 -10.715 125.285 ;
        RECT -11.045 122.235 -10.715 122.565 ;
        RECT -11.045 118.155 -10.715 118.485 ;
        RECT -11.045 114.075 -10.715 114.405 ;
        RECT -11.045 104.555 -10.715 104.885 ;
        RECT -11.045 103.195 -10.715 103.525 ;
        RECT -11.045 96.395 -10.715 96.725 ;
        RECT -11.045 93.675 -10.715 94.005 ;
        RECT -11.045 89.595 -10.715 89.925 ;
        RECT -11.045 85.515 -10.715 85.845 ;
        RECT -11.045 82.795 -10.715 83.125 ;
        RECT -11.045 75.995 -10.715 76.325 ;
        RECT -11.045 74.635 -10.715 74.965 ;
        RECT -11.045 65.115 -10.715 65.445 ;
        RECT -11.045 61.035 -10.715 61.365 ;
        RECT -11.045 56.955 -10.715 57.285 ;
        RECT -11.045 54.235 -10.715 54.565 ;
        RECT -11.045 47.435 -10.715 47.765 ;
        RECT -11.045 46.075 -10.715 46.405 ;
        RECT -11.045 43.355 -10.715 43.685 ;
        RECT -11.045 36.555 -10.715 36.885 ;
        RECT -11.045 33.835 -10.715 34.165 ;
        RECT -11.045 32.475 -10.715 32.805 ;
        RECT -11.045 28.395 -10.715 28.725 ;
        RECT -11.045 25.675 -10.715 26.005 ;
        RECT -11.045 18.875 -10.715 19.205 ;
        RECT -11.045 17.515 -10.715 17.845 ;
        RECT -11.045 14.795 -10.715 15.125 ;
        RECT -11.045 7.995 -10.715 8.325 ;
        RECT -11.045 5.275 -10.715 5.605 ;
        RECT -11.045 3.915 -10.715 4.245 ;
        RECT -11.045 2.555 -10.715 2.885 ;
        RECT -11.045 1.195 -10.715 1.525 ;
        RECT -11.045 -0.165 -10.715 0.165 ;
        RECT -11.045 -2.885 -10.715 -2.555 ;
        RECT -11.045 -4.245 -10.715 -3.915 ;
        RECT -11.045 -5.605 -10.715 -5.275 ;
        RECT -11.045 -6.965 -10.715 -6.635 ;
        RECT -11.045 -8.325 -10.715 -7.995 ;
        RECT -11.045 -9.685 -10.715 -9.355 ;
        RECT -11.045 -12.405 -10.715 -12.075 ;
        RECT -11.045 -13.765 -10.715 -13.435 ;
        RECT -11.045 -14.95 -10.715 -14.62 ;
        RECT -11.045 -17.845 -10.715 -17.515 ;
        RECT -11.045 -19.79 -10.715 -19.46 ;
        RECT -11.045 -26.005 -10.715 -25.675 ;
        RECT -11.045 -27.365 -10.715 -27.035 ;
        RECT -11.045 -28.725 -10.715 -28.395 ;
        RECT -11.045 -30.085 -10.715 -29.755 ;
        RECT -11.045 -31.445 -10.715 -31.115 ;
        RECT -11.045 -32.805 -10.715 -32.475 ;
        RECT -11.045 -36.885 -10.715 -36.555 ;
        RECT -11.045 -37.93 -10.715 -37.6 ;
        RECT -11.045 -40.965 -10.715 -40.635 ;
        RECT -11.045 -42.77 -10.715 -42.44 ;
        RECT -11.045 -43.685 -10.715 -43.355 ;
        RECT -11.045 -51.845 -10.715 -51.515 ;
        RECT -11.045 -53.205 -10.715 -52.875 ;
        RECT -11.045 -54.565 -10.715 -54.235 ;
        RECT -11.045 -55.925 -10.715 -55.595 ;
        RECT -11.045 -57.285 -10.715 -56.955 ;
        RECT -11.045 -58.645 -10.715 -58.315 ;
        RECT -11.045 -60.005 -10.715 -59.675 ;
        RECT -11.045 -61.365 -10.715 -61.035 ;
        RECT -11.045 -62.725 -10.715 -62.395 ;
        RECT -11.045 -64.085 -10.715 -63.755 ;
        RECT -11.045 -65.445 -10.715 -65.115 ;
        RECT -11.045 -66.805 -10.715 -66.475 ;
        RECT -11.045 -68.165 -10.715 -67.835 ;
        RECT -11.045 -69.525 -10.715 -69.195 ;
        RECT -11.045 -70.885 -10.715 -70.555 ;
        RECT -11.045 -72.245 -10.715 -71.915 ;
        RECT -11.045 -74.965 -10.715 -74.635 ;
        RECT -11.045 -76.71 -10.715 -76.38 ;
        RECT -11.045 -77.685 -10.715 -77.355 ;
        RECT -11.045 -79.045 -10.715 -78.715 ;
        RECT -11.045 -81.765 -10.715 -81.435 ;
        RECT -11.045 -83.125 -10.715 -82.795 ;
        RECT -11.045 -84.485 -10.715 -84.155 ;
        RECT -11.045 -85.25 -10.715 -84.92 ;
        RECT -11.045 -87.205 -10.715 -86.875 ;
        RECT -11.045 -89.925 -10.715 -89.595 ;
        RECT -11.045 -91.285 -10.715 -90.955 ;
        RECT -11.045 -92.645 -10.715 -92.315 ;
        RECT -11.045 -94.005 -10.715 -93.675 ;
        RECT -11.045 -96.725 -10.715 -96.395 ;
        RECT -11.045 -98.085 -10.715 -97.755 ;
        RECT -11.045 -98.89 -10.715 -98.56 ;
        RECT -11.045 -100.805 -10.715 -100.475 ;
        RECT -11.045 -102.165 -10.715 -101.835 ;
        RECT -11.045 -104.885 -10.715 -104.555 ;
        RECT -11.045 -106.245 -10.715 -105.915 ;
        RECT -11.045 -107.43 -10.715 -107.1 ;
        RECT -11.045 -113.045 -10.715 -112.715 ;
        RECT -11.045 -114.405 -10.715 -114.075 ;
        RECT -11.045 -115.765 -10.715 -115.435 ;
        RECT -11.045 -117.125 -10.715 -116.795 ;
        RECT -11.045 -119.845 -10.715 -119.515 ;
        RECT -11.045 -125.285 -10.715 -124.955 ;
        RECT -11.045 -126.645 -10.715 -126.315 ;
        RECT -11.045 -129.365 -10.715 -129.035 ;
        RECT -11.045 -130.725 -10.715 -130.395 ;
        RECT -11.045 -133.445 -10.715 -133.115 ;
        RECT -11.045 -134.805 -10.715 -134.475 ;
        RECT -11.045 -136.165 -10.715 -135.835 ;
        RECT -11.045 -137.525 -10.715 -137.195 ;
        RECT -11.045 -138.885 -10.715 -138.555 ;
        RECT -11.045 -140.245 -10.715 -139.915 ;
        RECT -11.045 -141.605 -10.715 -141.275 ;
        RECT -11.045 -145.685 -10.715 -145.355 ;
        RECT -11.045 -147.045 -10.715 -146.715 ;
        RECT -11.045 -148.405 -10.715 -148.075 ;
        RECT -11.045 -149.765 -10.715 -149.435 ;
        RECT -11.045 -151.125 -10.715 -150.795 ;
        RECT -11.045 -152.485 -10.715 -152.155 ;
        RECT -11.045 -153.845 -10.715 -153.515 ;
        RECT -11.045 -155.205 -10.715 -154.875 ;
        RECT -11.045 -156.565 -10.715 -156.235 ;
        RECT -11.045 -159.285 -10.715 -158.955 ;
        RECT -11.045 -160.645 -10.715 -160.315 ;
        RECT -11.045 -162.005 -10.715 -161.675 ;
        RECT -11.045 -163.365 -10.715 -163.035 ;
        RECT -11.045 -164.725 -10.715 -164.395 ;
        RECT -11.045 -166.085 -10.715 -165.755 ;
        RECT -11.045 -170.165 -10.715 -169.835 ;
        RECT -11.045 -174.245 -10.715 -173.915 ;
        RECT -11.045 -175.725 -10.715 -175.395 ;
        RECT -11.045 -176.965 -10.715 -176.635 ;
        RECT -11.045 -178.325 -10.715 -177.995 ;
        RECT -11.045 -180.57 -10.715 -179.44 ;
        RECT -11.04 -180.685 -10.72 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -9.685 241.32 -9.355 242.45 ;
        RECT -9.685 239.195 -9.355 239.525 ;
        RECT -9.685 237.835 -9.355 238.165 ;
        RECT -9.685 236.475 -9.355 236.805 ;
        RECT -9.685 235.115 -9.355 235.445 ;
        RECT -9.685 233.755 -9.355 234.085 ;
        RECT -9.685 232.395 -9.355 232.725 ;
        RECT -9.685 231.035 -9.355 231.365 ;
        RECT -9.685 221.515 -9.355 221.845 ;
        RECT -9.685 217.435 -9.355 217.765 ;
        RECT -9.685 213.355 -9.355 213.685 ;
        RECT -9.685 210.635 -9.355 210.965 ;
        RECT -9.685 203.835 -9.355 204.165 ;
        RECT -9.685 202.475 -9.355 202.805 ;
        RECT -9.685 199.755 -9.355 200.085 ;
        RECT -9.685 192.955 -9.355 193.285 ;
        RECT -9.685 190.235 -9.355 190.565 ;
        RECT -9.685 188.875 -9.355 189.205 ;
        RECT -9.685 184.795 -9.355 185.125 ;
        RECT -9.685 182.075 -9.355 182.405 ;
        RECT -9.685 175.275 -9.355 175.605 ;
        RECT -9.685 173.915 -9.355 174.245 ;
        RECT -9.685 171.195 -9.355 171.525 ;
        RECT -9.685 164.395 -9.355 164.725 ;
        RECT -9.685 161.675 -9.355 162.005 ;
        RECT -9.685 160.315 -9.355 160.645 ;
        RECT -9.685 153.515 -9.355 153.845 ;
        RECT -9.685 150.795 -9.355 151.125 ;
        RECT -9.685 146.715 -9.355 147.045 ;
        RECT -9.685 145.355 -9.355 145.685 ;
        RECT -9.685 142.635 -9.355 142.965 ;
        RECT -9.685 135.835 -9.355 136.165 ;
        RECT -9.685 133.115 -9.355 133.445 ;
        RECT -9.685 131.755 -9.355 132.085 ;
        RECT -9.685 124.955 -9.355 125.285 ;
        RECT -9.685 122.235 -9.355 122.565 ;
        RECT -9.685 118.155 -9.355 118.485 ;
        RECT -9.685 114.075 -9.355 114.405 ;
        RECT -9.685 104.555 -9.355 104.885 ;
        RECT -9.685 103.195 -9.355 103.525 ;
        RECT -9.685 96.395 -9.355 96.725 ;
        RECT -9.685 93.675 -9.355 94.005 ;
        RECT -9.685 89.595 -9.355 89.925 ;
        RECT -9.685 85.515 -9.355 85.845 ;
        RECT -9.685 82.795 -9.355 83.125 ;
        RECT -9.685 75.995 -9.355 76.325 ;
        RECT -9.685 74.635 -9.355 74.965 ;
        RECT -9.685 65.115 -9.355 65.445 ;
        RECT -9.685 61.035 -9.355 61.365 ;
        RECT -9.685 56.955 -9.355 57.285 ;
        RECT -9.685 54.235 -9.355 54.565 ;
        RECT -9.685 47.435 -9.355 47.765 ;
        RECT -9.685 46.075 -9.355 46.405 ;
        RECT -9.685 43.355 -9.355 43.685 ;
        RECT -9.685 36.555 -9.355 36.885 ;
        RECT -9.685 33.835 -9.355 34.165 ;
        RECT -9.685 32.475 -9.355 32.805 ;
        RECT -9.685 28.395 -9.355 28.725 ;
        RECT -9.685 25.675 -9.355 26.005 ;
        RECT -9.685 18.875 -9.355 19.205 ;
        RECT -9.685 17.515 -9.355 17.845 ;
        RECT -9.685 14.795 -9.355 15.125 ;
        RECT -9.685 7.995 -9.355 8.325 ;
        RECT -9.685 5.275 -9.355 5.605 ;
        RECT -9.685 3.915 -9.355 4.245 ;
        RECT -9.685 2.555 -9.355 2.885 ;
        RECT -9.685 1.195 -9.355 1.525 ;
        RECT -9.685 -0.165 -9.355 0.165 ;
        RECT -9.685 -2.885 -9.355 -2.555 ;
        RECT -9.685 -4.245 -9.355 -3.915 ;
        RECT -9.685 -5.605 -9.355 -5.275 ;
        RECT -9.685 -6.965 -9.355 -6.635 ;
        RECT -9.685 -8.325 -9.355 -7.995 ;
        RECT -9.685 -9.685 -9.355 -9.355 ;
        RECT -9.685 -12.405 -9.355 -12.075 ;
        RECT -9.685 -13.765 -9.355 -13.435 ;
        RECT -9.685 -17.845 -9.355 -17.515 ;
        RECT -9.685 -26.005 -9.355 -25.675 ;
        RECT -9.685 -27.365 -9.355 -27.035 ;
        RECT -9.685 -28.725 -9.355 -28.395 ;
        RECT -9.685 -30.085 -9.355 -29.755 ;
        RECT -9.685 -31.445 -9.355 -31.115 ;
        RECT -9.685 -32.805 -9.355 -32.475 ;
        RECT -9.685 -36.885 -9.355 -36.555 ;
        RECT -9.685 -40.965 -9.355 -40.635 ;
        RECT -9.685 -43.685 -9.355 -43.355 ;
        RECT -9.685 -51.845 -9.355 -51.515 ;
        RECT -9.685 -53.205 -9.355 -52.875 ;
        RECT -9.685 -54.565 -9.355 -54.235 ;
        RECT -9.685 -55.925 -9.355 -55.595 ;
        RECT -9.685 -57.285 -9.355 -56.955 ;
        RECT -9.685 -58.645 -9.355 -58.315 ;
        RECT -9.685 -60.005 -9.355 -59.675 ;
        RECT -9.685 -61.365 -9.355 -61.035 ;
        RECT -9.685 -62.725 -9.355 -62.395 ;
        RECT -9.685 -64.085 -9.355 -63.755 ;
        RECT -9.685 -65.445 -9.355 -65.115 ;
        RECT -9.685 -66.805 -9.355 -66.475 ;
        RECT -9.685 -68.165 -9.355 -67.835 ;
        RECT -9.685 -69.525 -9.355 -69.195 ;
        RECT -9.685 -70.885 -9.355 -70.555 ;
        RECT -9.685 -72.245 -9.355 -71.915 ;
        RECT -9.685 -74.965 -9.355 -74.635 ;
        RECT -9.685 -77.685 -9.355 -77.355 ;
        RECT -9.685 -79.045 -9.355 -78.715 ;
        RECT -9.685 -81.765 -9.355 -81.435 ;
        RECT -9.685 -83.125 -9.355 -82.795 ;
        RECT -9.685 -84.485 -9.355 -84.155 ;
        RECT -9.68 -85.84 -9.36 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -8.325 241.32 -7.995 242.45 ;
        RECT -8.325 239.195 -7.995 239.525 ;
        RECT -8.325 237.835 -7.995 238.165 ;
        RECT -8.325 236.475 -7.995 236.805 ;
        RECT -8.325 235.115 -7.995 235.445 ;
        RECT -8.325 233.755 -7.995 234.085 ;
        RECT -8.325 232.395 -7.995 232.725 ;
        RECT -8.325 231.035 -7.995 231.365 ;
        RECT -8.325 221.515 -7.995 221.845 ;
        RECT -8.325 217.435 -7.995 217.765 ;
        RECT -8.325 213.355 -7.995 213.685 ;
        RECT -8.325 210.635 -7.995 210.965 ;
        RECT -8.325 203.835 -7.995 204.165 ;
        RECT -8.325 202.475 -7.995 202.805 ;
        RECT -8.325 199.755 -7.995 200.085 ;
        RECT -8.325 192.955 -7.995 193.285 ;
        RECT -8.325 190.235 -7.995 190.565 ;
        RECT -8.325 188.875 -7.995 189.205 ;
        RECT -8.325 184.795 -7.995 185.125 ;
        RECT -8.325 182.075 -7.995 182.405 ;
        RECT -8.325 175.275 -7.995 175.605 ;
        RECT -8.325 173.915 -7.995 174.245 ;
        RECT -8.325 171.195 -7.995 171.525 ;
        RECT -8.325 164.395 -7.995 164.725 ;
        RECT -8.325 161.675 -7.995 162.005 ;
        RECT -8.325 160.315 -7.995 160.645 ;
        RECT -8.325 153.515 -7.995 153.845 ;
        RECT -8.325 150.795 -7.995 151.125 ;
        RECT -8.325 146.715 -7.995 147.045 ;
        RECT -8.325 145.355 -7.995 145.685 ;
        RECT -8.325 142.635 -7.995 142.965 ;
        RECT -8.325 135.835 -7.995 136.165 ;
        RECT -8.325 133.115 -7.995 133.445 ;
        RECT -8.325 131.755 -7.995 132.085 ;
        RECT -8.325 124.955 -7.995 125.285 ;
        RECT -8.325 122.235 -7.995 122.565 ;
        RECT -8.325 118.155 -7.995 118.485 ;
        RECT -8.325 114.075 -7.995 114.405 ;
        RECT -8.325 104.555 -7.995 104.885 ;
        RECT -8.325 103.195 -7.995 103.525 ;
        RECT -8.325 96.395 -7.995 96.725 ;
        RECT -8.325 93.675 -7.995 94.005 ;
        RECT -8.325 89.595 -7.995 89.925 ;
        RECT -8.325 85.515 -7.995 85.845 ;
        RECT -8.325 82.795 -7.995 83.125 ;
        RECT -8.325 75.995 -7.995 76.325 ;
        RECT -8.325 74.635 -7.995 74.965 ;
        RECT -8.325 65.115 -7.995 65.445 ;
        RECT -8.325 61.035 -7.995 61.365 ;
        RECT -8.325 56.955 -7.995 57.285 ;
        RECT -8.325 54.235 -7.995 54.565 ;
        RECT -8.325 47.435 -7.995 47.765 ;
        RECT -8.325 46.075 -7.995 46.405 ;
        RECT -8.325 43.355 -7.995 43.685 ;
        RECT -8.325 36.555 -7.995 36.885 ;
        RECT -8.325 33.835 -7.995 34.165 ;
        RECT -8.325 32.475 -7.995 32.805 ;
        RECT -8.325 28.395 -7.995 28.725 ;
        RECT -8.325 25.675 -7.995 26.005 ;
        RECT -8.325 18.875 -7.995 19.205 ;
        RECT -8.325 17.515 -7.995 17.845 ;
        RECT -8.325 14.795 -7.995 15.125 ;
        RECT -8.325 7.995 -7.995 8.325 ;
        RECT -8.325 5.275 -7.995 5.605 ;
        RECT -8.325 3.915 -7.995 4.245 ;
        RECT -8.325 2.555 -7.995 2.885 ;
        RECT -8.325 1.195 -7.995 1.525 ;
        RECT -8.325 -0.165 -7.995 0.165 ;
        RECT -8.32 -0.84 -8 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -8.325 -122.565 -7.995 -122.235 ;
        RECT -8.325 -123.925 -7.995 -123.595 ;
        RECT -8.325 -125.285 -7.995 -124.955 ;
        RECT -8.325 -126.645 -7.995 -126.315 ;
        RECT -8.325 -128.005 -7.995 -127.675 ;
        RECT -8.325 -129.365 -7.995 -129.035 ;
        RECT -8.325 -130.725 -7.995 -130.395 ;
        RECT -8.325 -132.085 -7.995 -131.755 ;
        RECT -8.325 -133.445 -7.995 -133.115 ;
        RECT -8.325 -134.805 -7.995 -134.475 ;
        RECT -8.325 -136.165 -7.995 -135.835 ;
        RECT -8.325 -137.525 -7.995 -137.195 ;
        RECT -8.325 -138.885 -7.995 -138.555 ;
        RECT -8.325 -140.245 -7.995 -139.915 ;
        RECT -8.325 -141.605 -7.995 -141.275 ;
        RECT -8.325 -142.965 -7.995 -142.635 ;
        RECT -8.325 -144.325 -7.995 -143.995 ;
        RECT -8.325 -145.685 -7.995 -145.355 ;
        RECT -8.325 -147.045 -7.995 -146.715 ;
        RECT -8.325 -148.405 -7.995 -148.075 ;
        RECT -8.325 -149.765 -7.995 -149.435 ;
        RECT -8.325 -151.125 -7.995 -150.795 ;
        RECT -8.325 -152.485 -7.995 -152.155 ;
        RECT -8.325 -153.845 -7.995 -153.515 ;
        RECT -8.325 -155.205 -7.995 -154.875 ;
        RECT -8.325 -156.565 -7.995 -156.235 ;
        RECT -8.325 -157.925 -7.995 -157.595 ;
        RECT -8.325 -159.285 -7.995 -158.955 ;
        RECT -8.325 -160.645 -7.995 -160.315 ;
        RECT -8.325 -162.005 -7.995 -161.675 ;
        RECT -8.325 -163.365 -7.995 -163.035 ;
        RECT -8.325 -164.725 -7.995 -164.395 ;
        RECT -8.325 -166.085 -7.995 -165.755 ;
        RECT -8.325 -167.445 -7.995 -167.115 ;
        RECT -8.325 -168.805 -7.995 -168.475 ;
        RECT -8.325 -170.165 -7.995 -169.835 ;
        RECT -8.325 -171.525 -7.995 -171.195 ;
        RECT -8.325 -172.885 -7.995 -172.555 ;
        RECT -8.325 -174.245 -7.995 -173.915 ;
        RECT -8.325 -175.605 -7.995 -175.275 ;
        RECT -8.325 -176.965 -7.995 -176.635 ;
        RECT -8.325 -178.325 -7.995 -177.995 ;
        RECT -8.325 -180.57 -7.995 -179.44 ;
        RECT -8.32 -180.685 -8 -121.56 ;
    END
    PORT
      LAYER met3 ;
        RECT -6.965 241.32 -6.635 242.45 ;
        RECT -6.965 239.195 -6.635 239.525 ;
        RECT -6.965 237.835 -6.635 238.165 ;
        RECT -6.965 236.475 -6.635 236.805 ;
        RECT -6.965 235.115 -6.635 235.445 ;
        RECT -6.965 233.755 -6.635 234.085 ;
        RECT -6.965 232.395 -6.635 232.725 ;
        RECT -6.965 231.035 -6.635 231.365 ;
        RECT -6.965 221.515 -6.635 221.845 ;
        RECT -6.965 217.435 -6.635 217.765 ;
        RECT -6.965 213.355 -6.635 213.685 ;
        RECT -6.965 210.635 -6.635 210.965 ;
        RECT -6.965 203.835 -6.635 204.165 ;
        RECT -6.965 202.475 -6.635 202.805 ;
        RECT -6.965 199.755 -6.635 200.085 ;
        RECT -6.965 192.955 -6.635 193.285 ;
        RECT -6.965 190.235 -6.635 190.565 ;
        RECT -6.965 188.875 -6.635 189.205 ;
        RECT -6.965 184.795 -6.635 185.125 ;
        RECT -6.965 182.075 -6.635 182.405 ;
        RECT -6.965 175.275 -6.635 175.605 ;
        RECT -6.965 173.915 -6.635 174.245 ;
        RECT -6.965 171.195 -6.635 171.525 ;
        RECT -6.965 164.395 -6.635 164.725 ;
        RECT -6.965 161.675 -6.635 162.005 ;
        RECT -6.965 160.315 -6.635 160.645 ;
        RECT -6.965 153.515 -6.635 153.845 ;
        RECT -6.965 150.795 -6.635 151.125 ;
        RECT -6.965 146.715 -6.635 147.045 ;
        RECT -6.965 145.355 -6.635 145.685 ;
        RECT -6.965 142.635 -6.635 142.965 ;
        RECT -6.965 135.835 -6.635 136.165 ;
        RECT -6.965 133.115 -6.635 133.445 ;
        RECT -6.965 131.755 -6.635 132.085 ;
        RECT -6.965 124.955 -6.635 125.285 ;
        RECT -6.965 122.235 -6.635 122.565 ;
        RECT -6.965 118.155 -6.635 118.485 ;
        RECT -6.965 114.075 -6.635 114.405 ;
        RECT -6.965 104.555 -6.635 104.885 ;
        RECT -6.965 103.195 -6.635 103.525 ;
        RECT -6.965 96.395 -6.635 96.725 ;
        RECT -6.965 93.675 -6.635 94.005 ;
        RECT -6.965 89.595 -6.635 89.925 ;
        RECT -6.965 85.515 -6.635 85.845 ;
        RECT -6.965 82.795 -6.635 83.125 ;
        RECT -6.965 75.995 -6.635 76.325 ;
        RECT -6.965 74.635 -6.635 74.965 ;
        RECT -6.965 65.115 -6.635 65.445 ;
        RECT -6.965 61.035 -6.635 61.365 ;
        RECT -6.965 56.955 -6.635 57.285 ;
        RECT -6.965 54.235 -6.635 54.565 ;
        RECT -6.965 47.435 -6.635 47.765 ;
        RECT -6.965 46.075 -6.635 46.405 ;
        RECT -6.965 43.355 -6.635 43.685 ;
        RECT -6.965 36.555 -6.635 36.885 ;
        RECT -6.965 33.835 -6.635 34.165 ;
        RECT -6.965 32.475 -6.635 32.805 ;
        RECT -6.965 28.395 -6.635 28.725 ;
        RECT -6.965 25.675 -6.635 26.005 ;
        RECT -6.965 18.875 -6.635 19.205 ;
        RECT -6.965 17.515 -6.635 17.845 ;
        RECT -6.965 14.795 -6.635 15.125 ;
        RECT -6.965 7.995 -6.635 8.325 ;
        RECT -6.965 5.275 -6.635 5.605 ;
        RECT -6.965 3.915 -6.635 4.245 ;
        RECT -6.965 2.555 -6.635 2.885 ;
        RECT -6.965 1.195 -6.635 1.525 ;
        RECT -6.965 -0.165 -6.635 0.165 ;
        RECT -6.965 -1.525 -6.635 -1.195 ;
        RECT -6.965 -2.885 -6.635 -2.555 ;
        RECT -6.965 -4.245 -6.635 -3.915 ;
        RECT -6.965 -5.605 -6.635 -5.275 ;
        RECT -6.965 -6.965 -6.635 -6.635 ;
        RECT -6.965 -8.325 -6.635 -7.995 ;
        RECT -6.965 -9.685 -6.635 -9.355 ;
        RECT -6.965 -12.405 -6.635 -12.075 ;
        RECT -6.965 -13.765 -6.635 -13.435 ;
        RECT -6.965 -15.125 -6.635 -14.795 ;
        RECT -6.965 -16.485 -6.635 -16.155 ;
        RECT -6.965 -17.845 -6.635 -17.515 ;
        RECT -6.965 -21.925 -6.635 -21.595 ;
        RECT -6.965 -23.285 -6.635 -22.955 ;
        RECT -6.965 -24.645 -6.635 -24.315 ;
        RECT -6.965 -26.005 -6.635 -25.675 ;
        RECT -6.965 -27.365 -6.635 -27.035 ;
        RECT -6.965 -28.725 -6.635 -28.395 ;
        RECT -6.965 -30.085 -6.635 -29.755 ;
        RECT -6.965 -31.445 -6.635 -31.115 ;
        RECT -6.965 -32.805 -6.635 -32.475 ;
        RECT -6.965 -34.165 -6.635 -33.835 ;
        RECT -6.965 -36.885 -6.635 -36.555 ;
        RECT -6.965 -38.245 -6.635 -37.915 ;
        RECT -6.965 -40.965 -6.635 -40.635 ;
        RECT -6.965 -42.325 -6.635 -41.995 ;
        RECT -6.965 -43.685 -6.635 -43.355 ;
        RECT -6.965 -45.045 -6.635 -44.715 ;
        RECT -6.965 -46.405 -6.635 -46.075 ;
        RECT -6.965 -47.765 -6.635 -47.435 ;
        RECT -6.965 -49.125 -6.635 -48.795 ;
        RECT -6.965 -51.845 -6.635 -51.515 ;
        RECT -6.965 -53.205 -6.635 -52.875 ;
        RECT -6.965 -54.565 -6.635 -54.235 ;
        RECT -6.965 -55.925 -6.635 -55.595 ;
        RECT -6.965 -57.285 -6.635 -56.955 ;
        RECT -6.965 -58.645 -6.635 -58.315 ;
        RECT -6.965 -60.005 -6.635 -59.675 ;
        RECT -6.965 -61.365 -6.635 -61.035 ;
        RECT -6.965 -62.725 -6.635 -62.395 ;
        RECT -6.965 -64.085 -6.635 -63.755 ;
        RECT -6.965 -65.445 -6.635 -65.115 ;
        RECT -6.965 -66.805 -6.635 -66.475 ;
        RECT -6.965 -68.165 -6.635 -67.835 ;
        RECT -6.965 -69.525 -6.635 -69.195 ;
        RECT -6.965 -70.885 -6.635 -70.555 ;
        RECT -6.965 -72.245 -6.635 -71.915 ;
        RECT -6.965 -73.605 -6.635 -73.275 ;
        RECT -6.965 -74.965 -6.635 -74.635 ;
        RECT -6.965 -76.325 -6.635 -75.995 ;
        RECT -6.965 -77.685 -6.635 -77.355 ;
        RECT -6.965 -79.045 -6.635 -78.715 ;
        RECT -6.965 -80.405 -6.635 -80.075 ;
        RECT -6.965 -81.765 -6.635 -81.435 ;
        RECT -6.965 -83.125 -6.635 -82.795 ;
        RECT -6.965 -84.485 -6.635 -84.155 ;
        RECT -6.965 -85.845 -6.635 -85.515 ;
        RECT -6.965 -87.205 -6.635 -86.875 ;
        RECT -6.965 -88.565 -6.635 -88.235 ;
        RECT -6.965 -89.925 -6.635 -89.595 ;
        RECT -6.965 -91.285 -6.635 -90.955 ;
        RECT -6.965 -92.645 -6.635 -92.315 ;
        RECT -6.965 -94.005 -6.635 -93.675 ;
        RECT -6.965 -95.365 -6.635 -95.035 ;
        RECT -6.965 -96.725 -6.635 -96.395 ;
        RECT -6.965 -98.085 -6.635 -97.755 ;
        RECT -6.965 -99.445 -6.635 -99.115 ;
        RECT -6.965 -100.805 -6.635 -100.475 ;
        RECT -6.965 -102.165 -6.635 -101.835 ;
        RECT -6.965 -103.525 -6.635 -103.195 ;
        RECT -6.965 -104.885 -6.635 -104.555 ;
        RECT -6.965 -106.245 -6.635 -105.915 ;
        RECT -6.965 -107.605 -6.635 -107.275 ;
        RECT -6.965 -108.965 -6.635 -108.635 ;
        RECT -6.965 -110.325 -6.635 -109.995 ;
        RECT -6.965 -111.685 -6.635 -111.355 ;
        RECT -6.965 -113.045 -6.635 -112.715 ;
        RECT -6.965 -114.405 -6.635 -114.075 ;
        RECT -6.965 -115.765 -6.635 -115.435 ;
        RECT -6.965 -117.125 -6.635 -116.795 ;
        RECT -6.965 -119.845 -6.635 -119.515 ;
        RECT -6.965 -121.205 -6.635 -120.875 ;
        RECT -6.965 -122.565 -6.635 -122.235 ;
        RECT -6.965 -123.925 -6.635 -123.595 ;
        RECT -6.965 -125.285 -6.635 -124.955 ;
        RECT -6.965 -126.645 -6.635 -126.315 ;
        RECT -6.965 -128.005 -6.635 -127.675 ;
        RECT -6.965 -129.365 -6.635 -129.035 ;
        RECT -6.965 -130.725 -6.635 -130.395 ;
        RECT -6.965 -132.085 -6.635 -131.755 ;
        RECT -6.965 -133.445 -6.635 -133.115 ;
        RECT -6.965 -134.805 -6.635 -134.475 ;
        RECT -6.965 -136.165 -6.635 -135.835 ;
        RECT -6.965 -137.525 -6.635 -137.195 ;
        RECT -6.965 -138.885 -6.635 -138.555 ;
        RECT -6.965 -140.245 -6.635 -139.915 ;
        RECT -6.965 -141.605 -6.635 -141.275 ;
        RECT -6.965 -142.965 -6.635 -142.635 ;
        RECT -6.965 -144.325 -6.635 -143.995 ;
        RECT -6.965 -145.685 -6.635 -145.355 ;
        RECT -6.965 -147.045 -6.635 -146.715 ;
        RECT -6.965 -148.405 -6.635 -148.075 ;
        RECT -6.965 -149.765 -6.635 -149.435 ;
        RECT -6.965 -151.125 -6.635 -150.795 ;
        RECT -6.965 -152.485 -6.635 -152.155 ;
        RECT -6.965 -153.845 -6.635 -153.515 ;
        RECT -6.965 -155.205 -6.635 -154.875 ;
        RECT -6.965 -156.565 -6.635 -156.235 ;
        RECT -6.965 -157.925 -6.635 -157.595 ;
        RECT -6.965 -159.285 -6.635 -158.955 ;
        RECT -6.965 -160.645 -6.635 -160.315 ;
        RECT -6.965 -162.005 -6.635 -161.675 ;
        RECT -6.965 -163.365 -6.635 -163.035 ;
        RECT -6.965 -164.725 -6.635 -164.395 ;
        RECT -6.965 -166.085 -6.635 -165.755 ;
        RECT -6.965 -167.445 -6.635 -167.115 ;
        RECT -6.965 -168.805 -6.635 -168.475 ;
        RECT -6.965 -170.165 -6.635 -169.835 ;
        RECT -6.965 -171.525 -6.635 -171.195 ;
        RECT -6.965 -172.885 -6.635 -172.555 ;
        RECT -6.965 -174.245 -6.635 -173.915 ;
        RECT -6.965 -175.605 -6.635 -175.275 ;
        RECT -6.965 -176.965 -6.635 -176.635 ;
        RECT -6.965 -178.325 -6.635 -177.995 ;
        RECT -6.965 -180.57 -6.635 -179.44 ;
        RECT -6.96 -180.685 -6.64 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -5.605 -108.965 -5.275 -108.635 ;
        RECT -5.605 -110.325 -5.275 -109.995 ;
        RECT -5.605 -111.685 -5.275 -111.355 ;
        RECT -5.605 -113.045 -5.275 -112.715 ;
        RECT -5.605 -114.405 -5.275 -114.075 ;
        RECT -5.605 -115.765 -5.275 -115.435 ;
        RECT -5.605 -117.125 -5.275 -116.795 ;
        RECT -5.605 -119.845 -5.275 -119.515 ;
        RECT -5.605 -121.205 -5.275 -120.875 ;
        RECT -5.605 -122.565 -5.275 -122.235 ;
        RECT -5.605 -123.925 -5.275 -123.595 ;
        RECT -5.605 -125.285 -5.275 -124.955 ;
        RECT -5.605 -126.645 -5.275 -126.315 ;
        RECT -5.605 -128.005 -5.275 -127.675 ;
        RECT -5.605 -129.365 -5.275 -129.035 ;
        RECT -5.605 -130.725 -5.275 -130.395 ;
        RECT -5.605 -132.085 -5.275 -131.755 ;
        RECT -5.605 -133.445 -5.275 -133.115 ;
        RECT -5.605 -134.805 -5.275 -134.475 ;
        RECT -5.605 -136.165 -5.275 -135.835 ;
        RECT -5.605 -137.525 -5.275 -137.195 ;
        RECT -5.605 -138.885 -5.275 -138.555 ;
        RECT -5.605 -140.245 -5.275 -139.915 ;
        RECT -5.605 -141.605 -5.275 -141.275 ;
        RECT -5.605 -142.965 -5.275 -142.635 ;
        RECT -5.605 -144.325 -5.275 -143.995 ;
        RECT -5.605 -145.685 -5.275 -145.355 ;
        RECT -5.605 -147.045 -5.275 -146.715 ;
        RECT -5.605 -148.405 -5.275 -148.075 ;
        RECT -5.605 -149.765 -5.275 -149.435 ;
        RECT -5.605 -151.125 -5.275 -150.795 ;
        RECT -5.605 -152.485 -5.275 -152.155 ;
        RECT -5.605 -153.845 -5.275 -153.515 ;
        RECT -5.605 -155.205 -5.275 -154.875 ;
        RECT -5.605 -156.565 -5.275 -156.235 ;
        RECT -5.605 -157.925 -5.275 -157.595 ;
        RECT -5.605 -159.285 -5.275 -158.955 ;
        RECT -5.605 -160.645 -5.275 -160.315 ;
        RECT -5.605 -162.005 -5.275 -161.675 ;
        RECT -5.605 -163.365 -5.275 -163.035 ;
        RECT -5.605 -164.725 -5.275 -164.395 ;
        RECT -5.605 -166.085 -5.275 -165.755 ;
        RECT -5.605 -167.445 -5.275 -167.115 ;
        RECT -5.605 -168.805 -5.275 -168.475 ;
        RECT -5.605 -170.165 -5.275 -169.835 ;
        RECT -5.605 -171.525 -5.275 -171.195 ;
        RECT -5.605 -172.885 -5.275 -172.555 ;
        RECT -5.605 -174.245 -5.275 -173.915 ;
        RECT -5.605 -175.605 -5.275 -175.275 ;
        RECT -5.605 -176.965 -5.275 -176.635 ;
        RECT -5.605 -178.325 -5.275 -177.995 ;
        RECT -5.605 -180.57 -5.275 -179.44 ;
        RECT -5.6 -180.685 -5.28 242.565 ;
        RECT -5.605 241.32 -5.275 242.45 ;
        RECT -5.605 239.195 -5.275 239.525 ;
        RECT -5.605 237.835 -5.275 238.165 ;
        RECT -5.605 235.975 -5.275 236.305 ;
        RECT -5.605 233.925 -5.275 234.255 ;
        RECT -5.605 231.995 -5.275 232.325 ;
        RECT -5.605 230.155 -5.275 230.485 ;
        RECT -5.605 228.665 -5.275 228.995 ;
        RECT -5.605 226.995 -5.275 227.325 ;
        RECT -5.605 225.505 -5.275 225.835 ;
        RECT -5.605 223.835 -5.275 224.165 ;
        RECT -5.605 222.345 -5.275 222.675 ;
        RECT -5.605 220.675 -5.275 221.005 ;
        RECT -5.605 219.185 -5.275 219.515 ;
        RECT -5.605 217.775 -5.275 218.105 ;
        RECT -5.605 215.935 -5.275 216.265 ;
        RECT -5.605 214.445 -5.275 214.775 ;
        RECT -5.605 212.775 -5.275 213.105 ;
        RECT -5.605 211.285 -5.275 211.615 ;
        RECT -5.605 209.615 -5.275 209.945 ;
        RECT -5.605 208.125 -5.275 208.455 ;
        RECT -5.605 206.455 -5.275 206.785 ;
        RECT -5.605 204.965 -5.275 205.295 ;
        RECT -5.605 203.555 -5.275 203.885 ;
        RECT -5.605 201.715 -5.275 202.045 ;
        RECT -5.605 200.225 -5.275 200.555 ;
        RECT -5.605 198.555 -5.275 198.885 ;
        RECT -5.605 197.065 -5.275 197.395 ;
        RECT -5.605 195.395 -5.275 195.725 ;
        RECT -5.605 193.905 -5.275 194.235 ;
        RECT -5.605 192.235 -5.275 192.565 ;
        RECT -5.605 190.745 -5.275 191.075 ;
        RECT -5.605 189.335 -5.275 189.665 ;
        RECT -5.605 187.495 -5.275 187.825 ;
        RECT -5.605 186.005 -5.275 186.335 ;
        RECT -5.605 184.335 -5.275 184.665 ;
        RECT -5.605 182.845 -5.275 183.175 ;
        RECT -5.605 181.175 -5.275 181.505 ;
        RECT -5.605 179.685 -5.275 180.015 ;
        RECT -5.605 178.015 -5.275 178.345 ;
        RECT -5.605 176.525 -5.275 176.855 ;
        RECT -5.605 175.115 -5.275 175.445 ;
        RECT -5.605 173.275 -5.275 173.605 ;
        RECT -5.605 171.785 -5.275 172.115 ;
        RECT -5.605 170.115 -5.275 170.445 ;
        RECT -5.605 168.625 -5.275 168.955 ;
        RECT -5.605 166.955 -5.275 167.285 ;
        RECT -5.605 165.465 -5.275 165.795 ;
        RECT -5.605 163.795 -5.275 164.125 ;
        RECT -5.605 162.305 -5.275 162.635 ;
        RECT -5.605 160.895 -5.275 161.225 ;
        RECT -5.605 159.055 -5.275 159.385 ;
        RECT -5.605 157.565 -5.275 157.895 ;
        RECT -5.605 155.895 -5.275 156.225 ;
        RECT -5.605 154.405 -5.275 154.735 ;
        RECT -5.605 152.735 -5.275 153.065 ;
        RECT -5.605 151.245 -5.275 151.575 ;
        RECT -5.605 149.575 -5.275 149.905 ;
        RECT -5.605 148.085 -5.275 148.415 ;
        RECT -5.605 146.675 -5.275 147.005 ;
        RECT -5.605 144.835 -5.275 145.165 ;
        RECT -5.605 143.345 -5.275 143.675 ;
        RECT -5.605 141.675 -5.275 142.005 ;
        RECT -5.605 140.185 -5.275 140.515 ;
        RECT -5.605 138.515 -5.275 138.845 ;
        RECT -5.605 137.025 -5.275 137.355 ;
        RECT -5.605 135.355 -5.275 135.685 ;
        RECT -5.605 133.865 -5.275 134.195 ;
        RECT -5.605 132.455 -5.275 132.785 ;
        RECT -5.605 130.615 -5.275 130.945 ;
        RECT -5.605 129.125 -5.275 129.455 ;
        RECT -5.605 127.455 -5.275 127.785 ;
        RECT -5.605 125.965 -5.275 126.295 ;
        RECT -5.605 124.295 -5.275 124.625 ;
        RECT -5.605 122.805 -5.275 123.135 ;
        RECT -5.605 121.135 -5.275 121.465 ;
        RECT -5.605 119.645 -5.275 119.975 ;
        RECT -5.605 118.235 -5.275 118.565 ;
        RECT -5.605 116.395 -5.275 116.725 ;
        RECT -5.605 114.905 -5.275 115.235 ;
        RECT -5.605 113.235 -5.275 113.565 ;
        RECT -5.605 111.745 -5.275 112.075 ;
        RECT -5.605 110.075 -5.275 110.405 ;
        RECT -5.605 108.585 -5.275 108.915 ;
        RECT -5.605 106.915 -5.275 107.245 ;
        RECT -5.605 105.425 -5.275 105.755 ;
        RECT -5.605 104.015 -5.275 104.345 ;
        RECT -5.605 102.175 -5.275 102.505 ;
        RECT -5.605 100.685 -5.275 101.015 ;
        RECT -5.605 99.015 -5.275 99.345 ;
        RECT -5.605 97.525 -5.275 97.855 ;
        RECT -5.605 95.855 -5.275 96.185 ;
        RECT -5.605 94.365 -5.275 94.695 ;
        RECT -5.605 92.695 -5.275 93.025 ;
        RECT -5.605 91.205 -5.275 91.535 ;
        RECT -5.605 89.795 -5.275 90.125 ;
        RECT -5.605 87.955 -5.275 88.285 ;
        RECT -5.605 86.465 -5.275 86.795 ;
        RECT -5.605 84.795 -5.275 85.125 ;
        RECT -5.605 83.305 -5.275 83.635 ;
        RECT -5.605 81.635 -5.275 81.965 ;
        RECT -5.605 80.145 -5.275 80.475 ;
        RECT -5.605 78.475 -5.275 78.805 ;
        RECT -5.605 76.985 -5.275 77.315 ;
        RECT -5.605 75.575 -5.275 75.905 ;
        RECT -5.605 73.735 -5.275 74.065 ;
        RECT -5.605 72.245 -5.275 72.575 ;
        RECT -5.605 70.575 -5.275 70.905 ;
        RECT -5.605 69.085 -5.275 69.415 ;
        RECT -5.605 67.415 -5.275 67.745 ;
        RECT -5.605 65.925 -5.275 66.255 ;
        RECT -5.605 64.255 -5.275 64.585 ;
        RECT -5.605 62.765 -5.275 63.095 ;
        RECT -5.605 61.355 -5.275 61.685 ;
        RECT -5.605 59.515 -5.275 59.845 ;
        RECT -5.605 58.025 -5.275 58.355 ;
        RECT -5.605 56.355 -5.275 56.685 ;
        RECT -5.605 54.865 -5.275 55.195 ;
        RECT -5.605 53.195 -5.275 53.525 ;
        RECT -5.605 51.705 -5.275 52.035 ;
        RECT -5.605 50.035 -5.275 50.365 ;
        RECT -5.605 48.545 -5.275 48.875 ;
        RECT -5.605 47.135 -5.275 47.465 ;
        RECT -5.605 45.295 -5.275 45.625 ;
        RECT -5.605 43.805 -5.275 44.135 ;
        RECT -5.605 42.135 -5.275 42.465 ;
        RECT -5.605 40.645 -5.275 40.975 ;
        RECT -5.605 38.975 -5.275 39.305 ;
        RECT -5.605 37.485 -5.275 37.815 ;
        RECT -5.605 35.815 -5.275 36.145 ;
        RECT -5.605 34.325 -5.275 34.655 ;
        RECT -5.605 32.915 -5.275 33.245 ;
        RECT -5.605 31.075 -5.275 31.405 ;
        RECT -5.605 29.585 -5.275 29.915 ;
        RECT -5.605 27.915 -5.275 28.245 ;
        RECT -5.605 26.425 -5.275 26.755 ;
        RECT -5.605 24.755 -5.275 25.085 ;
        RECT -5.605 23.265 -5.275 23.595 ;
        RECT -5.605 21.595 -5.275 21.925 ;
        RECT -5.605 20.105 -5.275 20.435 ;
        RECT -5.605 18.695 -5.275 19.025 ;
        RECT -5.605 16.855 -5.275 17.185 ;
        RECT -5.605 15.365 -5.275 15.695 ;
        RECT -5.605 13.695 -5.275 14.025 ;
        RECT -5.605 12.205 -5.275 12.535 ;
        RECT -5.605 10.535 -5.275 10.865 ;
        RECT -5.605 9.045 -5.275 9.375 ;
        RECT -5.605 7.375 -5.275 7.705 ;
        RECT -5.605 5.885 -5.275 6.215 ;
        RECT -5.605 4.475 -5.275 4.805 ;
        RECT -5.605 2.115 -5.275 2.445 ;
        RECT -5.605 0.06 -5.275 0.39 ;
        RECT -5.605 -1.525 -5.275 -1.195 ;
        RECT -5.605 -2.885 -5.275 -2.555 ;
        RECT -5.605 -4.245 -5.275 -3.915 ;
        RECT -5.605 -5.605 -5.275 -5.275 ;
        RECT -5.605 -6.965 -5.275 -6.635 ;
        RECT -5.605 -8.325 -5.275 -7.995 ;
        RECT -5.605 -9.685 -5.275 -9.355 ;
        RECT -5.605 -12.405 -5.275 -12.075 ;
        RECT -5.605 -13.765 -5.275 -13.435 ;
        RECT -5.605 -15.125 -5.275 -14.795 ;
        RECT -5.605 -16.485 -5.275 -16.155 ;
        RECT -5.605 -17.845 -5.275 -17.515 ;
        RECT -5.605 -21.925 -5.275 -21.595 ;
        RECT -5.605 -23.285 -5.275 -22.955 ;
        RECT -5.605 -24.645 -5.275 -24.315 ;
        RECT -5.605 -26.005 -5.275 -25.675 ;
        RECT -5.605 -27.365 -5.275 -27.035 ;
        RECT -5.605 -28.725 -5.275 -28.395 ;
        RECT -5.605 -30.085 -5.275 -29.755 ;
        RECT -5.605 -31.445 -5.275 -31.115 ;
        RECT -5.605 -32.805 -5.275 -32.475 ;
        RECT -5.605 -34.165 -5.275 -33.835 ;
        RECT -5.605 -36.885 -5.275 -36.555 ;
        RECT -5.605 -38.245 -5.275 -37.915 ;
        RECT -5.605 -40.965 -5.275 -40.635 ;
        RECT -5.605 -42.325 -5.275 -41.995 ;
        RECT -5.605 -43.685 -5.275 -43.355 ;
        RECT -5.605 -45.045 -5.275 -44.715 ;
        RECT -5.605 -46.405 -5.275 -46.075 ;
        RECT -5.605 -47.765 -5.275 -47.435 ;
        RECT -5.605 -49.125 -5.275 -48.795 ;
        RECT -5.605 -51.845 -5.275 -51.515 ;
        RECT -5.605 -53.205 -5.275 -52.875 ;
        RECT -5.605 -54.565 -5.275 -54.235 ;
        RECT -5.605 -55.925 -5.275 -55.595 ;
        RECT -5.605 -57.285 -5.275 -56.955 ;
        RECT -5.605 -58.645 -5.275 -58.315 ;
        RECT -5.605 -60.005 -5.275 -59.675 ;
        RECT -5.605 -61.365 -5.275 -61.035 ;
        RECT -5.605 -62.725 -5.275 -62.395 ;
        RECT -5.605 -64.085 -5.275 -63.755 ;
        RECT -5.605 -65.445 -5.275 -65.115 ;
        RECT -5.605 -66.805 -5.275 -66.475 ;
        RECT -5.605 -68.165 -5.275 -67.835 ;
        RECT -5.605 -69.525 -5.275 -69.195 ;
        RECT -5.605 -70.885 -5.275 -70.555 ;
        RECT -5.605 -72.245 -5.275 -71.915 ;
        RECT -5.605 -73.605 -5.275 -73.275 ;
        RECT -5.605 -74.965 -5.275 -74.635 ;
        RECT -5.605 -76.325 -5.275 -75.995 ;
        RECT -5.605 -77.685 -5.275 -77.355 ;
        RECT -5.605 -79.045 -5.275 -78.715 ;
        RECT -5.605 -80.405 -5.275 -80.075 ;
        RECT -5.605 -81.765 -5.275 -81.435 ;
        RECT -5.605 -83.125 -5.275 -82.795 ;
        RECT -5.605 -84.485 -5.275 -84.155 ;
        RECT -5.605 -85.845 -5.275 -85.515 ;
        RECT -5.605 -87.205 -5.275 -86.875 ;
        RECT -5.605 -88.565 -5.275 -88.235 ;
        RECT -5.605 -89.925 -5.275 -89.595 ;
        RECT -5.605 -91.285 -5.275 -90.955 ;
        RECT -5.605 -92.645 -5.275 -92.315 ;
        RECT -5.605 -94.005 -5.275 -93.675 ;
        RECT -5.605 -95.365 -5.275 -95.035 ;
        RECT -5.605 -96.725 -5.275 -96.395 ;
        RECT -5.605 -98.085 -5.275 -97.755 ;
        RECT -5.605 -99.445 -5.275 -99.115 ;
        RECT -5.605 -100.805 -5.275 -100.475 ;
        RECT -5.605 -102.165 -5.275 -101.835 ;
        RECT -5.605 -103.525 -5.275 -103.195 ;
        RECT -5.605 -104.885 -5.275 -104.555 ;
        RECT -5.605 -106.245 -5.275 -105.915 ;
        RECT -5.605 -107.605 -5.275 -107.275 ;
    END
    PORT
      LAYER met3 ;
        RECT -19.205 -27.365 -18.875 -27.035 ;
        RECT -19.205 -28.725 -18.875 -28.395 ;
        RECT -19.205 -30.085 -18.875 -29.755 ;
        RECT -19.205 -31.445 -18.875 -31.115 ;
        RECT -19.205 -32.805 -18.875 -32.475 ;
        RECT -19.205 -35.525 -18.875 -35.195 ;
        RECT -19.205 -36.885 -18.875 -36.555 ;
        RECT -19.205 -37.93 -18.875 -37.6 ;
        RECT -19.205 -40.965 -18.875 -40.635 ;
        RECT -19.205 -42.77 -18.875 -42.44 ;
        RECT -19.205 -43.685 -18.875 -43.355 ;
        RECT -19.205 -50.485 -18.875 -50.155 ;
        RECT -19.205 -51.845 -18.875 -51.515 ;
        RECT -19.205 -53.205 -18.875 -52.875 ;
        RECT -19.205 -54.565 -18.875 -54.235 ;
        RECT -19.205 -55.925 -18.875 -55.595 ;
        RECT -19.205 -57.285 -18.875 -56.955 ;
        RECT -19.205 -58.645 -18.875 -58.315 ;
        RECT -19.205 -60.005 -18.875 -59.675 ;
        RECT -19.205 -61.365 -18.875 -61.035 ;
        RECT -19.205 -62.725 -18.875 -62.395 ;
        RECT -19.205 -64.085 -18.875 -63.755 ;
        RECT -19.205 -65.445 -18.875 -65.115 ;
        RECT -19.205 -66.805 -18.875 -66.475 ;
        RECT -19.205 -68.165 -18.875 -67.835 ;
        RECT -19.205 -69.525 -18.875 -69.195 ;
        RECT -19.205 -70.885 -18.875 -70.555 ;
        RECT -19.205 -72.245 -18.875 -71.915 ;
        RECT -19.205 -74.965 -18.875 -74.635 ;
        RECT -19.205 -76.71 -18.875 -76.38 ;
        RECT -19.205 -77.685 -18.875 -77.355 ;
        RECT -19.205 -79.045 -18.875 -78.715 ;
        RECT -19.205 -81.765 -18.875 -81.435 ;
        RECT -19.205 -83.125 -18.875 -82.795 ;
        RECT -19.205 -84.485 -18.875 -84.155 ;
        RECT -19.205 -85.25 -18.875 -84.92 ;
        RECT -19.205 -87.205 -18.875 -86.875 ;
        RECT -19.205 -89.925 -18.875 -89.595 ;
        RECT -19.205 -91.285 -18.875 -90.955 ;
        RECT -19.205 -92.645 -18.875 -92.315 ;
        RECT -19.205 -94.005 -18.875 -93.675 ;
        RECT -19.205 -96.725 -18.875 -96.395 ;
        RECT -19.205 -98.085 -18.875 -97.755 ;
        RECT -19.205 -98.89 -18.875 -98.56 ;
        RECT -19.205 -100.805 -18.875 -100.475 ;
        RECT -19.205 -102.165 -18.875 -101.835 ;
        RECT -19.205 -104.885 -18.875 -104.555 ;
        RECT -19.205 -106.245 -18.875 -105.915 ;
        RECT -19.205 -107.43 -18.875 -107.1 ;
        RECT -19.205 -108.965 -18.875 -108.635 ;
        RECT -19.205 -113.045 -18.875 -112.715 ;
        RECT -19.205 -114.405 -18.875 -114.075 ;
        RECT -19.205 -115.765 -18.875 -115.435 ;
        RECT -19.205 -117.125 -18.875 -116.795 ;
        RECT -19.205 -125.285 -18.875 -124.955 ;
        RECT -19.205 -134.805 -18.875 -134.475 ;
        RECT -19.205 -138.885 -18.875 -138.555 ;
        RECT -19.205 -145.685 -18.875 -145.355 ;
        RECT -19.205 -151.125 -18.875 -150.795 ;
        RECT -19.205 -152.485 -18.875 -152.155 ;
        RECT -19.205 -156.565 -18.875 -156.235 ;
        RECT -19.205 -157.925 -18.875 -157.595 ;
        RECT -19.205 -159.285 -18.875 -158.955 ;
        RECT -19.205 -160.645 -18.875 -160.315 ;
        RECT -19.205 -162.005 -18.875 -161.675 ;
        RECT -19.205 -163.365 -18.875 -163.035 ;
        RECT -19.205 -164.725 -18.875 -164.395 ;
        RECT -19.205 -166.085 -18.875 -165.755 ;
        RECT -19.205 -167.445 -18.875 -167.115 ;
        RECT -19.205 -170.165 -18.875 -169.835 ;
        RECT -19.205 -172.885 -18.875 -172.555 ;
        RECT -19.205 -174.245 -18.875 -173.915 ;
        RECT -19.205 -175.725 -18.875 -175.395 ;
        RECT -19.205 -176.965 -18.875 -176.635 ;
        RECT -19.205 -178.325 -18.875 -177.995 ;
        RECT -19.205 -180.57 -18.875 -179.44 ;
        RECT -19.2 -180.685 -18.88 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT -17.845 241.32 -17.515 242.45 ;
        RECT -17.845 239.195 -17.515 239.525 ;
        RECT -17.845 237.835 -17.515 238.165 ;
        RECT -17.845 236.475 -17.515 236.805 ;
        RECT -17.845 235.115 -17.515 235.445 ;
        RECT -17.845 233.755 -17.515 234.085 ;
        RECT -17.845 232.395 -17.515 232.725 ;
        RECT -17.845 231.035 -17.515 231.365 ;
        RECT -17.845 229.675 -17.515 230.005 ;
        RECT -17.845 228.315 -17.515 228.645 ;
        RECT -17.845 226.955 -17.515 227.285 ;
        RECT -17.845 225.595 -17.515 225.925 ;
        RECT -17.845 224.235 -17.515 224.565 ;
        RECT -17.845 222.875 -17.515 223.205 ;
        RECT -17.845 221.515 -17.515 221.845 ;
        RECT -17.845 220.155 -17.515 220.485 ;
        RECT -17.845 218.795 -17.515 219.125 ;
        RECT -17.845 217.435 -17.515 217.765 ;
        RECT -17.845 216.075 -17.515 216.405 ;
        RECT -17.845 214.715 -17.515 215.045 ;
        RECT -17.845 213.355 -17.515 213.685 ;
        RECT -17.845 211.995 -17.515 212.325 ;
        RECT -17.845 210.635 -17.515 210.965 ;
        RECT -17.845 209.275 -17.515 209.605 ;
        RECT -17.845 207.915 -17.515 208.245 ;
        RECT -17.845 206.555 -17.515 206.885 ;
        RECT -17.845 205.195 -17.515 205.525 ;
        RECT -17.845 203.835 -17.515 204.165 ;
        RECT -17.845 202.475 -17.515 202.805 ;
        RECT -17.845 201.115 -17.515 201.445 ;
        RECT -17.845 199.755 -17.515 200.085 ;
        RECT -17.845 198.395 -17.515 198.725 ;
        RECT -17.845 197.035 -17.515 197.365 ;
        RECT -17.845 195.675 -17.515 196.005 ;
        RECT -17.845 194.315 -17.515 194.645 ;
        RECT -17.845 192.955 -17.515 193.285 ;
        RECT -17.845 191.595 -17.515 191.925 ;
        RECT -17.845 190.235 -17.515 190.565 ;
        RECT -17.845 188.875 -17.515 189.205 ;
        RECT -17.845 187.515 -17.515 187.845 ;
        RECT -17.845 186.155 -17.515 186.485 ;
        RECT -17.845 184.795 -17.515 185.125 ;
        RECT -17.845 183.435 -17.515 183.765 ;
        RECT -17.845 182.075 -17.515 182.405 ;
        RECT -17.845 180.715 -17.515 181.045 ;
        RECT -17.845 179.355 -17.515 179.685 ;
        RECT -17.845 177.995 -17.515 178.325 ;
        RECT -17.845 176.635 -17.515 176.965 ;
        RECT -17.845 175.275 -17.515 175.605 ;
        RECT -17.845 173.915 -17.515 174.245 ;
        RECT -17.845 172.555 -17.515 172.885 ;
        RECT -17.845 171.195 -17.515 171.525 ;
        RECT -17.845 169.835 -17.515 170.165 ;
        RECT -17.845 168.475 -17.515 168.805 ;
        RECT -17.845 167.115 -17.515 167.445 ;
        RECT -17.845 165.755 -17.515 166.085 ;
        RECT -17.845 164.395 -17.515 164.725 ;
        RECT -17.845 163.035 -17.515 163.365 ;
        RECT -17.845 161.675 -17.515 162.005 ;
        RECT -17.845 160.315 -17.515 160.645 ;
        RECT -17.845 158.955 -17.515 159.285 ;
        RECT -17.845 157.595 -17.515 157.925 ;
        RECT -17.845 156.235 -17.515 156.565 ;
        RECT -17.845 154.875 -17.515 155.205 ;
        RECT -17.845 153.515 -17.515 153.845 ;
        RECT -17.845 152.155 -17.515 152.485 ;
        RECT -17.845 150.795 -17.515 151.125 ;
        RECT -17.845 149.435 -17.515 149.765 ;
        RECT -17.845 148.075 -17.515 148.405 ;
        RECT -17.845 146.715 -17.515 147.045 ;
        RECT -17.845 145.355 -17.515 145.685 ;
        RECT -17.845 143.995 -17.515 144.325 ;
        RECT -17.845 142.635 -17.515 142.965 ;
        RECT -17.845 141.275 -17.515 141.605 ;
        RECT -17.845 139.915 -17.515 140.245 ;
        RECT -17.845 138.555 -17.515 138.885 ;
        RECT -17.845 137.195 -17.515 137.525 ;
        RECT -17.845 135.835 -17.515 136.165 ;
        RECT -17.845 134.475 -17.515 134.805 ;
        RECT -17.845 133.115 -17.515 133.445 ;
        RECT -17.845 131.755 -17.515 132.085 ;
        RECT -17.845 130.395 -17.515 130.725 ;
        RECT -17.845 129.035 -17.515 129.365 ;
        RECT -17.845 127.675 -17.515 128.005 ;
        RECT -17.845 126.315 -17.515 126.645 ;
        RECT -17.845 124.955 -17.515 125.285 ;
        RECT -17.845 123.595 -17.515 123.925 ;
        RECT -17.845 122.235 -17.515 122.565 ;
        RECT -17.845 120.875 -17.515 121.205 ;
        RECT -17.845 119.515 -17.515 119.845 ;
        RECT -17.845 118.155 -17.515 118.485 ;
        RECT -17.845 116.795 -17.515 117.125 ;
        RECT -17.845 115.435 -17.515 115.765 ;
        RECT -17.845 114.075 -17.515 114.405 ;
        RECT -17.845 112.715 -17.515 113.045 ;
        RECT -17.845 111.355 -17.515 111.685 ;
        RECT -17.845 109.995 -17.515 110.325 ;
        RECT -17.845 108.635 -17.515 108.965 ;
        RECT -17.845 107.275 -17.515 107.605 ;
        RECT -17.845 105.915 -17.515 106.245 ;
        RECT -17.845 104.555 -17.515 104.885 ;
        RECT -17.845 103.195 -17.515 103.525 ;
        RECT -17.845 101.835 -17.515 102.165 ;
        RECT -17.845 100.475 -17.515 100.805 ;
        RECT -17.845 99.115 -17.515 99.445 ;
        RECT -17.845 97.755 -17.515 98.085 ;
        RECT -17.845 96.395 -17.515 96.725 ;
        RECT -17.845 95.035 -17.515 95.365 ;
        RECT -17.845 93.675 -17.515 94.005 ;
        RECT -17.845 92.315 -17.515 92.645 ;
        RECT -17.845 90.955 -17.515 91.285 ;
        RECT -17.845 89.595 -17.515 89.925 ;
        RECT -17.845 88.235 -17.515 88.565 ;
        RECT -17.845 86.875 -17.515 87.205 ;
        RECT -17.845 85.515 -17.515 85.845 ;
        RECT -17.845 84.155 -17.515 84.485 ;
        RECT -17.845 82.795 -17.515 83.125 ;
        RECT -17.845 81.435 -17.515 81.765 ;
        RECT -17.845 80.075 -17.515 80.405 ;
        RECT -17.845 78.715 -17.515 79.045 ;
        RECT -17.845 77.355 -17.515 77.685 ;
        RECT -17.845 75.995 -17.515 76.325 ;
        RECT -17.845 74.635 -17.515 74.965 ;
        RECT -17.845 73.275 -17.515 73.605 ;
        RECT -17.845 71.915 -17.515 72.245 ;
        RECT -17.845 70.555 -17.515 70.885 ;
        RECT -17.845 69.195 -17.515 69.525 ;
        RECT -17.845 67.835 -17.515 68.165 ;
        RECT -17.845 66.475 -17.515 66.805 ;
        RECT -17.845 65.115 -17.515 65.445 ;
        RECT -17.845 63.755 -17.515 64.085 ;
        RECT -17.845 62.395 -17.515 62.725 ;
        RECT -17.845 61.035 -17.515 61.365 ;
        RECT -17.845 59.675 -17.515 60.005 ;
        RECT -17.845 58.315 -17.515 58.645 ;
        RECT -17.845 56.955 -17.515 57.285 ;
        RECT -17.845 55.595 -17.515 55.925 ;
        RECT -17.845 54.235 -17.515 54.565 ;
        RECT -17.845 52.875 -17.515 53.205 ;
        RECT -17.845 51.515 -17.515 51.845 ;
        RECT -17.845 50.155 -17.515 50.485 ;
        RECT -17.845 48.795 -17.515 49.125 ;
        RECT -17.845 47.435 -17.515 47.765 ;
        RECT -17.845 46.075 -17.515 46.405 ;
        RECT -17.845 44.715 -17.515 45.045 ;
        RECT -17.845 43.355 -17.515 43.685 ;
        RECT -17.845 41.995 -17.515 42.325 ;
        RECT -17.845 40.635 -17.515 40.965 ;
        RECT -17.845 39.275 -17.515 39.605 ;
        RECT -17.845 37.915 -17.515 38.245 ;
        RECT -17.845 36.555 -17.515 36.885 ;
        RECT -17.845 35.195 -17.515 35.525 ;
        RECT -17.845 33.835 -17.515 34.165 ;
        RECT -17.845 32.475 -17.515 32.805 ;
        RECT -17.845 31.115 -17.515 31.445 ;
        RECT -17.845 29.755 -17.515 30.085 ;
        RECT -17.845 28.395 -17.515 28.725 ;
        RECT -17.845 27.035 -17.515 27.365 ;
        RECT -17.845 25.675 -17.515 26.005 ;
        RECT -17.845 24.315 -17.515 24.645 ;
        RECT -17.845 22.955 -17.515 23.285 ;
        RECT -17.845 21.595 -17.515 21.925 ;
        RECT -17.845 20.235 -17.515 20.565 ;
        RECT -17.845 18.875 -17.515 19.205 ;
        RECT -17.845 17.515 -17.515 17.845 ;
        RECT -17.845 16.155 -17.515 16.485 ;
        RECT -17.845 14.795 -17.515 15.125 ;
        RECT -17.845 13.435 -17.515 13.765 ;
        RECT -17.845 12.075 -17.515 12.405 ;
        RECT -17.845 10.715 -17.515 11.045 ;
        RECT -17.845 9.355 -17.515 9.685 ;
        RECT -17.845 7.995 -17.515 8.325 ;
        RECT -17.845 6.635 -17.515 6.965 ;
        RECT -17.845 5.275 -17.515 5.605 ;
        RECT -17.845 3.915 -17.515 4.245 ;
        RECT -17.845 2.555 -17.515 2.885 ;
        RECT -17.845 1.195 -17.515 1.525 ;
        RECT -17.845 -0.165 -17.515 0.165 ;
        RECT -17.845 -2.885 -17.515 -2.555 ;
        RECT -17.845 -4.245 -17.515 -3.915 ;
        RECT -17.845 -8.325 -17.515 -7.995 ;
        RECT -17.845 -9.685 -17.515 -9.355 ;
        RECT -17.84 -11.04 -17.52 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -17.845 -27.365 -17.515 -27.035 ;
        RECT -17.845 -28.725 -17.515 -28.395 ;
        RECT -17.845 -30.085 -17.515 -29.755 ;
        RECT -17.845 -31.445 -17.515 -31.115 ;
        RECT -17.845 -32.805 -17.515 -32.475 ;
        RECT -17.845 -36.885 -17.515 -36.555 ;
        RECT -17.845 -37.93 -17.515 -37.6 ;
        RECT -17.845 -40.965 -17.515 -40.635 ;
        RECT -17.845 -42.77 -17.515 -42.44 ;
        RECT -17.845 -43.685 -17.515 -43.355 ;
        RECT -17.845 -50.485 -17.515 -50.155 ;
        RECT -17.845 -51.845 -17.515 -51.515 ;
        RECT -17.845 -53.205 -17.515 -52.875 ;
        RECT -17.845 -54.565 -17.515 -54.235 ;
        RECT -17.845 -55.925 -17.515 -55.595 ;
        RECT -17.845 -57.285 -17.515 -56.955 ;
        RECT -17.845 -58.645 -17.515 -58.315 ;
        RECT -17.845 -60.005 -17.515 -59.675 ;
        RECT -17.845 -61.365 -17.515 -61.035 ;
        RECT -17.845 -62.725 -17.515 -62.395 ;
        RECT -17.845 -64.085 -17.515 -63.755 ;
        RECT -17.845 -65.445 -17.515 -65.115 ;
        RECT -17.845 -66.805 -17.515 -66.475 ;
        RECT -17.845 -68.165 -17.515 -67.835 ;
        RECT -17.845 -69.525 -17.515 -69.195 ;
        RECT -17.845 -70.885 -17.515 -70.555 ;
        RECT -17.845 -72.245 -17.515 -71.915 ;
        RECT -17.845 -74.965 -17.515 -74.635 ;
        RECT -17.845 -76.71 -17.515 -76.38 ;
        RECT -17.845 -77.685 -17.515 -77.355 ;
        RECT -17.845 -79.045 -17.515 -78.715 ;
        RECT -17.845 -81.765 -17.515 -81.435 ;
        RECT -17.845 -83.125 -17.515 -82.795 ;
        RECT -17.845 -84.485 -17.515 -84.155 ;
        RECT -17.845 -85.25 -17.515 -84.92 ;
        RECT -17.845 -87.205 -17.515 -86.875 ;
        RECT -17.845 -89.925 -17.515 -89.595 ;
        RECT -17.845 -91.285 -17.515 -90.955 ;
        RECT -17.845 -92.645 -17.515 -92.315 ;
        RECT -17.845 -94.005 -17.515 -93.675 ;
        RECT -17.845 -96.725 -17.515 -96.395 ;
        RECT -17.845 -98.085 -17.515 -97.755 ;
        RECT -17.845 -98.89 -17.515 -98.56 ;
        RECT -17.845 -100.805 -17.515 -100.475 ;
        RECT -17.845 -102.165 -17.515 -101.835 ;
        RECT -17.845 -104.885 -17.515 -104.555 ;
        RECT -17.845 -106.245 -17.515 -105.915 ;
        RECT -17.845 -107.43 -17.515 -107.1 ;
        RECT -17.845 -114.405 -17.515 -114.075 ;
        RECT -17.845 -115.765 -17.515 -115.435 ;
        RECT -17.845 -117.125 -17.515 -116.795 ;
        RECT -17.845 -125.285 -17.515 -124.955 ;
        RECT -17.845 -138.885 -17.515 -138.555 ;
        RECT -17.845 -144.325 -17.515 -143.995 ;
        RECT -17.845 -145.685 -17.515 -145.355 ;
        RECT -17.845 -151.125 -17.515 -150.795 ;
        RECT -17.845 -152.485 -17.515 -152.155 ;
        RECT -17.845 -156.565 -17.515 -156.235 ;
        RECT -17.845 -157.925 -17.515 -157.595 ;
        RECT -17.845 -159.285 -17.515 -158.955 ;
        RECT -17.845 -160.645 -17.515 -160.315 ;
        RECT -17.845 -162.005 -17.515 -161.675 ;
        RECT -17.845 -163.365 -17.515 -163.035 ;
        RECT -17.845 -164.725 -17.515 -164.395 ;
        RECT -17.845 -166.085 -17.515 -165.755 ;
        RECT -17.845 -167.445 -17.515 -167.115 ;
        RECT -17.845 -170.165 -17.515 -169.835 ;
        RECT -17.845 -174.245 -17.515 -173.915 ;
        RECT -17.845 -175.725 -17.515 -175.395 ;
        RECT -17.845 -176.965 -17.515 -176.635 ;
        RECT -17.845 -178.325 -17.515 -177.995 ;
        RECT -17.845 -180.57 -17.515 -179.44 ;
        RECT -17.84 -180.685 -17.52 -26.36 ;
    END
    PORT
      LAYER met3 ;
        RECT -16.485 241.32 -16.155 242.45 ;
        RECT -16.485 239.195 -16.155 239.525 ;
        RECT -16.485 237.835 -16.155 238.165 ;
        RECT -16.485 236.475 -16.155 236.805 ;
        RECT -16.485 235.115 -16.155 235.445 ;
        RECT -16.485 233.755 -16.155 234.085 ;
        RECT -16.485 232.395 -16.155 232.725 ;
        RECT -16.485 231.035 -16.155 231.365 ;
        RECT -16.485 229.675 -16.155 230.005 ;
        RECT -16.485 228.315 -16.155 228.645 ;
        RECT -16.485 226.955 -16.155 227.285 ;
        RECT -16.485 225.595 -16.155 225.925 ;
        RECT -16.485 224.235 -16.155 224.565 ;
        RECT -16.485 222.875 -16.155 223.205 ;
        RECT -16.485 221.515 -16.155 221.845 ;
        RECT -16.485 220.155 -16.155 220.485 ;
        RECT -16.485 218.795 -16.155 219.125 ;
        RECT -16.485 217.435 -16.155 217.765 ;
        RECT -16.485 216.075 -16.155 216.405 ;
        RECT -16.485 214.715 -16.155 215.045 ;
        RECT -16.485 213.355 -16.155 213.685 ;
        RECT -16.485 211.995 -16.155 212.325 ;
        RECT -16.485 210.635 -16.155 210.965 ;
        RECT -16.485 209.275 -16.155 209.605 ;
        RECT -16.485 207.915 -16.155 208.245 ;
        RECT -16.485 206.555 -16.155 206.885 ;
        RECT -16.485 205.195 -16.155 205.525 ;
        RECT -16.485 203.835 -16.155 204.165 ;
        RECT -16.485 202.475 -16.155 202.805 ;
        RECT -16.485 201.115 -16.155 201.445 ;
        RECT -16.485 199.755 -16.155 200.085 ;
        RECT -16.485 198.395 -16.155 198.725 ;
        RECT -16.485 197.035 -16.155 197.365 ;
        RECT -16.485 195.675 -16.155 196.005 ;
        RECT -16.485 194.315 -16.155 194.645 ;
        RECT -16.485 192.955 -16.155 193.285 ;
        RECT -16.485 191.595 -16.155 191.925 ;
        RECT -16.485 190.235 -16.155 190.565 ;
        RECT -16.485 188.875 -16.155 189.205 ;
        RECT -16.485 187.515 -16.155 187.845 ;
        RECT -16.485 186.155 -16.155 186.485 ;
        RECT -16.485 184.795 -16.155 185.125 ;
        RECT -16.485 183.435 -16.155 183.765 ;
        RECT -16.485 182.075 -16.155 182.405 ;
        RECT -16.485 180.715 -16.155 181.045 ;
        RECT -16.485 179.355 -16.155 179.685 ;
        RECT -16.485 177.995 -16.155 178.325 ;
        RECT -16.485 176.635 -16.155 176.965 ;
        RECT -16.485 175.275 -16.155 175.605 ;
        RECT -16.485 173.915 -16.155 174.245 ;
        RECT -16.485 172.555 -16.155 172.885 ;
        RECT -16.485 171.195 -16.155 171.525 ;
        RECT -16.485 169.835 -16.155 170.165 ;
        RECT -16.485 168.475 -16.155 168.805 ;
        RECT -16.485 167.115 -16.155 167.445 ;
        RECT -16.485 165.755 -16.155 166.085 ;
        RECT -16.485 164.395 -16.155 164.725 ;
        RECT -16.485 163.035 -16.155 163.365 ;
        RECT -16.485 161.675 -16.155 162.005 ;
        RECT -16.485 160.315 -16.155 160.645 ;
        RECT -16.485 158.955 -16.155 159.285 ;
        RECT -16.485 157.595 -16.155 157.925 ;
        RECT -16.485 156.235 -16.155 156.565 ;
        RECT -16.485 154.875 -16.155 155.205 ;
        RECT -16.485 153.515 -16.155 153.845 ;
        RECT -16.485 152.155 -16.155 152.485 ;
        RECT -16.485 150.795 -16.155 151.125 ;
        RECT -16.485 149.435 -16.155 149.765 ;
        RECT -16.485 148.075 -16.155 148.405 ;
        RECT -16.485 146.715 -16.155 147.045 ;
        RECT -16.485 145.355 -16.155 145.685 ;
        RECT -16.485 143.995 -16.155 144.325 ;
        RECT -16.485 142.635 -16.155 142.965 ;
        RECT -16.485 141.275 -16.155 141.605 ;
        RECT -16.485 139.915 -16.155 140.245 ;
        RECT -16.485 138.555 -16.155 138.885 ;
        RECT -16.485 137.195 -16.155 137.525 ;
        RECT -16.485 135.835 -16.155 136.165 ;
        RECT -16.485 134.475 -16.155 134.805 ;
        RECT -16.485 133.115 -16.155 133.445 ;
        RECT -16.485 131.755 -16.155 132.085 ;
        RECT -16.485 130.395 -16.155 130.725 ;
        RECT -16.485 129.035 -16.155 129.365 ;
        RECT -16.485 127.675 -16.155 128.005 ;
        RECT -16.485 126.315 -16.155 126.645 ;
        RECT -16.485 124.955 -16.155 125.285 ;
        RECT -16.485 123.595 -16.155 123.925 ;
        RECT -16.485 122.235 -16.155 122.565 ;
        RECT -16.485 120.875 -16.155 121.205 ;
        RECT -16.485 119.515 -16.155 119.845 ;
        RECT -16.485 118.155 -16.155 118.485 ;
        RECT -16.485 116.795 -16.155 117.125 ;
        RECT -16.485 115.435 -16.155 115.765 ;
        RECT -16.485 114.075 -16.155 114.405 ;
        RECT -16.485 112.715 -16.155 113.045 ;
        RECT -16.485 111.355 -16.155 111.685 ;
        RECT -16.485 109.995 -16.155 110.325 ;
        RECT -16.485 108.635 -16.155 108.965 ;
        RECT -16.485 107.275 -16.155 107.605 ;
        RECT -16.485 105.915 -16.155 106.245 ;
        RECT -16.485 104.555 -16.155 104.885 ;
        RECT -16.485 103.195 -16.155 103.525 ;
        RECT -16.485 101.835 -16.155 102.165 ;
        RECT -16.485 100.475 -16.155 100.805 ;
        RECT -16.485 99.115 -16.155 99.445 ;
        RECT -16.485 97.755 -16.155 98.085 ;
        RECT -16.485 96.395 -16.155 96.725 ;
        RECT -16.485 95.035 -16.155 95.365 ;
        RECT -16.485 93.675 -16.155 94.005 ;
        RECT -16.485 92.315 -16.155 92.645 ;
        RECT -16.485 90.955 -16.155 91.285 ;
        RECT -16.485 89.595 -16.155 89.925 ;
        RECT -16.485 88.235 -16.155 88.565 ;
        RECT -16.485 86.875 -16.155 87.205 ;
        RECT -16.485 85.515 -16.155 85.845 ;
        RECT -16.485 84.155 -16.155 84.485 ;
        RECT -16.485 82.795 -16.155 83.125 ;
        RECT -16.485 81.435 -16.155 81.765 ;
        RECT -16.485 80.075 -16.155 80.405 ;
        RECT -16.485 78.715 -16.155 79.045 ;
        RECT -16.485 77.355 -16.155 77.685 ;
        RECT -16.485 75.995 -16.155 76.325 ;
        RECT -16.485 74.635 -16.155 74.965 ;
        RECT -16.485 73.275 -16.155 73.605 ;
        RECT -16.485 71.915 -16.155 72.245 ;
        RECT -16.485 70.555 -16.155 70.885 ;
        RECT -16.485 69.195 -16.155 69.525 ;
        RECT -16.485 67.835 -16.155 68.165 ;
        RECT -16.485 66.475 -16.155 66.805 ;
        RECT -16.485 65.115 -16.155 65.445 ;
        RECT -16.485 63.755 -16.155 64.085 ;
        RECT -16.485 62.395 -16.155 62.725 ;
        RECT -16.485 61.035 -16.155 61.365 ;
        RECT -16.485 59.675 -16.155 60.005 ;
        RECT -16.485 58.315 -16.155 58.645 ;
        RECT -16.485 56.955 -16.155 57.285 ;
        RECT -16.485 55.595 -16.155 55.925 ;
        RECT -16.485 54.235 -16.155 54.565 ;
        RECT -16.485 52.875 -16.155 53.205 ;
        RECT -16.485 51.515 -16.155 51.845 ;
        RECT -16.485 50.155 -16.155 50.485 ;
        RECT -16.485 48.795 -16.155 49.125 ;
        RECT -16.485 47.435 -16.155 47.765 ;
        RECT -16.485 46.075 -16.155 46.405 ;
        RECT -16.485 44.715 -16.155 45.045 ;
        RECT -16.485 43.355 -16.155 43.685 ;
        RECT -16.485 41.995 -16.155 42.325 ;
        RECT -16.485 40.635 -16.155 40.965 ;
        RECT -16.485 39.275 -16.155 39.605 ;
        RECT -16.485 37.915 -16.155 38.245 ;
        RECT -16.485 36.555 -16.155 36.885 ;
        RECT -16.485 35.195 -16.155 35.525 ;
        RECT -16.485 33.835 -16.155 34.165 ;
        RECT -16.485 32.475 -16.155 32.805 ;
        RECT -16.485 31.115 -16.155 31.445 ;
        RECT -16.485 29.755 -16.155 30.085 ;
        RECT -16.485 28.395 -16.155 28.725 ;
        RECT -16.485 27.035 -16.155 27.365 ;
        RECT -16.485 25.675 -16.155 26.005 ;
        RECT -16.485 24.315 -16.155 24.645 ;
        RECT -16.485 22.955 -16.155 23.285 ;
        RECT -16.485 21.595 -16.155 21.925 ;
        RECT -16.485 20.235 -16.155 20.565 ;
        RECT -16.485 18.875 -16.155 19.205 ;
        RECT -16.485 17.515 -16.155 17.845 ;
        RECT -16.485 16.155 -16.155 16.485 ;
        RECT -16.485 14.795 -16.155 15.125 ;
        RECT -16.485 13.435 -16.155 13.765 ;
        RECT -16.485 12.075 -16.155 12.405 ;
        RECT -16.485 10.715 -16.155 11.045 ;
        RECT -16.485 9.355 -16.155 9.685 ;
        RECT -16.485 7.995 -16.155 8.325 ;
        RECT -16.485 6.635 -16.155 6.965 ;
        RECT -16.485 5.275 -16.155 5.605 ;
        RECT -16.485 3.915 -16.155 4.245 ;
        RECT -16.485 2.555 -16.155 2.885 ;
        RECT -16.485 1.195 -16.155 1.525 ;
        RECT -16.485 -0.165 -16.155 0.165 ;
        RECT -16.485 -2.885 -16.155 -2.555 ;
        RECT -16.485 -4.245 -16.155 -3.915 ;
        RECT -16.485 -5.605 -16.155 -5.275 ;
        RECT -16.485 -8.325 -16.155 -7.995 ;
        RECT -16.485 -9.685 -16.155 -9.355 ;
        RECT -16.485 -12.405 -16.155 -12.075 ;
        RECT -16.48 -12.405 -16.16 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -16.485 -27.365 -16.155 -27.035 ;
        RECT -16.485 -28.725 -16.155 -28.395 ;
        RECT -16.485 -30.085 -16.155 -29.755 ;
        RECT -16.485 -31.445 -16.155 -31.115 ;
        RECT -16.485 -32.805 -16.155 -32.475 ;
        RECT -16.485 -36.885 -16.155 -36.555 ;
        RECT -16.485 -37.93 -16.155 -37.6 ;
        RECT -16.485 -40.965 -16.155 -40.635 ;
        RECT -16.485 -42.77 -16.155 -42.44 ;
        RECT -16.485 -43.685 -16.155 -43.355 ;
        RECT -16.485 -50.485 -16.155 -50.155 ;
        RECT -16.485 -51.845 -16.155 -51.515 ;
        RECT -16.485 -53.205 -16.155 -52.875 ;
        RECT -16.485 -54.565 -16.155 -54.235 ;
        RECT -16.485 -55.925 -16.155 -55.595 ;
        RECT -16.485 -57.285 -16.155 -56.955 ;
        RECT -16.485 -58.645 -16.155 -58.315 ;
        RECT -16.485 -60.005 -16.155 -59.675 ;
        RECT -16.485 -61.365 -16.155 -61.035 ;
        RECT -16.485 -62.725 -16.155 -62.395 ;
        RECT -16.485 -64.085 -16.155 -63.755 ;
        RECT -16.485 -65.445 -16.155 -65.115 ;
        RECT -16.485 -66.805 -16.155 -66.475 ;
        RECT -16.485 -68.165 -16.155 -67.835 ;
        RECT -16.485 -69.525 -16.155 -69.195 ;
        RECT -16.485 -70.885 -16.155 -70.555 ;
        RECT -16.485 -72.245 -16.155 -71.915 ;
        RECT -16.485 -74.965 -16.155 -74.635 ;
        RECT -16.485 -76.71 -16.155 -76.38 ;
        RECT -16.485 -77.685 -16.155 -77.355 ;
        RECT -16.485 -79.045 -16.155 -78.715 ;
        RECT -16.485 -81.765 -16.155 -81.435 ;
        RECT -16.485 -83.125 -16.155 -82.795 ;
        RECT -16.485 -84.485 -16.155 -84.155 ;
        RECT -16.485 -85.25 -16.155 -84.92 ;
        RECT -16.485 -87.205 -16.155 -86.875 ;
        RECT -16.485 -89.925 -16.155 -89.595 ;
        RECT -16.485 -91.285 -16.155 -90.955 ;
        RECT -16.485 -92.645 -16.155 -92.315 ;
        RECT -16.485 -94.005 -16.155 -93.675 ;
        RECT -16.485 -96.725 -16.155 -96.395 ;
        RECT -16.485 -98.085 -16.155 -97.755 ;
        RECT -16.485 -98.89 -16.155 -98.56 ;
        RECT -16.485 -100.805 -16.155 -100.475 ;
        RECT -16.485 -102.165 -16.155 -101.835 ;
        RECT -16.485 -104.885 -16.155 -104.555 ;
        RECT -16.485 -106.245 -16.155 -105.915 ;
        RECT -16.485 -107.43 -16.155 -107.1 ;
        RECT -16.48 -110.32 -16.16 -26.36 ;
    END
    PORT
      LAYER met3 ;
        RECT -16.485 -174.245 -16.155 -173.915 ;
        RECT -16.485 -176.965 -16.155 -176.635 ;
        RECT -16.485 -178.325 -16.155 -177.995 ;
        RECT -16.485 -180.57 -16.155 -179.44 ;
        RECT -16.48 -180.685 -16.16 -173.915 ;
    END
    PORT
      LAYER met3 ;
        RECT -15.125 241.32 -14.795 242.45 ;
        RECT -15.125 239.195 -14.795 239.525 ;
        RECT -15.125 237.835 -14.795 238.165 ;
        RECT -15.125 236.475 -14.795 236.805 ;
        RECT -15.125 235.115 -14.795 235.445 ;
        RECT -15.125 233.755 -14.795 234.085 ;
        RECT -15.125 232.395 -14.795 232.725 ;
        RECT -15.125 231.035 -14.795 231.365 ;
        RECT -15.125 229.675 -14.795 230.005 ;
        RECT -15.125 228.315 -14.795 228.645 ;
        RECT -15.125 226.955 -14.795 227.285 ;
        RECT -15.125 225.595 -14.795 225.925 ;
        RECT -15.125 224.235 -14.795 224.565 ;
        RECT -15.125 222.875 -14.795 223.205 ;
        RECT -15.125 221.515 -14.795 221.845 ;
        RECT -15.125 220.155 -14.795 220.485 ;
        RECT -15.125 218.795 -14.795 219.125 ;
        RECT -15.125 217.435 -14.795 217.765 ;
        RECT -15.125 216.075 -14.795 216.405 ;
        RECT -15.125 214.715 -14.795 215.045 ;
        RECT -15.125 213.355 -14.795 213.685 ;
        RECT -15.125 211.995 -14.795 212.325 ;
        RECT -15.125 210.635 -14.795 210.965 ;
        RECT -15.125 209.275 -14.795 209.605 ;
        RECT -15.125 207.915 -14.795 208.245 ;
        RECT -15.125 206.555 -14.795 206.885 ;
        RECT -15.125 205.195 -14.795 205.525 ;
        RECT -15.125 203.835 -14.795 204.165 ;
        RECT -15.125 202.475 -14.795 202.805 ;
        RECT -15.125 201.115 -14.795 201.445 ;
        RECT -15.125 199.755 -14.795 200.085 ;
        RECT -15.125 198.395 -14.795 198.725 ;
        RECT -15.125 197.035 -14.795 197.365 ;
        RECT -15.125 195.675 -14.795 196.005 ;
        RECT -15.125 194.315 -14.795 194.645 ;
        RECT -15.125 192.955 -14.795 193.285 ;
        RECT -15.125 191.595 -14.795 191.925 ;
        RECT -15.125 190.235 -14.795 190.565 ;
        RECT -15.125 188.875 -14.795 189.205 ;
        RECT -15.125 187.515 -14.795 187.845 ;
        RECT -15.125 186.155 -14.795 186.485 ;
        RECT -15.125 184.795 -14.795 185.125 ;
        RECT -15.125 183.435 -14.795 183.765 ;
        RECT -15.125 182.075 -14.795 182.405 ;
        RECT -15.125 180.715 -14.795 181.045 ;
        RECT -15.125 179.355 -14.795 179.685 ;
        RECT -15.125 177.995 -14.795 178.325 ;
        RECT -15.125 176.635 -14.795 176.965 ;
        RECT -15.125 175.275 -14.795 175.605 ;
        RECT -15.125 173.915 -14.795 174.245 ;
        RECT -15.125 172.555 -14.795 172.885 ;
        RECT -15.125 171.195 -14.795 171.525 ;
        RECT -15.125 169.835 -14.795 170.165 ;
        RECT -15.125 168.475 -14.795 168.805 ;
        RECT -15.125 167.115 -14.795 167.445 ;
        RECT -15.125 165.755 -14.795 166.085 ;
        RECT -15.125 164.395 -14.795 164.725 ;
        RECT -15.125 163.035 -14.795 163.365 ;
        RECT -15.125 161.675 -14.795 162.005 ;
        RECT -15.125 160.315 -14.795 160.645 ;
        RECT -15.125 158.955 -14.795 159.285 ;
        RECT -15.125 157.595 -14.795 157.925 ;
        RECT -15.125 156.235 -14.795 156.565 ;
        RECT -15.125 154.875 -14.795 155.205 ;
        RECT -15.125 153.515 -14.795 153.845 ;
        RECT -15.125 152.155 -14.795 152.485 ;
        RECT -15.125 150.795 -14.795 151.125 ;
        RECT -15.125 149.435 -14.795 149.765 ;
        RECT -15.125 148.075 -14.795 148.405 ;
        RECT -15.125 146.715 -14.795 147.045 ;
        RECT -15.125 145.355 -14.795 145.685 ;
        RECT -15.125 143.995 -14.795 144.325 ;
        RECT -15.125 142.635 -14.795 142.965 ;
        RECT -15.125 141.275 -14.795 141.605 ;
        RECT -15.125 139.915 -14.795 140.245 ;
        RECT -15.125 138.555 -14.795 138.885 ;
        RECT -15.125 137.195 -14.795 137.525 ;
        RECT -15.125 135.835 -14.795 136.165 ;
        RECT -15.125 134.475 -14.795 134.805 ;
        RECT -15.125 133.115 -14.795 133.445 ;
        RECT -15.125 131.755 -14.795 132.085 ;
        RECT -15.125 130.395 -14.795 130.725 ;
        RECT -15.125 129.035 -14.795 129.365 ;
        RECT -15.125 127.675 -14.795 128.005 ;
        RECT -15.125 126.315 -14.795 126.645 ;
        RECT -15.125 124.955 -14.795 125.285 ;
        RECT -15.125 123.595 -14.795 123.925 ;
        RECT -15.125 122.235 -14.795 122.565 ;
        RECT -15.125 120.875 -14.795 121.205 ;
        RECT -15.125 119.515 -14.795 119.845 ;
        RECT -15.125 118.155 -14.795 118.485 ;
        RECT -15.125 116.795 -14.795 117.125 ;
        RECT -15.125 115.435 -14.795 115.765 ;
        RECT -15.125 114.075 -14.795 114.405 ;
        RECT -15.125 112.715 -14.795 113.045 ;
        RECT -15.125 111.355 -14.795 111.685 ;
        RECT -15.125 109.995 -14.795 110.325 ;
        RECT -15.125 108.635 -14.795 108.965 ;
        RECT -15.125 107.275 -14.795 107.605 ;
        RECT -15.125 105.915 -14.795 106.245 ;
        RECT -15.125 104.555 -14.795 104.885 ;
        RECT -15.125 103.195 -14.795 103.525 ;
        RECT -15.125 101.835 -14.795 102.165 ;
        RECT -15.125 100.475 -14.795 100.805 ;
        RECT -15.125 99.115 -14.795 99.445 ;
        RECT -15.125 97.755 -14.795 98.085 ;
        RECT -15.125 96.395 -14.795 96.725 ;
        RECT -15.125 95.035 -14.795 95.365 ;
        RECT -15.125 93.675 -14.795 94.005 ;
        RECT -15.125 92.315 -14.795 92.645 ;
        RECT -15.125 90.955 -14.795 91.285 ;
        RECT -15.125 89.595 -14.795 89.925 ;
        RECT -15.125 88.235 -14.795 88.565 ;
        RECT -15.125 86.875 -14.795 87.205 ;
        RECT -15.125 85.515 -14.795 85.845 ;
        RECT -15.125 84.155 -14.795 84.485 ;
        RECT -15.125 82.795 -14.795 83.125 ;
        RECT -15.125 81.435 -14.795 81.765 ;
        RECT -15.125 80.075 -14.795 80.405 ;
        RECT -15.125 78.715 -14.795 79.045 ;
        RECT -15.125 77.355 -14.795 77.685 ;
        RECT -15.125 75.995 -14.795 76.325 ;
        RECT -15.125 74.635 -14.795 74.965 ;
        RECT -15.125 73.275 -14.795 73.605 ;
        RECT -15.125 71.915 -14.795 72.245 ;
        RECT -15.125 70.555 -14.795 70.885 ;
        RECT -15.125 69.195 -14.795 69.525 ;
        RECT -15.125 67.835 -14.795 68.165 ;
        RECT -15.125 66.475 -14.795 66.805 ;
        RECT -15.125 65.115 -14.795 65.445 ;
        RECT -15.125 63.755 -14.795 64.085 ;
        RECT -15.125 62.395 -14.795 62.725 ;
        RECT -15.125 61.035 -14.795 61.365 ;
        RECT -15.125 59.675 -14.795 60.005 ;
        RECT -15.125 58.315 -14.795 58.645 ;
        RECT -15.125 56.955 -14.795 57.285 ;
        RECT -15.125 55.595 -14.795 55.925 ;
        RECT -15.125 54.235 -14.795 54.565 ;
        RECT -15.125 52.875 -14.795 53.205 ;
        RECT -15.125 51.515 -14.795 51.845 ;
        RECT -15.125 50.155 -14.795 50.485 ;
        RECT -15.125 48.795 -14.795 49.125 ;
        RECT -15.125 47.435 -14.795 47.765 ;
        RECT -15.125 46.075 -14.795 46.405 ;
        RECT -15.125 44.715 -14.795 45.045 ;
        RECT -15.125 43.355 -14.795 43.685 ;
        RECT -15.125 41.995 -14.795 42.325 ;
        RECT -15.125 40.635 -14.795 40.965 ;
        RECT -15.125 39.275 -14.795 39.605 ;
        RECT -15.125 37.915 -14.795 38.245 ;
        RECT -15.125 36.555 -14.795 36.885 ;
        RECT -15.125 35.195 -14.795 35.525 ;
        RECT -15.125 33.835 -14.795 34.165 ;
        RECT -15.125 32.475 -14.795 32.805 ;
        RECT -15.125 31.115 -14.795 31.445 ;
        RECT -15.125 29.755 -14.795 30.085 ;
        RECT -15.125 28.395 -14.795 28.725 ;
        RECT -15.125 27.035 -14.795 27.365 ;
        RECT -15.125 25.675 -14.795 26.005 ;
        RECT -15.125 24.315 -14.795 24.645 ;
        RECT -15.125 22.955 -14.795 23.285 ;
        RECT -15.125 21.595 -14.795 21.925 ;
        RECT -15.125 20.235 -14.795 20.565 ;
        RECT -15.125 18.875 -14.795 19.205 ;
        RECT -15.125 17.515 -14.795 17.845 ;
        RECT -15.125 16.155 -14.795 16.485 ;
        RECT -15.125 14.795 -14.795 15.125 ;
        RECT -15.125 13.435 -14.795 13.765 ;
        RECT -15.125 12.075 -14.795 12.405 ;
        RECT -15.125 10.715 -14.795 11.045 ;
        RECT -15.125 9.355 -14.795 9.685 ;
        RECT -15.125 7.995 -14.795 8.325 ;
        RECT -15.125 6.635 -14.795 6.965 ;
        RECT -15.125 5.275 -14.795 5.605 ;
        RECT -15.125 3.915 -14.795 4.245 ;
        RECT -15.125 2.555 -14.795 2.885 ;
        RECT -15.125 1.195 -14.795 1.525 ;
        RECT -15.125 -0.165 -14.795 0.165 ;
        RECT -15.125 -2.885 -14.795 -2.555 ;
        RECT -15.125 -4.245 -14.795 -3.915 ;
        RECT -15.125 -5.605 -14.795 -5.275 ;
        RECT -15.125 -8.325 -14.795 -7.995 ;
        RECT -15.125 -9.685 -14.795 -9.355 ;
        RECT -15.125 -12.405 -14.795 -12.075 ;
        RECT -15.125 -14.95 -14.795 -14.62 ;
        RECT -15.125 -17.845 -14.795 -17.515 ;
        RECT -15.125 -19.79 -14.795 -19.46 ;
        RECT -15.125 -27.365 -14.795 -27.035 ;
        RECT -15.125 -28.725 -14.795 -28.395 ;
        RECT -15.125 -30.085 -14.795 -29.755 ;
        RECT -15.125 -31.445 -14.795 -31.115 ;
        RECT -15.125 -32.805 -14.795 -32.475 ;
        RECT -15.125 -36.885 -14.795 -36.555 ;
        RECT -15.125 -37.93 -14.795 -37.6 ;
        RECT -15.125 -40.965 -14.795 -40.635 ;
        RECT -15.125 -42.77 -14.795 -42.44 ;
        RECT -15.125 -43.685 -14.795 -43.355 ;
        RECT -15.125 -50.485 -14.795 -50.155 ;
        RECT -15.125 -51.845 -14.795 -51.515 ;
        RECT -15.125 -53.205 -14.795 -52.875 ;
        RECT -15.125 -54.565 -14.795 -54.235 ;
        RECT -15.125 -55.925 -14.795 -55.595 ;
        RECT -15.125 -57.285 -14.795 -56.955 ;
        RECT -15.125 -58.645 -14.795 -58.315 ;
        RECT -15.125 -60.005 -14.795 -59.675 ;
        RECT -15.125 -61.365 -14.795 -61.035 ;
        RECT -15.125 -62.725 -14.795 -62.395 ;
        RECT -15.125 -64.085 -14.795 -63.755 ;
        RECT -15.125 -65.445 -14.795 -65.115 ;
        RECT -15.125 -66.805 -14.795 -66.475 ;
        RECT -15.125 -68.165 -14.795 -67.835 ;
        RECT -15.125 -69.525 -14.795 -69.195 ;
        RECT -15.125 -70.885 -14.795 -70.555 ;
        RECT -15.125 -72.245 -14.795 -71.915 ;
        RECT -15.125 -74.965 -14.795 -74.635 ;
        RECT -15.125 -76.71 -14.795 -76.38 ;
        RECT -15.125 -77.685 -14.795 -77.355 ;
        RECT -15.125 -79.045 -14.795 -78.715 ;
        RECT -15.125 -81.765 -14.795 -81.435 ;
        RECT -15.125 -83.125 -14.795 -82.795 ;
        RECT -15.125 -84.485 -14.795 -84.155 ;
        RECT -15.125 -85.25 -14.795 -84.92 ;
        RECT -15.125 -87.205 -14.795 -86.875 ;
        RECT -15.125 -89.925 -14.795 -89.595 ;
        RECT -15.125 -91.285 -14.795 -90.955 ;
        RECT -15.125 -92.645 -14.795 -92.315 ;
        RECT -15.125 -94.005 -14.795 -93.675 ;
        RECT -15.125 -96.725 -14.795 -96.395 ;
        RECT -15.125 -98.085 -14.795 -97.755 ;
        RECT -15.125 -98.89 -14.795 -98.56 ;
        RECT -15.125 -100.805 -14.795 -100.475 ;
        RECT -15.125 -102.165 -14.795 -101.835 ;
        RECT -15.125 -104.885 -14.795 -104.555 ;
        RECT -15.125 -106.245 -14.795 -105.915 ;
        RECT -15.125 -107.43 -14.795 -107.1 ;
        RECT -15.12 -109.64 -14.8 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -15.125 -114.405 -14.795 -114.075 ;
        RECT -15.125 -115.765 -14.795 -115.435 ;
        RECT -15.125 -117.125 -14.795 -116.795 ;
        RECT -15.125 -121.205 -14.795 -120.875 ;
        RECT -15.125 -125.285 -14.795 -124.955 ;
        RECT -15.125 -128.005 -14.795 -127.675 ;
        RECT -15.125 -133.445 -14.795 -133.115 ;
        RECT -15.125 -136.165 -14.795 -135.835 ;
        RECT -15.125 -138.885 -14.795 -138.555 ;
        RECT -15.125 -141.605 -14.795 -141.275 ;
        RECT -15.125 -145.685 -14.795 -145.355 ;
        RECT -15.125 -147.045 -14.795 -146.715 ;
        RECT -15.125 -152.485 -14.795 -152.155 ;
        RECT -15.125 -156.565 -14.795 -156.235 ;
        RECT -15.125 -157.925 -14.795 -157.595 ;
        RECT -15.125 -159.285 -14.795 -158.955 ;
        RECT -15.125 -160.645 -14.795 -160.315 ;
        RECT -15.125 -162.005 -14.795 -161.675 ;
        RECT -15.125 -163.365 -14.795 -163.035 ;
        RECT -15.125 -164.725 -14.795 -164.395 ;
        RECT -15.125 -166.085 -14.795 -165.755 ;
        RECT -15.125 -167.445 -14.795 -167.115 ;
        RECT -15.125 -170.165 -14.795 -169.835 ;
        RECT -15.12 -172.2 -14.8 -113.4 ;
    END
    PORT
      LAYER met3 ;
        RECT -13.765 105.915 -13.435 106.245 ;
        RECT -13.765 104.555 -13.435 104.885 ;
        RECT -13.765 103.195 -13.435 103.525 ;
        RECT -13.765 101.835 -13.435 102.165 ;
        RECT -13.765 100.475 -13.435 100.805 ;
        RECT -13.765 99.115 -13.435 99.445 ;
        RECT -13.765 97.755 -13.435 98.085 ;
        RECT -13.765 96.395 -13.435 96.725 ;
        RECT -13.765 95.035 -13.435 95.365 ;
        RECT -13.765 93.675 -13.435 94.005 ;
        RECT -13.765 92.315 -13.435 92.645 ;
        RECT -13.765 90.955 -13.435 91.285 ;
        RECT -13.765 89.595 -13.435 89.925 ;
        RECT -13.765 88.235 -13.435 88.565 ;
        RECT -13.765 86.875 -13.435 87.205 ;
        RECT -13.765 85.515 -13.435 85.845 ;
        RECT -13.765 84.155 -13.435 84.485 ;
        RECT -13.765 82.795 -13.435 83.125 ;
        RECT -13.765 81.435 -13.435 81.765 ;
        RECT -13.765 80.075 -13.435 80.405 ;
        RECT -13.765 78.715 -13.435 79.045 ;
        RECT -13.765 77.355 -13.435 77.685 ;
        RECT -13.765 75.995 -13.435 76.325 ;
        RECT -13.765 74.635 -13.435 74.965 ;
        RECT -13.765 73.275 -13.435 73.605 ;
        RECT -13.765 71.915 -13.435 72.245 ;
        RECT -13.765 70.555 -13.435 70.885 ;
        RECT -13.765 69.195 -13.435 69.525 ;
        RECT -13.765 67.835 -13.435 68.165 ;
        RECT -13.765 66.475 -13.435 66.805 ;
        RECT -13.765 65.115 -13.435 65.445 ;
        RECT -13.765 63.755 -13.435 64.085 ;
        RECT -13.765 62.395 -13.435 62.725 ;
        RECT -13.765 61.035 -13.435 61.365 ;
        RECT -13.765 59.675 -13.435 60.005 ;
        RECT -13.765 58.315 -13.435 58.645 ;
        RECT -13.765 56.955 -13.435 57.285 ;
        RECT -13.765 55.595 -13.435 55.925 ;
        RECT -13.765 54.235 -13.435 54.565 ;
        RECT -13.765 52.875 -13.435 53.205 ;
        RECT -13.765 51.515 -13.435 51.845 ;
        RECT -13.765 50.155 -13.435 50.485 ;
        RECT -13.765 48.795 -13.435 49.125 ;
        RECT -13.765 47.435 -13.435 47.765 ;
        RECT -13.765 46.075 -13.435 46.405 ;
        RECT -13.765 44.715 -13.435 45.045 ;
        RECT -13.765 43.355 -13.435 43.685 ;
        RECT -13.765 41.995 -13.435 42.325 ;
        RECT -13.765 40.635 -13.435 40.965 ;
        RECT -13.765 39.275 -13.435 39.605 ;
        RECT -13.765 37.915 -13.435 38.245 ;
        RECT -13.765 36.555 -13.435 36.885 ;
        RECT -13.765 35.195 -13.435 35.525 ;
        RECT -13.765 33.835 -13.435 34.165 ;
        RECT -13.765 32.475 -13.435 32.805 ;
        RECT -13.765 31.115 -13.435 31.445 ;
        RECT -13.765 29.755 -13.435 30.085 ;
        RECT -13.765 28.395 -13.435 28.725 ;
        RECT -13.765 27.035 -13.435 27.365 ;
        RECT -13.765 25.675 -13.435 26.005 ;
        RECT -13.765 24.315 -13.435 24.645 ;
        RECT -13.765 22.955 -13.435 23.285 ;
        RECT -13.765 21.595 -13.435 21.925 ;
        RECT -13.765 20.235 -13.435 20.565 ;
        RECT -13.765 18.875 -13.435 19.205 ;
        RECT -13.765 17.515 -13.435 17.845 ;
        RECT -13.765 16.155 -13.435 16.485 ;
        RECT -13.765 14.795 -13.435 15.125 ;
        RECT -13.765 13.435 -13.435 13.765 ;
        RECT -13.765 12.075 -13.435 12.405 ;
        RECT -13.765 10.715 -13.435 11.045 ;
        RECT -13.765 9.355 -13.435 9.685 ;
        RECT -13.765 7.995 -13.435 8.325 ;
        RECT -13.765 6.635 -13.435 6.965 ;
        RECT -13.765 5.275 -13.435 5.605 ;
        RECT -13.765 3.915 -13.435 4.245 ;
        RECT -13.765 2.555 -13.435 2.885 ;
        RECT -13.765 1.195 -13.435 1.525 ;
        RECT -13.765 -0.165 -13.435 0.165 ;
        RECT -13.765 -2.885 -13.435 -2.555 ;
        RECT -13.765 -4.245 -13.435 -3.915 ;
        RECT -13.765 -5.605 -13.435 -5.275 ;
        RECT -13.765 -8.325 -13.435 -7.995 ;
        RECT -13.765 -9.685 -13.435 -9.355 ;
        RECT -13.765 -12.405 -13.435 -12.075 ;
        RECT -13.765 -14.95 -13.435 -14.62 ;
        RECT -13.765 -17.845 -13.435 -17.515 ;
        RECT -13.765 -19.79 -13.435 -19.46 ;
        RECT -13.765 -27.365 -13.435 -27.035 ;
        RECT -13.765 -28.725 -13.435 -28.395 ;
        RECT -13.765 -30.085 -13.435 -29.755 ;
        RECT -13.765 -31.445 -13.435 -31.115 ;
        RECT -13.765 -32.805 -13.435 -32.475 ;
        RECT -13.765 -36.885 -13.435 -36.555 ;
        RECT -13.765 -37.93 -13.435 -37.6 ;
        RECT -13.765 -40.965 -13.435 -40.635 ;
        RECT -13.765 -42.77 -13.435 -42.44 ;
        RECT -13.765 -43.685 -13.435 -43.355 ;
        RECT -13.765 -50.485 -13.435 -50.155 ;
        RECT -13.765 -51.845 -13.435 -51.515 ;
        RECT -13.765 -53.205 -13.435 -52.875 ;
        RECT -13.765 -54.565 -13.435 -54.235 ;
        RECT -13.765 -55.925 -13.435 -55.595 ;
        RECT -13.765 -57.285 -13.435 -56.955 ;
        RECT -13.765 -58.645 -13.435 -58.315 ;
        RECT -13.765 -60.005 -13.435 -59.675 ;
        RECT -13.765 -61.365 -13.435 -61.035 ;
        RECT -13.765 -62.725 -13.435 -62.395 ;
        RECT -13.765 -64.085 -13.435 -63.755 ;
        RECT -13.765 -65.445 -13.435 -65.115 ;
        RECT -13.765 -66.805 -13.435 -66.475 ;
        RECT -13.765 -68.165 -13.435 -67.835 ;
        RECT -13.765 -69.525 -13.435 -69.195 ;
        RECT -13.765 -70.885 -13.435 -70.555 ;
        RECT -13.765 -72.245 -13.435 -71.915 ;
        RECT -13.765 -74.965 -13.435 -74.635 ;
        RECT -13.765 -76.71 -13.435 -76.38 ;
        RECT -13.765 -77.685 -13.435 -77.355 ;
        RECT -13.765 -79.045 -13.435 -78.715 ;
        RECT -13.765 -81.765 -13.435 -81.435 ;
        RECT -13.765 -83.125 -13.435 -82.795 ;
        RECT -13.765 -84.485 -13.435 -84.155 ;
        RECT -13.765 -85.25 -13.435 -84.92 ;
        RECT -13.765 -87.205 -13.435 -86.875 ;
        RECT -13.765 -89.925 -13.435 -89.595 ;
        RECT -13.765 -91.285 -13.435 -90.955 ;
        RECT -13.765 -92.645 -13.435 -92.315 ;
        RECT -13.765 -94.005 -13.435 -93.675 ;
        RECT -13.765 -96.725 -13.435 -96.395 ;
        RECT -13.765 -98.085 -13.435 -97.755 ;
        RECT -13.765 -98.89 -13.435 -98.56 ;
        RECT -13.765 -100.805 -13.435 -100.475 ;
        RECT -13.765 -102.165 -13.435 -101.835 ;
        RECT -13.765 -104.885 -13.435 -104.555 ;
        RECT -13.765 -106.245 -13.435 -105.915 ;
        RECT -13.765 -107.43 -13.435 -107.1 ;
        RECT -13.765 -113.045 -13.435 -112.715 ;
        RECT -13.765 -114.405 -13.435 -114.075 ;
        RECT -13.765 -115.765 -13.435 -115.435 ;
        RECT -13.765 -117.125 -13.435 -116.795 ;
        RECT -13.765 -119.845 -13.435 -119.515 ;
        RECT -13.765 -121.205 -13.435 -120.875 ;
        RECT -13.765 -125.285 -13.435 -124.955 ;
        RECT -13.765 -129.365 -13.435 -129.035 ;
        RECT -13.765 -133.445 -13.435 -133.115 ;
        RECT -13.765 -136.165 -13.435 -135.835 ;
        RECT -13.765 -138.885 -13.435 -138.555 ;
        RECT -13.765 -141.605 -13.435 -141.275 ;
        RECT -13.765 -145.685 -13.435 -145.355 ;
        RECT -13.765 -147.045 -13.435 -146.715 ;
        RECT -13.765 -149.765 -13.435 -149.435 ;
        RECT -13.765 -152.485 -13.435 -152.155 ;
        RECT -13.765 -156.565 -13.435 -156.235 ;
        RECT -13.765 -157.925 -13.435 -157.595 ;
        RECT -13.765 -159.285 -13.435 -158.955 ;
        RECT -13.765 -160.645 -13.435 -160.315 ;
        RECT -13.765 -162.005 -13.435 -161.675 ;
        RECT -13.765 -163.365 -13.435 -163.035 ;
        RECT -13.765 -164.725 -13.435 -164.395 ;
        RECT -13.765 -166.085 -13.435 -165.755 ;
        RECT -13.765 -170.165 -13.435 -169.835 ;
        RECT -13.765 -172.885 -13.435 -172.555 ;
        RECT -13.765 -174.245 -13.435 -173.915 ;
        RECT -13.765 -175.725 -13.435 -175.395 ;
        RECT -13.765 -176.965 -13.435 -176.635 ;
        RECT -13.765 -178.325 -13.435 -177.995 ;
        RECT -13.765 -180.57 -13.435 -179.44 ;
        RECT -13.76 -180.685 -13.44 242.565 ;
        RECT -13.765 241.32 -13.435 242.45 ;
        RECT -13.765 239.195 -13.435 239.525 ;
        RECT -13.765 237.835 -13.435 238.165 ;
        RECT -13.765 236.475 -13.435 236.805 ;
        RECT -13.765 235.115 -13.435 235.445 ;
        RECT -13.765 233.755 -13.435 234.085 ;
        RECT -13.765 232.395 -13.435 232.725 ;
        RECT -13.765 231.035 -13.435 231.365 ;
        RECT -13.765 229.675 -13.435 230.005 ;
        RECT -13.765 228.315 -13.435 228.645 ;
        RECT -13.765 226.955 -13.435 227.285 ;
        RECT -13.765 225.595 -13.435 225.925 ;
        RECT -13.765 224.235 -13.435 224.565 ;
        RECT -13.765 222.875 -13.435 223.205 ;
        RECT -13.765 221.515 -13.435 221.845 ;
        RECT -13.765 220.155 -13.435 220.485 ;
        RECT -13.765 218.795 -13.435 219.125 ;
        RECT -13.765 217.435 -13.435 217.765 ;
        RECT -13.765 216.075 -13.435 216.405 ;
        RECT -13.765 214.715 -13.435 215.045 ;
        RECT -13.765 213.355 -13.435 213.685 ;
        RECT -13.765 211.995 -13.435 212.325 ;
        RECT -13.765 210.635 -13.435 210.965 ;
        RECT -13.765 209.275 -13.435 209.605 ;
        RECT -13.765 207.915 -13.435 208.245 ;
        RECT -13.765 206.555 -13.435 206.885 ;
        RECT -13.765 205.195 -13.435 205.525 ;
        RECT -13.765 203.835 -13.435 204.165 ;
        RECT -13.765 202.475 -13.435 202.805 ;
        RECT -13.765 201.115 -13.435 201.445 ;
        RECT -13.765 199.755 -13.435 200.085 ;
        RECT -13.765 198.395 -13.435 198.725 ;
        RECT -13.765 197.035 -13.435 197.365 ;
        RECT -13.765 195.675 -13.435 196.005 ;
        RECT -13.765 194.315 -13.435 194.645 ;
        RECT -13.765 192.955 -13.435 193.285 ;
        RECT -13.765 191.595 -13.435 191.925 ;
        RECT -13.765 190.235 -13.435 190.565 ;
        RECT -13.765 188.875 -13.435 189.205 ;
        RECT -13.765 187.515 -13.435 187.845 ;
        RECT -13.765 186.155 -13.435 186.485 ;
        RECT -13.765 184.795 -13.435 185.125 ;
        RECT -13.765 183.435 -13.435 183.765 ;
        RECT -13.765 182.075 -13.435 182.405 ;
        RECT -13.765 180.715 -13.435 181.045 ;
        RECT -13.765 179.355 -13.435 179.685 ;
        RECT -13.765 177.995 -13.435 178.325 ;
        RECT -13.765 176.635 -13.435 176.965 ;
        RECT -13.765 175.275 -13.435 175.605 ;
        RECT -13.765 173.915 -13.435 174.245 ;
        RECT -13.765 172.555 -13.435 172.885 ;
        RECT -13.765 171.195 -13.435 171.525 ;
        RECT -13.765 169.835 -13.435 170.165 ;
        RECT -13.765 168.475 -13.435 168.805 ;
        RECT -13.765 167.115 -13.435 167.445 ;
        RECT -13.765 165.755 -13.435 166.085 ;
        RECT -13.765 164.395 -13.435 164.725 ;
        RECT -13.765 163.035 -13.435 163.365 ;
        RECT -13.765 161.675 -13.435 162.005 ;
        RECT -13.765 160.315 -13.435 160.645 ;
        RECT -13.765 158.955 -13.435 159.285 ;
        RECT -13.765 157.595 -13.435 157.925 ;
        RECT -13.765 156.235 -13.435 156.565 ;
        RECT -13.765 154.875 -13.435 155.205 ;
        RECT -13.765 153.515 -13.435 153.845 ;
        RECT -13.765 152.155 -13.435 152.485 ;
        RECT -13.765 150.795 -13.435 151.125 ;
        RECT -13.765 149.435 -13.435 149.765 ;
        RECT -13.765 148.075 -13.435 148.405 ;
        RECT -13.765 146.715 -13.435 147.045 ;
        RECT -13.765 145.355 -13.435 145.685 ;
        RECT -13.765 143.995 -13.435 144.325 ;
        RECT -13.765 142.635 -13.435 142.965 ;
        RECT -13.765 141.275 -13.435 141.605 ;
        RECT -13.765 139.915 -13.435 140.245 ;
        RECT -13.765 138.555 -13.435 138.885 ;
        RECT -13.765 137.195 -13.435 137.525 ;
        RECT -13.765 135.835 -13.435 136.165 ;
        RECT -13.765 134.475 -13.435 134.805 ;
        RECT -13.765 133.115 -13.435 133.445 ;
        RECT -13.765 131.755 -13.435 132.085 ;
        RECT -13.765 130.395 -13.435 130.725 ;
        RECT -13.765 129.035 -13.435 129.365 ;
        RECT -13.765 127.675 -13.435 128.005 ;
        RECT -13.765 126.315 -13.435 126.645 ;
        RECT -13.765 124.955 -13.435 125.285 ;
        RECT -13.765 123.595 -13.435 123.925 ;
        RECT -13.765 122.235 -13.435 122.565 ;
        RECT -13.765 120.875 -13.435 121.205 ;
        RECT -13.765 119.515 -13.435 119.845 ;
        RECT -13.765 118.155 -13.435 118.485 ;
        RECT -13.765 116.795 -13.435 117.125 ;
        RECT -13.765 115.435 -13.435 115.765 ;
        RECT -13.765 114.075 -13.435 114.405 ;
        RECT -13.765 112.715 -13.435 113.045 ;
        RECT -13.765 111.355 -13.435 111.685 ;
        RECT -13.765 109.995 -13.435 110.325 ;
        RECT -13.765 108.635 -13.435 108.965 ;
        RECT -13.765 107.275 -13.435 107.605 ;
    END
    PORT
      LAYER met3 ;
        RECT -23.285 241.32 -22.955 242.45 ;
        RECT -23.285 239.195 -22.955 239.525 ;
        RECT -23.285 237.835 -22.955 238.165 ;
        RECT -23.285 236.475 -22.955 236.805 ;
        RECT -23.285 235.115 -22.955 235.445 ;
        RECT -23.285 233.755 -22.955 234.085 ;
        RECT -23.285 232.395 -22.955 232.725 ;
        RECT -23.285 231.035 -22.955 231.365 ;
        RECT -23.285 229.675 -22.955 230.005 ;
        RECT -23.285 228.315 -22.955 228.645 ;
        RECT -23.285 226.955 -22.955 227.285 ;
        RECT -23.285 225.595 -22.955 225.925 ;
        RECT -23.285 224.235 -22.955 224.565 ;
        RECT -23.285 222.875 -22.955 223.205 ;
        RECT -23.285 221.515 -22.955 221.845 ;
        RECT -23.285 220.155 -22.955 220.485 ;
        RECT -23.285 218.795 -22.955 219.125 ;
        RECT -23.285 217.435 -22.955 217.765 ;
        RECT -23.285 216.075 -22.955 216.405 ;
        RECT -23.285 214.715 -22.955 215.045 ;
        RECT -23.285 213.355 -22.955 213.685 ;
        RECT -23.285 211.995 -22.955 212.325 ;
        RECT -23.285 210.635 -22.955 210.965 ;
        RECT -23.285 209.275 -22.955 209.605 ;
        RECT -23.285 207.915 -22.955 208.245 ;
        RECT -23.285 206.555 -22.955 206.885 ;
        RECT -23.285 205.195 -22.955 205.525 ;
        RECT -23.285 203.835 -22.955 204.165 ;
        RECT -23.285 202.475 -22.955 202.805 ;
        RECT -23.285 201.115 -22.955 201.445 ;
        RECT -23.285 199.755 -22.955 200.085 ;
        RECT -23.285 198.395 -22.955 198.725 ;
        RECT -23.285 197.035 -22.955 197.365 ;
        RECT -23.285 195.675 -22.955 196.005 ;
        RECT -23.285 194.315 -22.955 194.645 ;
        RECT -23.285 192.955 -22.955 193.285 ;
        RECT -23.285 191.595 -22.955 191.925 ;
        RECT -23.285 190.235 -22.955 190.565 ;
        RECT -23.285 188.875 -22.955 189.205 ;
        RECT -23.285 187.515 -22.955 187.845 ;
        RECT -23.285 186.155 -22.955 186.485 ;
        RECT -23.285 184.795 -22.955 185.125 ;
        RECT -23.285 183.435 -22.955 183.765 ;
        RECT -23.285 182.075 -22.955 182.405 ;
        RECT -23.285 180.715 -22.955 181.045 ;
        RECT -23.285 179.355 -22.955 179.685 ;
        RECT -23.285 177.995 -22.955 178.325 ;
        RECT -23.285 176.635 -22.955 176.965 ;
        RECT -23.285 175.275 -22.955 175.605 ;
        RECT -23.285 173.915 -22.955 174.245 ;
        RECT -23.285 172.555 -22.955 172.885 ;
        RECT -23.285 171.195 -22.955 171.525 ;
        RECT -23.285 169.835 -22.955 170.165 ;
        RECT -23.285 168.475 -22.955 168.805 ;
        RECT -23.285 167.115 -22.955 167.445 ;
        RECT -23.285 165.755 -22.955 166.085 ;
        RECT -23.285 164.395 -22.955 164.725 ;
        RECT -23.285 163.035 -22.955 163.365 ;
        RECT -23.285 161.675 -22.955 162.005 ;
        RECT -23.285 160.315 -22.955 160.645 ;
        RECT -23.285 158.955 -22.955 159.285 ;
        RECT -23.285 157.595 -22.955 157.925 ;
        RECT -23.285 156.235 -22.955 156.565 ;
        RECT -23.285 154.875 -22.955 155.205 ;
        RECT -23.285 153.515 -22.955 153.845 ;
        RECT -23.285 152.155 -22.955 152.485 ;
        RECT -23.285 150.795 -22.955 151.125 ;
        RECT -23.285 149.435 -22.955 149.765 ;
        RECT -23.285 148.075 -22.955 148.405 ;
        RECT -23.285 146.715 -22.955 147.045 ;
        RECT -23.285 145.355 -22.955 145.685 ;
        RECT -23.285 143.995 -22.955 144.325 ;
        RECT -23.285 142.635 -22.955 142.965 ;
        RECT -23.285 141.275 -22.955 141.605 ;
        RECT -23.285 139.915 -22.955 140.245 ;
        RECT -23.285 138.555 -22.955 138.885 ;
        RECT -23.285 137.195 -22.955 137.525 ;
        RECT -23.285 135.835 -22.955 136.165 ;
        RECT -23.285 134.475 -22.955 134.805 ;
        RECT -23.285 133.115 -22.955 133.445 ;
        RECT -23.285 131.755 -22.955 132.085 ;
        RECT -23.285 130.395 -22.955 130.725 ;
        RECT -23.285 129.035 -22.955 129.365 ;
        RECT -23.285 127.675 -22.955 128.005 ;
        RECT -23.285 126.315 -22.955 126.645 ;
        RECT -23.285 124.955 -22.955 125.285 ;
        RECT -23.285 123.595 -22.955 123.925 ;
        RECT -23.285 122.235 -22.955 122.565 ;
        RECT -23.285 120.875 -22.955 121.205 ;
        RECT -23.285 119.515 -22.955 119.845 ;
        RECT -23.285 118.155 -22.955 118.485 ;
        RECT -23.285 116.795 -22.955 117.125 ;
        RECT -23.285 115.435 -22.955 115.765 ;
        RECT -23.285 114.075 -22.955 114.405 ;
        RECT -23.285 112.715 -22.955 113.045 ;
        RECT -23.285 111.355 -22.955 111.685 ;
        RECT -23.285 109.995 -22.955 110.325 ;
        RECT -23.285 108.635 -22.955 108.965 ;
        RECT -23.285 107.275 -22.955 107.605 ;
        RECT -23.285 105.915 -22.955 106.245 ;
        RECT -23.285 104.555 -22.955 104.885 ;
        RECT -23.285 103.195 -22.955 103.525 ;
        RECT -23.285 101.835 -22.955 102.165 ;
        RECT -23.285 100.475 -22.955 100.805 ;
        RECT -23.285 99.115 -22.955 99.445 ;
        RECT -23.285 97.755 -22.955 98.085 ;
        RECT -23.285 96.395 -22.955 96.725 ;
        RECT -23.285 95.035 -22.955 95.365 ;
        RECT -23.285 93.675 -22.955 94.005 ;
        RECT -23.285 92.315 -22.955 92.645 ;
        RECT -23.285 90.955 -22.955 91.285 ;
        RECT -23.285 89.595 -22.955 89.925 ;
        RECT -23.285 88.235 -22.955 88.565 ;
        RECT -23.285 86.875 -22.955 87.205 ;
        RECT -23.285 85.515 -22.955 85.845 ;
        RECT -23.285 84.155 -22.955 84.485 ;
        RECT -23.285 82.795 -22.955 83.125 ;
        RECT -23.285 81.435 -22.955 81.765 ;
        RECT -23.285 80.075 -22.955 80.405 ;
        RECT -23.285 78.715 -22.955 79.045 ;
        RECT -23.285 77.355 -22.955 77.685 ;
        RECT -23.285 75.995 -22.955 76.325 ;
        RECT -23.285 74.635 -22.955 74.965 ;
        RECT -23.285 73.275 -22.955 73.605 ;
        RECT -23.285 71.915 -22.955 72.245 ;
        RECT -23.285 70.555 -22.955 70.885 ;
        RECT -23.285 69.195 -22.955 69.525 ;
        RECT -23.285 67.835 -22.955 68.165 ;
        RECT -23.285 66.475 -22.955 66.805 ;
        RECT -23.285 65.115 -22.955 65.445 ;
        RECT -23.285 63.755 -22.955 64.085 ;
        RECT -23.285 62.395 -22.955 62.725 ;
        RECT -23.285 61.035 -22.955 61.365 ;
        RECT -23.285 59.675 -22.955 60.005 ;
        RECT -23.285 58.315 -22.955 58.645 ;
        RECT -23.285 56.955 -22.955 57.285 ;
        RECT -23.285 55.595 -22.955 55.925 ;
        RECT -23.285 54.235 -22.955 54.565 ;
        RECT -23.285 52.875 -22.955 53.205 ;
        RECT -23.285 51.515 -22.955 51.845 ;
        RECT -23.285 50.155 -22.955 50.485 ;
        RECT -23.285 48.795 -22.955 49.125 ;
        RECT -23.285 47.435 -22.955 47.765 ;
        RECT -23.285 46.075 -22.955 46.405 ;
        RECT -23.285 44.715 -22.955 45.045 ;
        RECT -23.285 43.355 -22.955 43.685 ;
        RECT -23.285 41.995 -22.955 42.325 ;
        RECT -23.285 40.635 -22.955 40.965 ;
        RECT -23.285 39.275 -22.955 39.605 ;
        RECT -23.285 37.915 -22.955 38.245 ;
        RECT -23.285 36.555 -22.955 36.885 ;
        RECT -23.285 35.195 -22.955 35.525 ;
        RECT -23.285 33.835 -22.955 34.165 ;
        RECT -23.285 32.475 -22.955 32.805 ;
        RECT -23.285 31.115 -22.955 31.445 ;
        RECT -23.285 29.755 -22.955 30.085 ;
        RECT -23.285 28.395 -22.955 28.725 ;
        RECT -23.285 27.035 -22.955 27.365 ;
        RECT -23.285 25.675 -22.955 26.005 ;
        RECT -23.285 24.315 -22.955 24.645 ;
        RECT -23.285 22.955 -22.955 23.285 ;
        RECT -23.285 21.595 -22.955 21.925 ;
        RECT -23.285 20.235 -22.955 20.565 ;
        RECT -23.285 18.875 -22.955 19.205 ;
        RECT -23.285 17.515 -22.955 17.845 ;
        RECT -23.285 16.155 -22.955 16.485 ;
        RECT -23.285 14.795 -22.955 15.125 ;
        RECT -23.285 13.435 -22.955 13.765 ;
        RECT -23.285 12.075 -22.955 12.405 ;
        RECT -23.285 10.715 -22.955 11.045 ;
        RECT -23.285 9.355 -22.955 9.685 ;
        RECT -23.285 7.995 -22.955 8.325 ;
        RECT -23.285 6.635 -22.955 6.965 ;
        RECT -23.285 5.275 -22.955 5.605 ;
        RECT -23.285 3.915 -22.955 4.245 ;
        RECT -23.285 2.555 -22.955 2.885 ;
        RECT -23.285 1.195 -22.955 1.525 ;
        RECT -23.285 -0.165 -22.955 0.165 ;
        RECT -23.285 -2.885 -22.955 -2.555 ;
        RECT -23.285 -8.325 -22.955 -7.995 ;
        RECT -23.285 -9.685 -22.955 -9.355 ;
        RECT -23.285 -14.95 -22.955 -14.62 ;
        RECT -23.285 -17.845 -22.955 -17.515 ;
        RECT -23.285 -19.79 -22.955 -19.46 ;
        RECT -23.285 -20.565 -22.955 -20.235 ;
        RECT -23.285 -28.725 -22.955 -28.395 ;
        RECT -23.285 -31.445 -22.955 -31.115 ;
        RECT -23.285 -32.805 -22.955 -32.475 ;
        RECT -23.285 -35.525 -22.955 -35.195 ;
        RECT -23.285 -36.885 -22.955 -36.555 ;
        RECT -23.285 -37.93 -22.955 -37.6 ;
        RECT -23.285 -40.965 -22.955 -40.635 ;
        RECT -23.285 -42.77 -22.955 -42.44 ;
        RECT -23.285 -43.685 -22.955 -43.355 ;
        RECT -23.285 -50.485 -22.955 -50.155 ;
        RECT -23.285 -51.845 -22.955 -51.515 ;
        RECT -23.285 -53.205 -22.955 -52.875 ;
        RECT -23.285 -54.565 -22.955 -54.235 ;
        RECT -23.285 -55.925 -22.955 -55.595 ;
        RECT -23.285 -57.285 -22.955 -56.955 ;
        RECT -23.285 -58.645 -22.955 -58.315 ;
        RECT -23.285 -60.005 -22.955 -59.675 ;
        RECT -23.285 -61.365 -22.955 -61.035 ;
        RECT -23.285 -64.085 -22.955 -63.755 ;
        RECT -23.285 -65.445 -22.955 -65.115 ;
        RECT -23.285 -66.805 -22.955 -66.475 ;
        RECT -23.285 -68.165 -22.955 -67.835 ;
        RECT -23.285 -69.525 -22.955 -69.195 ;
        RECT -23.285 -70.885 -22.955 -70.555 ;
        RECT -23.285 -72.245 -22.955 -71.915 ;
        RECT -23.285 -73.605 -22.955 -73.275 ;
        RECT -23.285 -74.965 -22.955 -74.635 ;
        RECT -23.285 -76.325 -22.955 -75.995 ;
        RECT -23.285 -77.685 -22.955 -77.355 ;
        RECT -23.285 -79.045 -22.955 -78.715 ;
        RECT -23.285 -80.405 -22.955 -80.075 ;
        RECT -23.285 -81.765 -22.955 -81.435 ;
        RECT -23.285 -83.125 -22.955 -82.795 ;
        RECT -23.285 -84.485 -22.955 -84.155 ;
        RECT -23.285 -85.845 -22.955 -85.515 ;
        RECT -23.285 -87.205 -22.955 -86.875 ;
        RECT -23.285 -88.565 -22.955 -88.235 ;
        RECT -23.285 -89.925 -22.955 -89.595 ;
        RECT -23.285 -91.285 -22.955 -90.955 ;
        RECT -23.285 -92.645 -22.955 -92.315 ;
        RECT -23.285 -94.005 -22.955 -93.675 ;
        RECT -23.285 -95.365 -22.955 -95.035 ;
        RECT -23.285 -96.725 -22.955 -96.395 ;
        RECT -23.285 -98.085 -22.955 -97.755 ;
        RECT -23.285 -99.445 -22.955 -99.115 ;
        RECT -23.285 -100.805 -22.955 -100.475 ;
        RECT -23.285 -102.165 -22.955 -101.835 ;
        RECT -23.285 -103.525 -22.955 -103.195 ;
        RECT -23.285 -104.885 -22.955 -104.555 ;
        RECT -23.285 -106.245 -22.955 -105.915 ;
        RECT -23.285 -107.605 -22.955 -107.275 ;
        RECT -23.285 -108.965 -22.955 -108.635 ;
        RECT -23.285 -111.685 -22.955 -111.355 ;
        RECT -23.28 -111.685 -22.96 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -23.285 -174.245 -22.955 -173.915 ;
        RECT -23.285 -175.725 -22.955 -175.395 ;
        RECT -23.285 -176.965 -22.955 -176.635 ;
        RECT -23.285 -178.325 -22.955 -177.995 ;
        RECT -23.285 -180.57 -22.955 -179.44 ;
        RECT -23.28 -180.685 -22.96 -172.56 ;
    END
    PORT
      LAYER met3 ;
        RECT -21.925 241.32 -21.595 242.45 ;
        RECT -21.925 239.195 -21.595 239.525 ;
        RECT -21.925 237.835 -21.595 238.165 ;
        RECT -21.925 236.475 -21.595 236.805 ;
        RECT -21.925 235.115 -21.595 235.445 ;
        RECT -21.925 233.755 -21.595 234.085 ;
        RECT -21.925 232.395 -21.595 232.725 ;
        RECT -21.925 231.035 -21.595 231.365 ;
        RECT -21.925 229.675 -21.595 230.005 ;
        RECT -21.925 228.315 -21.595 228.645 ;
        RECT -21.925 226.955 -21.595 227.285 ;
        RECT -21.925 225.595 -21.595 225.925 ;
        RECT -21.925 224.235 -21.595 224.565 ;
        RECT -21.925 222.875 -21.595 223.205 ;
        RECT -21.925 221.515 -21.595 221.845 ;
        RECT -21.925 220.155 -21.595 220.485 ;
        RECT -21.925 218.795 -21.595 219.125 ;
        RECT -21.925 217.435 -21.595 217.765 ;
        RECT -21.925 216.075 -21.595 216.405 ;
        RECT -21.925 214.715 -21.595 215.045 ;
        RECT -21.925 213.355 -21.595 213.685 ;
        RECT -21.925 211.995 -21.595 212.325 ;
        RECT -21.925 210.635 -21.595 210.965 ;
        RECT -21.925 209.275 -21.595 209.605 ;
        RECT -21.925 207.915 -21.595 208.245 ;
        RECT -21.925 206.555 -21.595 206.885 ;
        RECT -21.925 205.195 -21.595 205.525 ;
        RECT -21.925 203.835 -21.595 204.165 ;
        RECT -21.925 202.475 -21.595 202.805 ;
        RECT -21.925 201.115 -21.595 201.445 ;
        RECT -21.925 199.755 -21.595 200.085 ;
        RECT -21.925 198.395 -21.595 198.725 ;
        RECT -21.925 197.035 -21.595 197.365 ;
        RECT -21.925 195.675 -21.595 196.005 ;
        RECT -21.925 194.315 -21.595 194.645 ;
        RECT -21.925 192.955 -21.595 193.285 ;
        RECT -21.925 191.595 -21.595 191.925 ;
        RECT -21.925 190.235 -21.595 190.565 ;
        RECT -21.925 188.875 -21.595 189.205 ;
        RECT -21.925 187.515 -21.595 187.845 ;
        RECT -21.925 186.155 -21.595 186.485 ;
        RECT -21.925 184.795 -21.595 185.125 ;
        RECT -21.925 183.435 -21.595 183.765 ;
        RECT -21.925 182.075 -21.595 182.405 ;
        RECT -21.925 180.715 -21.595 181.045 ;
        RECT -21.925 179.355 -21.595 179.685 ;
        RECT -21.925 177.995 -21.595 178.325 ;
        RECT -21.925 176.635 -21.595 176.965 ;
        RECT -21.925 175.275 -21.595 175.605 ;
        RECT -21.925 173.915 -21.595 174.245 ;
        RECT -21.925 172.555 -21.595 172.885 ;
        RECT -21.925 171.195 -21.595 171.525 ;
        RECT -21.925 169.835 -21.595 170.165 ;
        RECT -21.925 168.475 -21.595 168.805 ;
        RECT -21.925 167.115 -21.595 167.445 ;
        RECT -21.925 165.755 -21.595 166.085 ;
        RECT -21.925 164.395 -21.595 164.725 ;
        RECT -21.925 163.035 -21.595 163.365 ;
        RECT -21.925 161.675 -21.595 162.005 ;
        RECT -21.925 160.315 -21.595 160.645 ;
        RECT -21.925 158.955 -21.595 159.285 ;
        RECT -21.925 157.595 -21.595 157.925 ;
        RECT -21.925 156.235 -21.595 156.565 ;
        RECT -21.925 154.875 -21.595 155.205 ;
        RECT -21.925 153.515 -21.595 153.845 ;
        RECT -21.925 152.155 -21.595 152.485 ;
        RECT -21.925 150.795 -21.595 151.125 ;
        RECT -21.925 149.435 -21.595 149.765 ;
        RECT -21.925 148.075 -21.595 148.405 ;
        RECT -21.925 146.715 -21.595 147.045 ;
        RECT -21.925 145.355 -21.595 145.685 ;
        RECT -21.925 143.995 -21.595 144.325 ;
        RECT -21.925 142.635 -21.595 142.965 ;
        RECT -21.925 141.275 -21.595 141.605 ;
        RECT -21.925 139.915 -21.595 140.245 ;
        RECT -21.925 138.555 -21.595 138.885 ;
        RECT -21.925 137.195 -21.595 137.525 ;
        RECT -21.925 135.835 -21.595 136.165 ;
        RECT -21.925 134.475 -21.595 134.805 ;
        RECT -21.925 133.115 -21.595 133.445 ;
        RECT -21.925 131.755 -21.595 132.085 ;
        RECT -21.925 130.395 -21.595 130.725 ;
        RECT -21.925 129.035 -21.595 129.365 ;
        RECT -21.925 127.675 -21.595 128.005 ;
        RECT -21.925 126.315 -21.595 126.645 ;
        RECT -21.925 124.955 -21.595 125.285 ;
        RECT -21.925 123.595 -21.595 123.925 ;
        RECT -21.925 122.235 -21.595 122.565 ;
        RECT -21.925 120.875 -21.595 121.205 ;
        RECT -21.925 119.515 -21.595 119.845 ;
        RECT -21.925 118.155 -21.595 118.485 ;
        RECT -21.925 116.795 -21.595 117.125 ;
        RECT -21.925 115.435 -21.595 115.765 ;
        RECT -21.925 114.075 -21.595 114.405 ;
        RECT -21.925 112.715 -21.595 113.045 ;
        RECT -21.925 111.355 -21.595 111.685 ;
        RECT -21.925 109.995 -21.595 110.325 ;
        RECT -21.925 108.635 -21.595 108.965 ;
        RECT -21.925 107.275 -21.595 107.605 ;
        RECT -21.925 105.915 -21.595 106.245 ;
        RECT -21.925 104.555 -21.595 104.885 ;
        RECT -21.925 103.195 -21.595 103.525 ;
        RECT -21.925 101.835 -21.595 102.165 ;
        RECT -21.925 100.475 -21.595 100.805 ;
        RECT -21.925 99.115 -21.595 99.445 ;
        RECT -21.925 97.755 -21.595 98.085 ;
        RECT -21.925 96.395 -21.595 96.725 ;
        RECT -21.925 95.035 -21.595 95.365 ;
        RECT -21.925 93.675 -21.595 94.005 ;
        RECT -21.925 92.315 -21.595 92.645 ;
        RECT -21.925 90.955 -21.595 91.285 ;
        RECT -21.925 89.595 -21.595 89.925 ;
        RECT -21.925 88.235 -21.595 88.565 ;
        RECT -21.925 86.875 -21.595 87.205 ;
        RECT -21.925 85.515 -21.595 85.845 ;
        RECT -21.925 84.155 -21.595 84.485 ;
        RECT -21.925 82.795 -21.595 83.125 ;
        RECT -21.925 81.435 -21.595 81.765 ;
        RECT -21.925 80.075 -21.595 80.405 ;
        RECT -21.925 78.715 -21.595 79.045 ;
        RECT -21.925 77.355 -21.595 77.685 ;
        RECT -21.925 75.995 -21.595 76.325 ;
        RECT -21.925 74.635 -21.595 74.965 ;
        RECT -21.925 73.275 -21.595 73.605 ;
        RECT -21.925 71.915 -21.595 72.245 ;
        RECT -21.925 70.555 -21.595 70.885 ;
        RECT -21.925 69.195 -21.595 69.525 ;
        RECT -21.925 67.835 -21.595 68.165 ;
        RECT -21.925 66.475 -21.595 66.805 ;
        RECT -21.925 65.115 -21.595 65.445 ;
        RECT -21.925 63.755 -21.595 64.085 ;
        RECT -21.925 62.395 -21.595 62.725 ;
        RECT -21.925 61.035 -21.595 61.365 ;
        RECT -21.925 59.675 -21.595 60.005 ;
        RECT -21.925 58.315 -21.595 58.645 ;
        RECT -21.925 56.955 -21.595 57.285 ;
        RECT -21.925 55.595 -21.595 55.925 ;
        RECT -21.925 54.235 -21.595 54.565 ;
        RECT -21.925 52.875 -21.595 53.205 ;
        RECT -21.925 51.515 -21.595 51.845 ;
        RECT -21.925 50.155 -21.595 50.485 ;
        RECT -21.925 48.795 -21.595 49.125 ;
        RECT -21.925 47.435 -21.595 47.765 ;
        RECT -21.925 46.075 -21.595 46.405 ;
        RECT -21.925 44.715 -21.595 45.045 ;
        RECT -21.925 43.355 -21.595 43.685 ;
        RECT -21.925 41.995 -21.595 42.325 ;
        RECT -21.925 40.635 -21.595 40.965 ;
        RECT -21.925 39.275 -21.595 39.605 ;
        RECT -21.925 37.915 -21.595 38.245 ;
        RECT -21.925 36.555 -21.595 36.885 ;
        RECT -21.925 35.195 -21.595 35.525 ;
        RECT -21.925 33.835 -21.595 34.165 ;
        RECT -21.925 32.475 -21.595 32.805 ;
        RECT -21.925 31.115 -21.595 31.445 ;
        RECT -21.925 29.755 -21.595 30.085 ;
        RECT -21.925 28.395 -21.595 28.725 ;
        RECT -21.925 27.035 -21.595 27.365 ;
        RECT -21.925 25.675 -21.595 26.005 ;
        RECT -21.925 24.315 -21.595 24.645 ;
        RECT -21.925 22.955 -21.595 23.285 ;
        RECT -21.925 21.595 -21.595 21.925 ;
        RECT -21.925 20.235 -21.595 20.565 ;
        RECT -21.925 18.875 -21.595 19.205 ;
        RECT -21.925 17.515 -21.595 17.845 ;
        RECT -21.925 16.155 -21.595 16.485 ;
        RECT -21.925 14.795 -21.595 15.125 ;
        RECT -21.925 13.435 -21.595 13.765 ;
        RECT -21.925 12.075 -21.595 12.405 ;
        RECT -21.925 10.715 -21.595 11.045 ;
        RECT -21.925 9.355 -21.595 9.685 ;
        RECT -21.925 7.995 -21.595 8.325 ;
        RECT -21.925 6.635 -21.595 6.965 ;
        RECT -21.925 5.275 -21.595 5.605 ;
        RECT -21.925 3.915 -21.595 4.245 ;
        RECT -21.925 2.555 -21.595 2.885 ;
        RECT -21.925 1.195 -21.595 1.525 ;
        RECT -21.925 -0.165 -21.595 0.165 ;
        RECT -21.925 -2.885 -21.595 -2.555 ;
        RECT -21.925 -8.325 -21.595 -7.995 ;
        RECT -21.925 -9.685 -21.595 -9.355 ;
        RECT -21.925 -14.95 -21.595 -14.62 ;
        RECT -21.925 -17.845 -21.595 -17.515 ;
        RECT -21.925 -19.79 -21.595 -19.46 ;
        RECT -21.925 -20.565 -21.595 -20.235 ;
        RECT -21.92 -23.96 -21.6 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -21.925 -64.085 -21.595 -63.755 ;
        RECT -21.925 -65.445 -21.595 -65.115 ;
        RECT -21.925 -66.805 -21.595 -66.475 ;
        RECT -21.925 -68.165 -21.595 -67.835 ;
        RECT -21.925 -69.525 -21.595 -69.195 ;
        RECT -21.925 -70.885 -21.595 -70.555 ;
        RECT -21.925 -72.245 -21.595 -71.915 ;
        RECT -21.925 -73.605 -21.595 -73.275 ;
        RECT -21.925 -74.965 -21.595 -74.635 ;
        RECT -21.925 -76.325 -21.595 -75.995 ;
        RECT -21.925 -77.685 -21.595 -77.355 ;
        RECT -21.925 -79.045 -21.595 -78.715 ;
        RECT -21.925 -80.405 -21.595 -80.075 ;
        RECT -21.925 -81.765 -21.595 -81.435 ;
        RECT -21.925 -83.125 -21.595 -82.795 ;
        RECT -21.925 -84.485 -21.595 -84.155 ;
        RECT -21.925 -85.845 -21.595 -85.515 ;
        RECT -21.925 -87.205 -21.595 -86.875 ;
        RECT -21.925 -88.565 -21.595 -88.235 ;
        RECT -21.925 -89.925 -21.595 -89.595 ;
        RECT -21.925 -91.285 -21.595 -90.955 ;
        RECT -21.925 -92.645 -21.595 -92.315 ;
        RECT -21.925 -94.005 -21.595 -93.675 ;
        RECT -21.925 -95.365 -21.595 -95.035 ;
        RECT -21.925 -96.725 -21.595 -96.395 ;
        RECT -21.925 -98.085 -21.595 -97.755 ;
        RECT -21.925 -99.445 -21.595 -99.115 ;
        RECT -21.925 -100.805 -21.595 -100.475 ;
        RECT -21.925 -102.165 -21.595 -101.835 ;
        RECT -21.925 -103.525 -21.595 -103.195 ;
        RECT -21.925 -104.885 -21.595 -104.555 ;
        RECT -21.925 -106.245 -21.595 -105.915 ;
        RECT -21.925 -107.605 -21.595 -107.275 ;
        RECT -21.925 -108.965 -21.595 -108.635 ;
        RECT -21.925 -111.685 -21.595 -111.355 ;
        RECT -21.925 -113.045 -21.595 -112.715 ;
        RECT -21.925 -114.405 -21.595 -114.075 ;
        RECT -21.925 -115.765 -21.595 -115.435 ;
        RECT -21.925 -117.125 -21.595 -116.795 ;
        RECT -21.925 -118.485 -21.595 -118.155 ;
        RECT -21.925 -122.565 -21.595 -122.235 ;
        RECT -21.925 -123.925 -21.595 -123.595 ;
        RECT -21.925 -125.285 -21.595 -124.955 ;
        RECT -21.925 -128.005 -21.595 -127.675 ;
        RECT -21.925 -134.805 -21.595 -134.475 ;
        RECT -21.925 -138.885 -21.595 -138.555 ;
        RECT -21.925 -141.605 -21.595 -141.275 ;
        RECT -21.925 -142.965 -21.595 -142.635 ;
        RECT -21.925 -145.685 -21.595 -145.355 ;
        RECT -21.925 -147.045 -21.595 -146.715 ;
        RECT -21.925 -151.125 -21.595 -150.795 ;
        RECT -21.925 -152.485 -21.595 -152.155 ;
        RECT -21.925 -156.565 -21.595 -156.235 ;
        RECT -21.925 -157.925 -21.595 -157.595 ;
        RECT -21.925 -159.285 -21.595 -158.955 ;
        RECT -21.925 -160.645 -21.595 -160.315 ;
        RECT -21.925 -162.005 -21.595 -161.675 ;
        RECT -21.925 -163.365 -21.595 -163.035 ;
        RECT -21.925 -164.725 -21.595 -164.395 ;
        RECT -21.925 -166.085 -21.595 -165.755 ;
        RECT -21.925 -167.445 -21.595 -167.115 ;
        RECT -21.925 -170.165 -21.595 -169.835 ;
        RECT -21.925 -174.245 -21.595 -173.915 ;
        RECT -21.925 -175.725 -21.595 -175.395 ;
        RECT -21.925 -176.965 -21.595 -176.635 ;
        RECT -21.925 -178.325 -21.595 -177.995 ;
        RECT -21.925 -180.57 -21.595 -179.44 ;
        RECT -21.92 -180.685 -21.6 -63.755 ;
    END
    PORT
      LAYER met3 ;
        RECT -20.565 241.32 -20.235 242.45 ;
        RECT -20.565 239.195 -20.235 239.525 ;
        RECT -20.565 237.835 -20.235 238.165 ;
        RECT -20.565 236.475 -20.235 236.805 ;
        RECT -20.565 235.115 -20.235 235.445 ;
        RECT -20.565 233.755 -20.235 234.085 ;
        RECT -20.565 232.395 -20.235 232.725 ;
        RECT -20.565 231.035 -20.235 231.365 ;
        RECT -20.565 229.675 -20.235 230.005 ;
        RECT -20.565 228.315 -20.235 228.645 ;
        RECT -20.565 226.955 -20.235 227.285 ;
        RECT -20.565 225.595 -20.235 225.925 ;
        RECT -20.565 224.235 -20.235 224.565 ;
        RECT -20.565 222.875 -20.235 223.205 ;
        RECT -20.565 221.515 -20.235 221.845 ;
        RECT -20.565 220.155 -20.235 220.485 ;
        RECT -20.565 218.795 -20.235 219.125 ;
        RECT -20.565 217.435 -20.235 217.765 ;
        RECT -20.565 216.075 -20.235 216.405 ;
        RECT -20.565 214.715 -20.235 215.045 ;
        RECT -20.565 213.355 -20.235 213.685 ;
        RECT -20.565 211.995 -20.235 212.325 ;
        RECT -20.565 210.635 -20.235 210.965 ;
        RECT -20.565 209.275 -20.235 209.605 ;
        RECT -20.565 207.915 -20.235 208.245 ;
        RECT -20.565 206.555 -20.235 206.885 ;
        RECT -20.565 205.195 -20.235 205.525 ;
        RECT -20.565 203.835 -20.235 204.165 ;
        RECT -20.565 202.475 -20.235 202.805 ;
        RECT -20.565 201.115 -20.235 201.445 ;
        RECT -20.565 199.755 -20.235 200.085 ;
        RECT -20.565 198.395 -20.235 198.725 ;
        RECT -20.565 197.035 -20.235 197.365 ;
        RECT -20.565 195.675 -20.235 196.005 ;
        RECT -20.565 194.315 -20.235 194.645 ;
        RECT -20.565 192.955 -20.235 193.285 ;
        RECT -20.565 191.595 -20.235 191.925 ;
        RECT -20.565 190.235 -20.235 190.565 ;
        RECT -20.565 188.875 -20.235 189.205 ;
        RECT -20.565 187.515 -20.235 187.845 ;
        RECT -20.565 186.155 -20.235 186.485 ;
        RECT -20.565 184.795 -20.235 185.125 ;
        RECT -20.565 183.435 -20.235 183.765 ;
        RECT -20.565 182.075 -20.235 182.405 ;
        RECT -20.565 180.715 -20.235 181.045 ;
        RECT -20.565 179.355 -20.235 179.685 ;
        RECT -20.565 177.995 -20.235 178.325 ;
        RECT -20.565 176.635 -20.235 176.965 ;
        RECT -20.565 175.275 -20.235 175.605 ;
        RECT -20.565 173.915 -20.235 174.245 ;
        RECT -20.565 172.555 -20.235 172.885 ;
        RECT -20.565 171.195 -20.235 171.525 ;
        RECT -20.565 169.835 -20.235 170.165 ;
        RECT -20.565 168.475 -20.235 168.805 ;
        RECT -20.565 167.115 -20.235 167.445 ;
        RECT -20.565 165.755 -20.235 166.085 ;
        RECT -20.565 164.395 -20.235 164.725 ;
        RECT -20.565 163.035 -20.235 163.365 ;
        RECT -20.565 161.675 -20.235 162.005 ;
        RECT -20.565 160.315 -20.235 160.645 ;
        RECT -20.565 158.955 -20.235 159.285 ;
        RECT -20.565 157.595 -20.235 157.925 ;
        RECT -20.565 156.235 -20.235 156.565 ;
        RECT -20.565 154.875 -20.235 155.205 ;
        RECT -20.565 153.515 -20.235 153.845 ;
        RECT -20.565 152.155 -20.235 152.485 ;
        RECT -20.565 150.795 -20.235 151.125 ;
        RECT -20.565 149.435 -20.235 149.765 ;
        RECT -20.565 148.075 -20.235 148.405 ;
        RECT -20.565 146.715 -20.235 147.045 ;
        RECT -20.565 145.355 -20.235 145.685 ;
        RECT -20.565 143.995 -20.235 144.325 ;
        RECT -20.565 142.635 -20.235 142.965 ;
        RECT -20.565 141.275 -20.235 141.605 ;
        RECT -20.565 139.915 -20.235 140.245 ;
        RECT -20.565 138.555 -20.235 138.885 ;
        RECT -20.565 137.195 -20.235 137.525 ;
        RECT -20.565 135.835 -20.235 136.165 ;
        RECT -20.565 134.475 -20.235 134.805 ;
        RECT -20.565 133.115 -20.235 133.445 ;
        RECT -20.565 131.755 -20.235 132.085 ;
        RECT -20.565 130.395 -20.235 130.725 ;
        RECT -20.565 129.035 -20.235 129.365 ;
        RECT -20.565 127.675 -20.235 128.005 ;
        RECT -20.565 126.315 -20.235 126.645 ;
        RECT -20.565 124.955 -20.235 125.285 ;
        RECT -20.565 123.595 -20.235 123.925 ;
        RECT -20.565 122.235 -20.235 122.565 ;
        RECT -20.565 120.875 -20.235 121.205 ;
        RECT -20.565 119.515 -20.235 119.845 ;
        RECT -20.565 118.155 -20.235 118.485 ;
        RECT -20.565 116.795 -20.235 117.125 ;
        RECT -20.565 115.435 -20.235 115.765 ;
        RECT -20.565 114.075 -20.235 114.405 ;
        RECT -20.565 112.715 -20.235 113.045 ;
        RECT -20.565 111.355 -20.235 111.685 ;
        RECT -20.565 109.995 -20.235 110.325 ;
        RECT -20.565 108.635 -20.235 108.965 ;
        RECT -20.565 107.275 -20.235 107.605 ;
        RECT -20.565 105.915 -20.235 106.245 ;
        RECT -20.565 104.555 -20.235 104.885 ;
        RECT -20.565 103.195 -20.235 103.525 ;
        RECT -20.565 101.835 -20.235 102.165 ;
        RECT -20.565 100.475 -20.235 100.805 ;
        RECT -20.565 99.115 -20.235 99.445 ;
        RECT -20.565 97.755 -20.235 98.085 ;
        RECT -20.565 96.395 -20.235 96.725 ;
        RECT -20.565 95.035 -20.235 95.365 ;
        RECT -20.565 93.675 -20.235 94.005 ;
        RECT -20.565 92.315 -20.235 92.645 ;
        RECT -20.565 90.955 -20.235 91.285 ;
        RECT -20.565 89.595 -20.235 89.925 ;
        RECT -20.565 88.235 -20.235 88.565 ;
        RECT -20.565 86.875 -20.235 87.205 ;
        RECT -20.565 85.515 -20.235 85.845 ;
        RECT -20.565 84.155 -20.235 84.485 ;
        RECT -20.565 82.795 -20.235 83.125 ;
        RECT -20.565 81.435 -20.235 81.765 ;
        RECT -20.565 80.075 -20.235 80.405 ;
        RECT -20.565 78.715 -20.235 79.045 ;
        RECT -20.565 77.355 -20.235 77.685 ;
        RECT -20.565 75.995 -20.235 76.325 ;
        RECT -20.565 74.635 -20.235 74.965 ;
        RECT -20.565 73.275 -20.235 73.605 ;
        RECT -20.565 71.915 -20.235 72.245 ;
        RECT -20.565 70.555 -20.235 70.885 ;
        RECT -20.565 69.195 -20.235 69.525 ;
        RECT -20.565 67.835 -20.235 68.165 ;
        RECT -20.565 66.475 -20.235 66.805 ;
        RECT -20.565 65.115 -20.235 65.445 ;
        RECT -20.565 63.755 -20.235 64.085 ;
        RECT -20.565 62.395 -20.235 62.725 ;
        RECT -20.565 61.035 -20.235 61.365 ;
        RECT -20.565 59.675 -20.235 60.005 ;
        RECT -20.565 58.315 -20.235 58.645 ;
        RECT -20.565 56.955 -20.235 57.285 ;
        RECT -20.565 55.595 -20.235 55.925 ;
        RECT -20.565 54.235 -20.235 54.565 ;
        RECT -20.565 52.875 -20.235 53.205 ;
        RECT -20.565 51.515 -20.235 51.845 ;
        RECT -20.565 50.155 -20.235 50.485 ;
        RECT -20.565 48.795 -20.235 49.125 ;
        RECT -20.565 47.435 -20.235 47.765 ;
        RECT -20.565 46.075 -20.235 46.405 ;
        RECT -20.565 44.715 -20.235 45.045 ;
        RECT -20.565 43.355 -20.235 43.685 ;
        RECT -20.565 41.995 -20.235 42.325 ;
        RECT -20.565 40.635 -20.235 40.965 ;
        RECT -20.565 39.275 -20.235 39.605 ;
        RECT -20.565 37.915 -20.235 38.245 ;
        RECT -20.565 36.555 -20.235 36.885 ;
        RECT -20.565 35.195 -20.235 35.525 ;
        RECT -20.565 33.835 -20.235 34.165 ;
        RECT -20.565 32.475 -20.235 32.805 ;
        RECT -20.565 31.115 -20.235 31.445 ;
        RECT -20.565 29.755 -20.235 30.085 ;
        RECT -20.565 28.395 -20.235 28.725 ;
        RECT -20.565 27.035 -20.235 27.365 ;
        RECT -20.565 25.675 -20.235 26.005 ;
        RECT -20.565 24.315 -20.235 24.645 ;
        RECT -20.565 22.955 -20.235 23.285 ;
        RECT -20.565 21.595 -20.235 21.925 ;
        RECT -20.565 20.235 -20.235 20.565 ;
        RECT -20.565 18.875 -20.235 19.205 ;
        RECT -20.565 17.515 -20.235 17.845 ;
        RECT -20.565 16.155 -20.235 16.485 ;
        RECT -20.565 14.795 -20.235 15.125 ;
        RECT -20.565 13.435 -20.235 13.765 ;
        RECT -20.565 12.075 -20.235 12.405 ;
        RECT -20.565 10.715 -20.235 11.045 ;
        RECT -20.565 9.355 -20.235 9.685 ;
        RECT -20.565 7.995 -20.235 8.325 ;
        RECT -20.565 6.635 -20.235 6.965 ;
        RECT -20.565 5.275 -20.235 5.605 ;
        RECT -20.565 3.915 -20.235 4.245 ;
        RECT -20.565 2.555 -20.235 2.885 ;
        RECT -20.565 1.195 -20.235 1.525 ;
        RECT -20.565 -0.165 -20.235 0.165 ;
        RECT -20.565 -2.885 -20.235 -2.555 ;
        RECT -20.565 -4.245 -20.235 -3.915 ;
        RECT -20.565 -8.325 -20.235 -7.995 ;
        RECT -20.565 -9.685 -20.235 -9.355 ;
        RECT -20.565 -14.95 -20.235 -14.62 ;
        RECT -20.565 -17.845 -20.235 -17.515 ;
        RECT -20.565 -19.79 -20.235 -19.46 ;
        RECT -20.565 -20.565 -20.235 -20.235 ;
        RECT -20.56 -22.6 -20.24 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -20.565 -28.725 -20.235 -28.395 ;
        RECT -20.565 -30.085 -20.235 -29.755 ;
        RECT -20.565 -31.445 -20.235 -31.115 ;
        RECT -20.565 -32.805 -20.235 -32.475 ;
        RECT -20.565 -35.525 -20.235 -35.195 ;
        RECT -20.565 -36.885 -20.235 -36.555 ;
        RECT -20.565 -37.93 -20.235 -37.6 ;
        RECT -20.565 -40.965 -20.235 -40.635 ;
        RECT -20.565 -42.77 -20.235 -42.44 ;
        RECT -20.565 -43.685 -20.235 -43.355 ;
        RECT -20.565 -50.485 -20.235 -50.155 ;
        RECT -20.565 -51.845 -20.235 -51.515 ;
        RECT -20.565 -53.205 -20.235 -52.875 ;
        RECT -20.565 -54.565 -20.235 -54.235 ;
        RECT -20.565 -55.925 -20.235 -55.595 ;
        RECT -20.565 -57.285 -20.235 -56.955 ;
        RECT -20.565 -58.645 -20.235 -58.315 ;
        RECT -20.565 -60.005 -20.235 -59.675 ;
        RECT -20.565 -61.365 -20.235 -61.035 ;
        RECT -20.565 -62.725 -20.235 -62.395 ;
        RECT -20.565 -64.085 -20.235 -63.755 ;
        RECT -20.565 -65.445 -20.235 -65.115 ;
        RECT -20.565 -66.805 -20.235 -66.475 ;
        RECT -20.565 -68.165 -20.235 -67.835 ;
        RECT -20.565 -69.525 -20.235 -69.195 ;
        RECT -20.565 -70.885 -20.235 -70.555 ;
        RECT -20.565 -72.245 -20.235 -71.915 ;
        RECT -20.565 -74.965 -20.235 -74.635 ;
        RECT -20.565 -77.685 -20.235 -77.355 ;
        RECT -20.565 -79.045 -20.235 -78.715 ;
        RECT -20.565 -81.765 -20.235 -81.435 ;
        RECT -20.565 -83.125 -20.235 -82.795 ;
        RECT -20.565 -84.485 -20.235 -84.155 ;
        RECT -20.565 -87.205 -20.235 -86.875 ;
        RECT -20.565 -89.925 -20.235 -89.595 ;
        RECT -20.565 -91.285 -20.235 -90.955 ;
        RECT -20.565 -92.645 -20.235 -92.315 ;
        RECT -20.565 -94.005 -20.235 -93.675 ;
        RECT -20.565 -96.725 -20.235 -96.395 ;
        RECT -20.565 -98.085 -20.235 -97.755 ;
        RECT -20.565 -100.805 -20.235 -100.475 ;
        RECT -20.565 -102.165 -20.235 -101.835 ;
        RECT -20.565 -104.885 -20.235 -104.555 ;
        RECT -20.565 -106.245 -20.235 -105.915 ;
        RECT -20.565 -108.965 -20.235 -108.635 ;
        RECT -20.565 -113.045 -20.235 -112.715 ;
        RECT -20.565 -114.405 -20.235 -114.075 ;
        RECT -20.565 -115.765 -20.235 -115.435 ;
        RECT -20.565 -117.125 -20.235 -116.795 ;
        RECT -20.565 -118.485 -20.235 -118.155 ;
        RECT -20.565 -123.925 -20.235 -123.595 ;
        RECT -20.565 -125.285 -20.235 -124.955 ;
        RECT -20.565 -128.005 -20.235 -127.675 ;
        RECT -20.565 -134.805 -20.235 -134.475 ;
        RECT -20.565 -138.885 -20.235 -138.555 ;
        RECT -20.565 -142.965 -20.235 -142.635 ;
        RECT -20.565 -145.685 -20.235 -145.355 ;
        RECT -20.565 -147.045 -20.235 -146.715 ;
        RECT -20.565 -151.125 -20.235 -150.795 ;
        RECT -20.565 -152.485 -20.235 -152.155 ;
        RECT -20.565 -156.565 -20.235 -156.235 ;
        RECT -20.565 -157.925 -20.235 -157.595 ;
        RECT -20.565 -159.285 -20.235 -158.955 ;
        RECT -20.565 -160.645 -20.235 -160.315 ;
        RECT -20.565 -162.005 -20.235 -161.675 ;
        RECT -20.565 -163.365 -20.235 -163.035 ;
        RECT -20.565 -164.725 -20.235 -164.395 ;
        RECT -20.565 -166.085 -20.235 -165.755 ;
        RECT -20.565 -167.445 -20.235 -167.115 ;
        RECT -20.565 -170.165 -20.235 -169.835 ;
        RECT -20.565 -172.885 -20.235 -172.555 ;
        RECT -20.565 -174.245 -20.235 -173.915 ;
        RECT -20.565 -175.725 -20.235 -175.395 ;
        RECT -20.565 -176.965 -20.235 -176.635 ;
        RECT -20.565 -178.325 -20.235 -177.995 ;
        RECT -20.565 -180.57 -20.235 -179.44 ;
        RECT -20.56 -180.685 -20.24 -28.395 ;
    END
    PORT
      LAYER met3 ;
        RECT -19.205 241.32 -18.875 242.45 ;
        RECT -19.205 239.195 -18.875 239.525 ;
        RECT -19.205 237.835 -18.875 238.165 ;
        RECT -19.205 236.475 -18.875 236.805 ;
        RECT -19.205 235.115 -18.875 235.445 ;
        RECT -19.205 233.755 -18.875 234.085 ;
        RECT -19.205 232.395 -18.875 232.725 ;
        RECT -19.205 231.035 -18.875 231.365 ;
        RECT -19.205 229.675 -18.875 230.005 ;
        RECT -19.205 228.315 -18.875 228.645 ;
        RECT -19.205 226.955 -18.875 227.285 ;
        RECT -19.205 225.595 -18.875 225.925 ;
        RECT -19.205 224.235 -18.875 224.565 ;
        RECT -19.205 222.875 -18.875 223.205 ;
        RECT -19.205 221.515 -18.875 221.845 ;
        RECT -19.205 220.155 -18.875 220.485 ;
        RECT -19.205 218.795 -18.875 219.125 ;
        RECT -19.205 217.435 -18.875 217.765 ;
        RECT -19.205 216.075 -18.875 216.405 ;
        RECT -19.205 214.715 -18.875 215.045 ;
        RECT -19.205 213.355 -18.875 213.685 ;
        RECT -19.205 211.995 -18.875 212.325 ;
        RECT -19.205 210.635 -18.875 210.965 ;
        RECT -19.205 209.275 -18.875 209.605 ;
        RECT -19.205 207.915 -18.875 208.245 ;
        RECT -19.205 206.555 -18.875 206.885 ;
        RECT -19.205 205.195 -18.875 205.525 ;
        RECT -19.205 203.835 -18.875 204.165 ;
        RECT -19.205 202.475 -18.875 202.805 ;
        RECT -19.205 201.115 -18.875 201.445 ;
        RECT -19.205 199.755 -18.875 200.085 ;
        RECT -19.205 198.395 -18.875 198.725 ;
        RECT -19.205 197.035 -18.875 197.365 ;
        RECT -19.205 195.675 -18.875 196.005 ;
        RECT -19.205 194.315 -18.875 194.645 ;
        RECT -19.205 192.955 -18.875 193.285 ;
        RECT -19.205 191.595 -18.875 191.925 ;
        RECT -19.205 190.235 -18.875 190.565 ;
        RECT -19.205 188.875 -18.875 189.205 ;
        RECT -19.205 187.515 -18.875 187.845 ;
        RECT -19.205 186.155 -18.875 186.485 ;
        RECT -19.205 184.795 -18.875 185.125 ;
        RECT -19.205 183.435 -18.875 183.765 ;
        RECT -19.205 182.075 -18.875 182.405 ;
        RECT -19.205 180.715 -18.875 181.045 ;
        RECT -19.205 179.355 -18.875 179.685 ;
        RECT -19.205 177.995 -18.875 178.325 ;
        RECT -19.205 176.635 -18.875 176.965 ;
        RECT -19.205 175.275 -18.875 175.605 ;
        RECT -19.205 173.915 -18.875 174.245 ;
        RECT -19.205 172.555 -18.875 172.885 ;
        RECT -19.205 171.195 -18.875 171.525 ;
        RECT -19.205 169.835 -18.875 170.165 ;
        RECT -19.205 168.475 -18.875 168.805 ;
        RECT -19.205 167.115 -18.875 167.445 ;
        RECT -19.205 165.755 -18.875 166.085 ;
        RECT -19.205 164.395 -18.875 164.725 ;
        RECT -19.205 163.035 -18.875 163.365 ;
        RECT -19.205 161.675 -18.875 162.005 ;
        RECT -19.205 160.315 -18.875 160.645 ;
        RECT -19.205 158.955 -18.875 159.285 ;
        RECT -19.205 157.595 -18.875 157.925 ;
        RECT -19.205 156.235 -18.875 156.565 ;
        RECT -19.205 154.875 -18.875 155.205 ;
        RECT -19.205 153.515 -18.875 153.845 ;
        RECT -19.205 152.155 -18.875 152.485 ;
        RECT -19.205 150.795 -18.875 151.125 ;
        RECT -19.205 149.435 -18.875 149.765 ;
        RECT -19.205 148.075 -18.875 148.405 ;
        RECT -19.205 146.715 -18.875 147.045 ;
        RECT -19.205 145.355 -18.875 145.685 ;
        RECT -19.205 143.995 -18.875 144.325 ;
        RECT -19.205 142.635 -18.875 142.965 ;
        RECT -19.205 141.275 -18.875 141.605 ;
        RECT -19.205 139.915 -18.875 140.245 ;
        RECT -19.205 138.555 -18.875 138.885 ;
        RECT -19.205 137.195 -18.875 137.525 ;
        RECT -19.205 135.835 -18.875 136.165 ;
        RECT -19.205 134.475 -18.875 134.805 ;
        RECT -19.205 133.115 -18.875 133.445 ;
        RECT -19.205 131.755 -18.875 132.085 ;
        RECT -19.205 130.395 -18.875 130.725 ;
        RECT -19.205 129.035 -18.875 129.365 ;
        RECT -19.205 127.675 -18.875 128.005 ;
        RECT -19.205 126.315 -18.875 126.645 ;
        RECT -19.205 124.955 -18.875 125.285 ;
        RECT -19.205 123.595 -18.875 123.925 ;
        RECT -19.205 122.235 -18.875 122.565 ;
        RECT -19.205 120.875 -18.875 121.205 ;
        RECT -19.205 119.515 -18.875 119.845 ;
        RECT -19.205 118.155 -18.875 118.485 ;
        RECT -19.205 116.795 -18.875 117.125 ;
        RECT -19.205 115.435 -18.875 115.765 ;
        RECT -19.205 114.075 -18.875 114.405 ;
        RECT -19.205 112.715 -18.875 113.045 ;
        RECT -19.205 111.355 -18.875 111.685 ;
        RECT -19.205 109.995 -18.875 110.325 ;
        RECT -19.205 108.635 -18.875 108.965 ;
        RECT -19.205 107.275 -18.875 107.605 ;
        RECT -19.205 105.915 -18.875 106.245 ;
        RECT -19.205 104.555 -18.875 104.885 ;
        RECT -19.205 103.195 -18.875 103.525 ;
        RECT -19.205 101.835 -18.875 102.165 ;
        RECT -19.205 100.475 -18.875 100.805 ;
        RECT -19.205 99.115 -18.875 99.445 ;
        RECT -19.205 97.755 -18.875 98.085 ;
        RECT -19.205 96.395 -18.875 96.725 ;
        RECT -19.205 95.035 -18.875 95.365 ;
        RECT -19.205 93.675 -18.875 94.005 ;
        RECT -19.205 92.315 -18.875 92.645 ;
        RECT -19.205 90.955 -18.875 91.285 ;
        RECT -19.205 89.595 -18.875 89.925 ;
        RECT -19.205 88.235 -18.875 88.565 ;
        RECT -19.205 86.875 -18.875 87.205 ;
        RECT -19.205 85.515 -18.875 85.845 ;
        RECT -19.205 84.155 -18.875 84.485 ;
        RECT -19.205 82.795 -18.875 83.125 ;
        RECT -19.205 81.435 -18.875 81.765 ;
        RECT -19.205 80.075 -18.875 80.405 ;
        RECT -19.205 78.715 -18.875 79.045 ;
        RECT -19.205 77.355 -18.875 77.685 ;
        RECT -19.205 75.995 -18.875 76.325 ;
        RECT -19.205 74.635 -18.875 74.965 ;
        RECT -19.205 73.275 -18.875 73.605 ;
        RECT -19.205 71.915 -18.875 72.245 ;
        RECT -19.205 70.555 -18.875 70.885 ;
        RECT -19.205 69.195 -18.875 69.525 ;
        RECT -19.205 67.835 -18.875 68.165 ;
        RECT -19.205 66.475 -18.875 66.805 ;
        RECT -19.205 65.115 -18.875 65.445 ;
        RECT -19.205 63.755 -18.875 64.085 ;
        RECT -19.205 62.395 -18.875 62.725 ;
        RECT -19.205 61.035 -18.875 61.365 ;
        RECT -19.205 59.675 -18.875 60.005 ;
        RECT -19.205 58.315 -18.875 58.645 ;
        RECT -19.205 56.955 -18.875 57.285 ;
        RECT -19.205 55.595 -18.875 55.925 ;
        RECT -19.205 54.235 -18.875 54.565 ;
        RECT -19.205 52.875 -18.875 53.205 ;
        RECT -19.205 51.515 -18.875 51.845 ;
        RECT -19.205 50.155 -18.875 50.485 ;
        RECT -19.205 48.795 -18.875 49.125 ;
        RECT -19.205 47.435 -18.875 47.765 ;
        RECT -19.205 46.075 -18.875 46.405 ;
        RECT -19.205 44.715 -18.875 45.045 ;
        RECT -19.205 43.355 -18.875 43.685 ;
        RECT -19.205 41.995 -18.875 42.325 ;
        RECT -19.205 40.635 -18.875 40.965 ;
        RECT -19.205 39.275 -18.875 39.605 ;
        RECT -19.205 37.915 -18.875 38.245 ;
        RECT -19.205 36.555 -18.875 36.885 ;
        RECT -19.205 35.195 -18.875 35.525 ;
        RECT -19.205 33.835 -18.875 34.165 ;
        RECT -19.205 32.475 -18.875 32.805 ;
        RECT -19.205 31.115 -18.875 31.445 ;
        RECT -19.205 29.755 -18.875 30.085 ;
        RECT -19.205 28.395 -18.875 28.725 ;
        RECT -19.205 27.035 -18.875 27.365 ;
        RECT -19.205 25.675 -18.875 26.005 ;
        RECT -19.205 24.315 -18.875 24.645 ;
        RECT -19.205 22.955 -18.875 23.285 ;
        RECT -19.205 21.595 -18.875 21.925 ;
        RECT -19.205 20.235 -18.875 20.565 ;
        RECT -19.205 18.875 -18.875 19.205 ;
        RECT -19.205 17.515 -18.875 17.845 ;
        RECT -19.205 16.155 -18.875 16.485 ;
        RECT -19.205 14.795 -18.875 15.125 ;
        RECT -19.205 13.435 -18.875 13.765 ;
        RECT -19.205 12.075 -18.875 12.405 ;
        RECT -19.205 10.715 -18.875 11.045 ;
        RECT -19.205 9.355 -18.875 9.685 ;
        RECT -19.205 7.995 -18.875 8.325 ;
        RECT -19.205 6.635 -18.875 6.965 ;
        RECT -19.205 5.275 -18.875 5.605 ;
        RECT -19.205 3.915 -18.875 4.245 ;
        RECT -19.205 2.555 -18.875 2.885 ;
        RECT -19.205 1.195 -18.875 1.525 ;
        RECT -19.205 -0.165 -18.875 0.165 ;
        RECT -19.205 -2.885 -18.875 -2.555 ;
        RECT -19.205 -4.245 -18.875 -3.915 ;
        RECT -19.205 -8.325 -18.875 -7.995 ;
        RECT -19.205 -9.685 -18.875 -9.355 ;
        RECT -19.205 -14.95 -18.875 -14.62 ;
        RECT -19.205 -17.845 -18.875 -17.515 ;
        RECT -19.205 -19.79 -18.875 -19.46 ;
        RECT -19.205 -20.565 -18.875 -20.235 ;
        RECT -19.2 -21.92 -18.88 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -28.725 -68.165 -28.395 -67.835 ;
        RECT -28.725 -69.525 -28.395 -69.195 ;
        RECT -28.725 -70.885 -28.395 -70.555 ;
        RECT -28.725 -72.245 -28.395 -71.915 ;
        RECT -28.725 -73.605 -28.395 -73.275 ;
        RECT -28.725 -74.965 -28.395 -74.635 ;
        RECT -28.725 -76.325 -28.395 -75.995 ;
        RECT -28.725 -77.685 -28.395 -77.355 ;
        RECT -28.725 -79.045 -28.395 -78.715 ;
        RECT -28.725 -80.405 -28.395 -80.075 ;
        RECT -28.725 -81.765 -28.395 -81.435 ;
        RECT -28.725 -83.125 -28.395 -82.795 ;
        RECT -28.725 -84.485 -28.395 -84.155 ;
        RECT -28.725 -85.845 -28.395 -85.515 ;
        RECT -28.725 -87.205 -28.395 -86.875 ;
        RECT -28.725 -88.565 -28.395 -88.235 ;
        RECT -28.725 -89.925 -28.395 -89.595 ;
        RECT -28.725 -92.645 -28.395 -92.315 ;
        RECT -28.725 -94.005 -28.395 -93.675 ;
        RECT -28.725 -95.365 -28.395 -95.035 ;
        RECT -28.725 -96.725 -28.395 -96.395 ;
        RECT -28.725 -98.73 -28.395 -98.4 ;
        RECT -28.725 -99.445 -28.395 -99.115 ;
        RECT -28.725 -102.165 -28.395 -101.835 ;
        RECT -28.725 -103.525 -28.395 -103.195 ;
        RECT -28.725 -104.885 -28.395 -104.555 ;
        RECT -28.725 -106.87 -28.395 -106.54 ;
        RECT -28.725 -107.605 -28.395 -107.275 ;
        RECT -28.725 -108.965 -28.395 -108.635 ;
        RECT -28.725 -113.045 -28.395 -112.715 ;
        RECT -28.725 -114.405 -28.395 -114.075 ;
        RECT -28.725 -115.765 -28.395 -115.435 ;
        RECT -28.725 -117.125 -28.395 -116.795 ;
        RECT -28.725 -118.485 -28.395 -118.155 ;
        RECT -28.725 -122.565 -28.395 -122.235 ;
        RECT -28.725 -125.285 -28.395 -124.955 ;
        RECT -28.725 -126.645 -28.395 -126.315 ;
        RECT -28.725 -128.005 -28.395 -127.675 ;
        RECT -28.725 -129.365 -28.395 -129.035 ;
        RECT -28.725 -133.445 -28.395 -133.115 ;
        RECT -28.725 -134.805 -28.395 -134.475 ;
        RECT -28.725 -136.165 -28.395 -135.835 ;
        RECT -28.725 -138.885 -28.395 -138.555 ;
        RECT -28.725 -141.605 -28.395 -141.275 ;
        RECT -28.725 -142.965 -28.395 -142.635 ;
        RECT -28.725 -144.325 -28.395 -143.995 ;
        RECT -28.725 -145.685 -28.395 -145.355 ;
        RECT -28.725 -147.045 -28.395 -146.715 ;
        RECT -28.725 -148.405 -28.395 -148.075 ;
        RECT -28.725 -151.125 -28.395 -150.795 ;
        RECT -28.725 -152.485 -28.395 -152.155 ;
        RECT -28.725 -156.565 -28.395 -156.235 ;
        RECT -28.725 -157.925 -28.395 -157.595 ;
        RECT -28.725 -159.285 -28.395 -158.955 ;
        RECT -28.725 -160.645 -28.395 -160.315 ;
        RECT -28.725 -162.005 -28.395 -161.675 ;
        RECT -28.725 -163.365 -28.395 -163.035 ;
        RECT -28.725 -164.725 -28.395 -164.395 ;
        RECT -28.725 -166.085 -28.395 -165.755 ;
        RECT -28.725 -167.445 -28.395 -167.115 ;
        RECT -28.725 -170.165 -28.395 -169.835 ;
        RECT -28.725 -174.245 -28.395 -173.915 ;
        RECT -28.725 -176.965 -28.395 -176.635 ;
        RECT -28.725 -178.325 -28.395 -177.995 ;
        RECT -28.725 -180.57 -28.395 -179.44 ;
        RECT -28.72 -180.685 -28.4 -67.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -27.365 241.32 -27.035 242.45 ;
        RECT -27.365 239.195 -27.035 239.525 ;
        RECT -27.365 237.835 -27.035 238.165 ;
        RECT -27.365 236.475 -27.035 236.805 ;
        RECT -27.365 235.115 -27.035 235.445 ;
        RECT -27.365 233.755 -27.035 234.085 ;
        RECT -27.365 232.395 -27.035 232.725 ;
        RECT -27.365 231.035 -27.035 231.365 ;
        RECT -27.365 229.675 -27.035 230.005 ;
        RECT -27.365 228.315 -27.035 228.645 ;
        RECT -27.365 226.955 -27.035 227.285 ;
        RECT -27.365 225.595 -27.035 225.925 ;
        RECT -27.365 224.235 -27.035 224.565 ;
        RECT -27.365 222.875 -27.035 223.205 ;
        RECT -27.365 221.515 -27.035 221.845 ;
        RECT -27.365 220.155 -27.035 220.485 ;
        RECT -27.365 218.795 -27.035 219.125 ;
        RECT -27.365 217.435 -27.035 217.765 ;
        RECT -27.365 216.075 -27.035 216.405 ;
        RECT -27.365 214.715 -27.035 215.045 ;
        RECT -27.365 213.355 -27.035 213.685 ;
        RECT -27.365 211.995 -27.035 212.325 ;
        RECT -27.365 210.635 -27.035 210.965 ;
        RECT -27.365 209.275 -27.035 209.605 ;
        RECT -27.365 207.915 -27.035 208.245 ;
        RECT -27.365 206.555 -27.035 206.885 ;
        RECT -27.365 205.195 -27.035 205.525 ;
        RECT -27.365 203.835 -27.035 204.165 ;
        RECT -27.365 202.475 -27.035 202.805 ;
        RECT -27.365 201.115 -27.035 201.445 ;
        RECT -27.365 199.755 -27.035 200.085 ;
        RECT -27.365 198.395 -27.035 198.725 ;
        RECT -27.365 197.035 -27.035 197.365 ;
        RECT -27.365 195.675 -27.035 196.005 ;
        RECT -27.365 194.315 -27.035 194.645 ;
        RECT -27.365 192.955 -27.035 193.285 ;
        RECT -27.365 191.595 -27.035 191.925 ;
        RECT -27.365 190.235 -27.035 190.565 ;
        RECT -27.365 188.875 -27.035 189.205 ;
        RECT -27.365 187.515 -27.035 187.845 ;
        RECT -27.365 186.155 -27.035 186.485 ;
        RECT -27.365 184.795 -27.035 185.125 ;
        RECT -27.365 183.435 -27.035 183.765 ;
        RECT -27.365 182.075 -27.035 182.405 ;
        RECT -27.365 180.715 -27.035 181.045 ;
        RECT -27.365 179.355 -27.035 179.685 ;
        RECT -27.365 177.995 -27.035 178.325 ;
        RECT -27.365 176.635 -27.035 176.965 ;
        RECT -27.365 175.275 -27.035 175.605 ;
        RECT -27.365 173.915 -27.035 174.245 ;
        RECT -27.365 172.555 -27.035 172.885 ;
        RECT -27.365 171.195 -27.035 171.525 ;
        RECT -27.365 169.835 -27.035 170.165 ;
        RECT -27.365 168.475 -27.035 168.805 ;
        RECT -27.365 167.115 -27.035 167.445 ;
        RECT -27.365 165.755 -27.035 166.085 ;
        RECT -27.365 164.395 -27.035 164.725 ;
        RECT -27.365 163.035 -27.035 163.365 ;
        RECT -27.365 161.675 -27.035 162.005 ;
        RECT -27.365 160.315 -27.035 160.645 ;
        RECT -27.365 158.955 -27.035 159.285 ;
        RECT -27.365 157.595 -27.035 157.925 ;
        RECT -27.365 156.235 -27.035 156.565 ;
        RECT -27.365 154.875 -27.035 155.205 ;
        RECT -27.365 153.515 -27.035 153.845 ;
        RECT -27.365 152.155 -27.035 152.485 ;
        RECT -27.365 150.795 -27.035 151.125 ;
        RECT -27.365 149.435 -27.035 149.765 ;
        RECT -27.365 148.075 -27.035 148.405 ;
        RECT -27.365 146.715 -27.035 147.045 ;
        RECT -27.365 145.355 -27.035 145.685 ;
        RECT -27.365 143.995 -27.035 144.325 ;
        RECT -27.365 142.635 -27.035 142.965 ;
        RECT -27.365 141.275 -27.035 141.605 ;
        RECT -27.365 139.915 -27.035 140.245 ;
        RECT -27.365 138.555 -27.035 138.885 ;
        RECT -27.365 137.195 -27.035 137.525 ;
        RECT -27.365 135.835 -27.035 136.165 ;
        RECT -27.365 134.475 -27.035 134.805 ;
        RECT -27.365 133.115 -27.035 133.445 ;
        RECT -27.365 131.755 -27.035 132.085 ;
        RECT -27.365 130.395 -27.035 130.725 ;
        RECT -27.365 129.035 -27.035 129.365 ;
        RECT -27.365 127.675 -27.035 128.005 ;
        RECT -27.365 126.315 -27.035 126.645 ;
        RECT -27.365 124.955 -27.035 125.285 ;
        RECT -27.365 123.595 -27.035 123.925 ;
        RECT -27.365 122.235 -27.035 122.565 ;
        RECT -27.365 120.875 -27.035 121.205 ;
        RECT -27.365 119.515 -27.035 119.845 ;
        RECT -27.365 118.155 -27.035 118.485 ;
        RECT -27.365 116.795 -27.035 117.125 ;
        RECT -27.365 115.435 -27.035 115.765 ;
        RECT -27.365 114.075 -27.035 114.405 ;
        RECT -27.365 112.715 -27.035 113.045 ;
        RECT -27.365 111.355 -27.035 111.685 ;
        RECT -27.365 109.995 -27.035 110.325 ;
        RECT -27.365 108.635 -27.035 108.965 ;
        RECT -27.365 107.275 -27.035 107.605 ;
        RECT -27.365 105.915 -27.035 106.245 ;
        RECT -27.365 104.555 -27.035 104.885 ;
        RECT -27.365 103.195 -27.035 103.525 ;
        RECT -27.365 101.835 -27.035 102.165 ;
        RECT -27.365 100.475 -27.035 100.805 ;
        RECT -27.365 99.115 -27.035 99.445 ;
        RECT -27.365 97.755 -27.035 98.085 ;
        RECT -27.365 96.395 -27.035 96.725 ;
        RECT -27.365 95.035 -27.035 95.365 ;
        RECT -27.365 93.675 -27.035 94.005 ;
        RECT -27.365 92.315 -27.035 92.645 ;
        RECT -27.365 90.955 -27.035 91.285 ;
        RECT -27.365 89.595 -27.035 89.925 ;
        RECT -27.365 88.235 -27.035 88.565 ;
        RECT -27.365 86.875 -27.035 87.205 ;
        RECT -27.365 85.515 -27.035 85.845 ;
        RECT -27.365 84.155 -27.035 84.485 ;
        RECT -27.365 82.795 -27.035 83.125 ;
        RECT -27.365 81.435 -27.035 81.765 ;
        RECT -27.365 80.075 -27.035 80.405 ;
        RECT -27.365 78.715 -27.035 79.045 ;
        RECT -27.365 77.355 -27.035 77.685 ;
        RECT -27.365 75.995 -27.035 76.325 ;
        RECT -27.365 74.635 -27.035 74.965 ;
        RECT -27.365 73.275 -27.035 73.605 ;
        RECT -27.365 71.915 -27.035 72.245 ;
        RECT -27.365 70.555 -27.035 70.885 ;
        RECT -27.365 69.195 -27.035 69.525 ;
        RECT -27.365 67.835 -27.035 68.165 ;
        RECT -27.365 66.475 -27.035 66.805 ;
        RECT -27.365 65.115 -27.035 65.445 ;
        RECT -27.365 63.755 -27.035 64.085 ;
        RECT -27.365 62.395 -27.035 62.725 ;
        RECT -27.365 61.035 -27.035 61.365 ;
        RECT -27.365 59.675 -27.035 60.005 ;
        RECT -27.365 58.315 -27.035 58.645 ;
        RECT -27.365 56.955 -27.035 57.285 ;
        RECT -27.365 55.595 -27.035 55.925 ;
        RECT -27.365 54.235 -27.035 54.565 ;
        RECT -27.365 52.875 -27.035 53.205 ;
        RECT -27.365 51.515 -27.035 51.845 ;
        RECT -27.365 50.155 -27.035 50.485 ;
        RECT -27.365 48.795 -27.035 49.125 ;
        RECT -27.365 47.435 -27.035 47.765 ;
        RECT -27.365 46.075 -27.035 46.405 ;
        RECT -27.365 44.715 -27.035 45.045 ;
        RECT -27.365 43.355 -27.035 43.685 ;
        RECT -27.365 41.995 -27.035 42.325 ;
        RECT -27.365 40.635 -27.035 40.965 ;
        RECT -27.365 39.275 -27.035 39.605 ;
        RECT -27.365 37.915 -27.035 38.245 ;
        RECT -27.365 36.555 -27.035 36.885 ;
        RECT -27.365 35.195 -27.035 35.525 ;
        RECT -27.365 33.835 -27.035 34.165 ;
        RECT -27.365 32.475 -27.035 32.805 ;
        RECT -27.365 31.115 -27.035 31.445 ;
        RECT -27.365 29.755 -27.035 30.085 ;
        RECT -27.365 28.395 -27.035 28.725 ;
        RECT -27.365 27.035 -27.035 27.365 ;
        RECT -27.365 25.675 -27.035 26.005 ;
        RECT -27.365 24.315 -27.035 24.645 ;
        RECT -27.365 22.955 -27.035 23.285 ;
        RECT -27.365 21.595 -27.035 21.925 ;
        RECT -27.365 20.235 -27.035 20.565 ;
        RECT -27.365 18.875 -27.035 19.205 ;
        RECT -27.365 17.515 -27.035 17.845 ;
        RECT -27.365 16.155 -27.035 16.485 ;
        RECT -27.365 14.795 -27.035 15.125 ;
        RECT -27.365 13.435 -27.035 13.765 ;
        RECT -27.365 12.075 -27.035 12.405 ;
        RECT -27.365 10.715 -27.035 11.045 ;
        RECT -27.365 9.355 -27.035 9.685 ;
        RECT -27.365 7.995 -27.035 8.325 ;
        RECT -27.365 6.635 -27.035 6.965 ;
        RECT -27.365 5.275 -27.035 5.605 ;
        RECT -27.365 3.915 -27.035 4.245 ;
        RECT -27.365 2.555 -27.035 2.885 ;
        RECT -27.365 1.195 -27.035 1.525 ;
        RECT -27.365 -0.165 -27.035 0.165 ;
        RECT -27.365 -8.325 -27.035 -7.995 ;
        RECT -27.365 -9.685 -27.035 -9.355 ;
        RECT -27.365 -14.95 -27.035 -14.62 ;
        RECT -27.365 -17.845 -27.035 -17.515 ;
        RECT -27.365 -19.79 -27.035 -19.46 ;
        RECT -27.365 -20.565 -27.035 -20.235 ;
        RECT -27.365 -28.725 -27.035 -28.395 ;
        RECT -27.365 -31.445 -27.035 -31.115 ;
        RECT -27.365 -32.805 -27.035 -32.475 ;
        RECT -27.365 -35.525 -27.035 -35.195 ;
        RECT -27.365 -36.885 -27.035 -36.555 ;
        RECT -27.365 -37.93 -27.035 -37.6 ;
        RECT -27.365 -40.965 -27.035 -40.635 ;
        RECT -27.365 -42.77 -27.035 -42.44 ;
        RECT -27.365 -43.685 -27.035 -43.355 ;
        RECT -27.365 -50.485 -27.035 -50.155 ;
        RECT -27.365 -51.845 -27.035 -51.515 ;
        RECT -27.365 -54.565 -27.035 -54.235 ;
        RECT -27.365 -55.925 -27.035 -55.595 ;
        RECT -27.365 -60.005 -27.035 -59.675 ;
        RECT -27.365 -66.805 -27.035 -66.475 ;
        RECT -27.365 -68.165 -27.035 -67.835 ;
        RECT -27.365 -69.525 -27.035 -69.195 ;
        RECT -27.365 -70.885 -27.035 -70.555 ;
        RECT -27.365 -72.245 -27.035 -71.915 ;
        RECT -27.365 -73.605 -27.035 -73.275 ;
        RECT -27.365 -74.965 -27.035 -74.635 ;
        RECT -27.365 -76.325 -27.035 -75.995 ;
        RECT -27.365 -77.685 -27.035 -77.355 ;
        RECT -27.365 -79.045 -27.035 -78.715 ;
        RECT -27.365 -80.405 -27.035 -80.075 ;
        RECT -27.365 -81.765 -27.035 -81.435 ;
        RECT -27.365 -83.125 -27.035 -82.795 ;
        RECT -27.365 -84.485 -27.035 -84.155 ;
        RECT -27.365 -85.845 -27.035 -85.515 ;
        RECT -27.365 -87.205 -27.035 -86.875 ;
        RECT -27.365 -88.565 -27.035 -88.235 ;
        RECT -27.365 -89.925 -27.035 -89.595 ;
        RECT -27.365 -92.645 -27.035 -92.315 ;
        RECT -27.365 -94.005 -27.035 -93.675 ;
        RECT -27.365 -95.365 -27.035 -95.035 ;
        RECT -27.365 -96.725 -27.035 -96.395 ;
        RECT -27.365 -98.73 -27.035 -98.4 ;
        RECT -27.365 -99.445 -27.035 -99.115 ;
        RECT -27.365 -102.165 -27.035 -101.835 ;
        RECT -27.365 -103.525 -27.035 -103.195 ;
        RECT -27.365 -104.885 -27.035 -104.555 ;
        RECT -27.365 -106.87 -27.035 -106.54 ;
        RECT -27.365 -107.605 -27.035 -107.275 ;
        RECT -27.365 -108.965 -27.035 -108.635 ;
        RECT -27.365 -113.045 -27.035 -112.715 ;
        RECT -27.365 -114.405 -27.035 -114.075 ;
        RECT -27.365 -115.765 -27.035 -115.435 ;
        RECT -27.365 -117.125 -27.035 -116.795 ;
        RECT -27.365 -118.485 -27.035 -118.155 ;
        RECT -27.365 -122.565 -27.035 -122.235 ;
        RECT -27.365 -125.285 -27.035 -124.955 ;
        RECT -27.365 -126.645 -27.035 -126.315 ;
        RECT -27.365 -128.005 -27.035 -127.675 ;
        RECT -27.365 -129.365 -27.035 -129.035 ;
        RECT -27.365 -133.445 -27.035 -133.115 ;
        RECT -27.365 -134.805 -27.035 -134.475 ;
        RECT -27.365 -136.165 -27.035 -135.835 ;
        RECT -27.365 -138.885 -27.035 -138.555 ;
        RECT -27.365 -141.605 -27.035 -141.275 ;
        RECT -27.365 -142.965 -27.035 -142.635 ;
        RECT -27.365 -144.325 -27.035 -143.995 ;
        RECT -27.365 -145.685 -27.035 -145.355 ;
        RECT -27.365 -147.045 -27.035 -146.715 ;
        RECT -27.365 -148.405 -27.035 -148.075 ;
        RECT -27.365 -151.125 -27.035 -150.795 ;
        RECT -27.365 -152.485 -27.035 -152.155 ;
        RECT -27.365 -156.565 -27.035 -156.235 ;
        RECT -27.365 -157.925 -27.035 -157.595 ;
        RECT -27.365 -159.285 -27.035 -158.955 ;
        RECT -27.365 -160.645 -27.035 -160.315 ;
        RECT -27.365 -162.005 -27.035 -161.675 ;
        RECT -27.365 -163.365 -27.035 -163.035 ;
        RECT -27.365 -164.725 -27.035 -164.395 ;
        RECT -27.365 -166.085 -27.035 -165.755 ;
        RECT -27.365 -167.445 -27.035 -167.115 ;
        RECT -27.365 -170.165 -27.035 -169.835 ;
        RECT -27.365 -174.245 -27.035 -173.915 ;
        RECT -27.365 -175.725 -27.035 -175.395 ;
        RECT -27.365 -176.965 -27.035 -176.635 ;
        RECT -27.365 -178.325 -27.035 -177.995 ;
        RECT -27.365 -180.57 -27.035 -179.44 ;
        RECT -27.36 -180.685 -27.04 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -26.005 241.32 -25.675 242.45 ;
        RECT -26.005 239.195 -25.675 239.525 ;
        RECT -26.005 237.835 -25.675 238.165 ;
        RECT -26.005 236.475 -25.675 236.805 ;
        RECT -26.005 235.115 -25.675 235.445 ;
        RECT -26.005 233.755 -25.675 234.085 ;
        RECT -26.005 232.395 -25.675 232.725 ;
        RECT -26.005 231.035 -25.675 231.365 ;
        RECT -26.005 229.675 -25.675 230.005 ;
        RECT -26.005 228.315 -25.675 228.645 ;
        RECT -26.005 226.955 -25.675 227.285 ;
        RECT -26.005 225.595 -25.675 225.925 ;
        RECT -26.005 224.235 -25.675 224.565 ;
        RECT -26.005 222.875 -25.675 223.205 ;
        RECT -26.005 221.515 -25.675 221.845 ;
        RECT -26.005 220.155 -25.675 220.485 ;
        RECT -26.005 218.795 -25.675 219.125 ;
        RECT -26.005 217.435 -25.675 217.765 ;
        RECT -26.005 216.075 -25.675 216.405 ;
        RECT -26.005 214.715 -25.675 215.045 ;
        RECT -26.005 213.355 -25.675 213.685 ;
        RECT -26.005 211.995 -25.675 212.325 ;
        RECT -26.005 210.635 -25.675 210.965 ;
        RECT -26.005 209.275 -25.675 209.605 ;
        RECT -26.005 207.915 -25.675 208.245 ;
        RECT -26.005 206.555 -25.675 206.885 ;
        RECT -26.005 205.195 -25.675 205.525 ;
        RECT -26.005 203.835 -25.675 204.165 ;
        RECT -26.005 202.475 -25.675 202.805 ;
        RECT -26.005 201.115 -25.675 201.445 ;
        RECT -26.005 199.755 -25.675 200.085 ;
        RECT -26.005 198.395 -25.675 198.725 ;
        RECT -26.005 197.035 -25.675 197.365 ;
        RECT -26.005 195.675 -25.675 196.005 ;
        RECT -26.005 194.315 -25.675 194.645 ;
        RECT -26.005 192.955 -25.675 193.285 ;
        RECT -26.005 191.595 -25.675 191.925 ;
        RECT -26.005 190.235 -25.675 190.565 ;
        RECT -26.005 188.875 -25.675 189.205 ;
        RECT -26.005 187.515 -25.675 187.845 ;
        RECT -26.005 186.155 -25.675 186.485 ;
        RECT -26.005 184.795 -25.675 185.125 ;
        RECT -26.005 183.435 -25.675 183.765 ;
        RECT -26.005 182.075 -25.675 182.405 ;
        RECT -26.005 180.715 -25.675 181.045 ;
        RECT -26.005 179.355 -25.675 179.685 ;
        RECT -26.005 177.995 -25.675 178.325 ;
        RECT -26.005 176.635 -25.675 176.965 ;
        RECT -26.005 175.275 -25.675 175.605 ;
        RECT -26.005 173.915 -25.675 174.245 ;
        RECT -26.005 172.555 -25.675 172.885 ;
        RECT -26.005 171.195 -25.675 171.525 ;
        RECT -26.005 169.835 -25.675 170.165 ;
        RECT -26.005 168.475 -25.675 168.805 ;
        RECT -26.005 167.115 -25.675 167.445 ;
        RECT -26.005 165.755 -25.675 166.085 ;
        RECT -26.005 164.395 -25.675 164.725 ;
        RECT -26.005 163.035 -25.675 163.365 ;
        RECT -26.005 161.675 -25.675 162.005 ;
        RECT -26.005 160.315 -25.675 160.645 ;
        RECT -26.005 158.955 -25.675 159.285 ;
        RECT -26.005 157.595 -25.675 157.925 ;
        RECT -26.005 156.235 -25.675 156.565 ;
        RECT -26.005 154.875 -25.675 155.205 ;
        RECT -26.005 153.515 -25.675 153.845 ;
        RECT -26.005 152.155 -25.675 152.485 ;
        RECT -26.005 150.795 -25.675 151.125 ;
        RECT -26.005 149.435 -25.675 149.765 ;
        RECT -26.005 148.075 -25.675 148.405 ;
        RECT -26.005 146.715 -25.675 147.045 ;
        RECT -26.005 145.355 -25.675 145.685 ;
        RECT -26.005 143.995 -25.675 144.325 ;
        RECT -26.005 142.635 -25.675 142.965 ;
        RECT -26.005 141.275 -25.675 141.605 ;
        RECT -26.005 139.915 -25.675 140.245 ;
        RECT -26.005 138.555 -25.675 138.885 ;
        RECT -26.005 137.195 -25.675 137.525 ;
        RECT -26.005 135.835 -25.675 136.165 ;
        RECT -26.005 134.475 -25.675 134.805 ;
        RECT -26.005 133.115 -25.675 133.445 ;
        RECT -26.005 131.755 -25.675 132.085 ;
        RECT -26.005 130.395 -25.675 130.725 ;
        RECT -26.005 129.035 -25.675 129.365 ;
        RECT -26.005 127.675 -25.675 128.005 ;
        RECT -26.005 126.315 -25.675 126.645 ;
        RECT -26.005 124.955 -25.675 125.285 ;
        RECT -26.005 123.595 -25.675 123.925 ;
        RECT -26.005 122.235 -25.675 122.565 ;
        RECT -26.005 120.875 -25.675 121.205 ;
        RECT -26.005 119.515 -25.675 119.845 ;
        RECT -26.005 118.155 -25.675 118.485 ;
        RECT -26.005 116.795 -25.675 117.125 ;
        RECT -26.005 115.435 -25.675 115.765 ;
        RECT -26.005 114.075 -25.675 114.405 ;
        RECT -26.005 112.715 -25.675 113.045 ;
        RECT -26.005 111.355 -25.675 111.685 ;
        RECT -26.005 109.995 -25.675 110.325 ;
        RECT -26.005 108.635 -25.675 108.965 ;
        RECT -26.005 107.275 -25.675 107.605 ;
        RECT -26.005 105.915 -25.675 106.245 ;
        RECT -26.005 104.555 -25.675 104.885 ;
        RECT -26.005 103.195 -25.675 103.525 ;
        RECT -26.005 101.835 -25.675 102.165 ;
        RECT -26.005 100.475 -25.675 100.805 ;
        RECT -26.005 99.115 -25.675 99.445 ;
        RECT -26.005 97.755 -25.675 98.085 ;
        RECT -26.005 96.395 -25.675 96.725 ;
        RECT -26.005 95.035 -25.675 95.365 ;
        RECT -26.005 93.675 -25.675 94.005 ;
        RECT -26.005 92.315 -25.675 92.645 ;
        RECT -26.005 90.955 -25.675 91.285 ;
        RECT -26.005 89.595 -25.675 89.925 ;
        RECT -26.005 88.235 -25.675 88.565 ;
        RECT -26.005 86.875 -25.675 87.205 ;
        RECT -26.005 85.515 -25.675 85.845 ;
        RECT -26.005 84.155 -25.675 84.485 ;
        RECT -26.005 82.795 -25.675 83.125 ;
        RECT -26.005 81.435 -25.675 81.765 ;
        RECT -26.005 80.075 -25.675 80.405 ;
        RECT -26.005 78.715 -25.675 79.045 ;
        RECT -26.005 77.355 -25.675 77.685 ;
        RECT -26.005 75.995 -25.675 76.325 ;
        RECT -26.005 74.635 -25.675 74.965 ;
        RECT -26.005 73.275 -25.675 73.605 ;
        RECT -26.005 71.915 -25.675 72.245 ;
        RECT -26.005 70.555 -25.675 70.885 ;
        RECT -26.005 69.195 -25.675 69.525 ;
        RECT -26.005 67.835 -25.675 68.165 ;
        RECT -26.005 66.475 -25.675 66.805 ;
        RECT -26.005 65.115 -25.675 65.445 ;
        RECT -26.005 63.755 -25.675 64.085 ;
        RECT -26.005 62.395 -25.675 62.725 ;
        RECT -26.005 61.035 -25.675 61.365 ;
        RECT -26.005 59.675 -25.675 60.005 ;
        RECT -26.005 58.315 -25.675 58.645 ;
        RECT -26.005 56.955 -25.675 57.285 ;
        RECT -26.005 55.595 -25.675 55.925 ;
        RECT -26.005 54.235 -25.675 54.565 ;
        RECT -26.005 52.875 -25.675 53.205 ;
        RECT -26.005 51.515 -25.675 51.845 ;
        RECT -26.005 50.155 -25.675 50.485 ;
        RECT -26.005 48.795 -25.675 49.125 ;
        RECT -26.005 47.435 -25.675 47.765 ;
        RECT -26.005 46.075 -25.675 46.405 ;
        RECT -26.005 44.715 -25.675 45.045 ;
        RECT -26.005 43.355 -25.675 43.685 ;
        RECT -26.005 41.995 -25.675 42.325 ;
        RECT -26.005 40.635 -25.675 40.965 ;
        RECT -26.005 39.275 -25.675 39.605 ;
        RECT -26.005 37.915 -25.675 38.245 ;
        RECT -26.005 36.555 -25.675 36.885 ;
        RECT -26.005 35.195 -25.675 35.525 ;
        RECT -26.005 33.835 -25.675 34.165 ;
        RECT -26.005 32.475 -25.675 32.805 ;
        RECT -26.005 31.115 -25.675 31.445 ;
        RECT -26.005 29.755 -25.675 30.085 ;
        RECT -26.005 28.395 -25.675 28.725 ;
        RECT -26.005 27.035 -25.675 27.365 ;
        RECT -26.005 25.675 -25.675 26.005 ;
        RECT -26.005 24.315 -25.675 24.645 ;
        RECT -26.005 22.955 -25.675 23.285 ;
        RECT -26.005 21.595 -25.675 21.925 ;
        RECT -26.005 20.235 -25.675 20.565 ;
        RECT -26.005 18.875 -25.675 19.205 ;
        RECT -26.005 17.515 -25.675 17.845 ;
        RECT -26.005 16.155 -25.675 16.485 ;
        RECT -26.005 14.795 -25.675 15.125 ;
        RECT -26.005 13.435 -25.675 13.765 ;
        RECT -26.005 12.075 -25.675 12.405 ;
        RECT -26.005 10.715 -25.675 11.045 ;
        RECT -26.005 9.355 -25.675 9.685 ;
        RECT -26.005 7.995 -25.675 8.325 ;
        RECT -26.005 6.635 -25.675 6.965 ;
        RECT -26.005 5.275 -25.675 5.605 ;
        RECT -26.005 3.915 -25.675 4.245 ;
        RECT -26.005 2.555 -25.675 2.885 ;
        RECT -26.005 1.195 -25.675 1.525 ;
        RECT -26.005 -0.165 -25.675 0.165 ;
        RECT -26.005 -2.885 -25.675 -2.555 ;
        RECT -26.005 -8.325 -25.675 -7.995 ;
        RECT -26.005 -9.685 -25.675 -9.355 ;
        RECT -26.005 -14.95 -25.675 -14.62 ;
        RECT -26.005 -17.845 -25.675 -17.515 ;
        RECT -26.005 -19.79 -25.675 -19.46 ;
        RECT -26.005 -20.565 -25.675 -20.235 ;
        RECT -26.005 -28.725 -25.675 -28.395 ;
        RECT -26.005 -31.445 -25.675 -31.115 ;
        RECT -26.005 -32.805 -25.675 -32.475 ;
        RECT -26.005 -35.525 -25.675 -35.195 ;
        RECT -26.005 -36.885 -25.675 -36.555 ;
        RECT -26.005 -37.93 -25.675 -37.6 ;
        RECT -26.005 -40.965 -25.675 -40.635 ;
        RECT -26.005 -42.77 -25.675 -42.44 ;
        RECT -26.005 -43.685 -25.675 -43.355 ;
        RECT -26.005 -50.485 -25.675 -50.155 ;
        RECT -26.005 -51.845 -25.675 -51.515 ;
        RECT -26.005 -54.565 -25.675 -54.235 ;
        RECT -26.005 -55.925 -25.675 -55.595 ;
        RECT -26.005 -60.005 -25.675 -59.675 ;
        RECT -26.005 -66.805 -25.675 -66.475 ;
        RECT -26.005 -68.165 -25.675 -67.835 ;
        RECT -26.005 -69.525 -25.675 -69.195 ;
        RECT -26.005 -70.885 -25.675 -70.555 ;
        RECT -26.005 -72.245 -25.675 -71.915 ;
        RECT -26.005 -73.605 -25.675 -73.275 ;
        RECT -26.005 -74.965 -25.675 -74.635 ;
        RECT -26.005 -76.325 -25.675 -75.995 ;
        RECT -26.005 -77.685 -25.675 -77.355 ;
        RECT -26.005 -79.045 -25.675 -78.715 ;
        RECT -26.005 -80.405 -25.675 -80.075 ;
        RECT -26.005 -81.765 -25.675 -81.435 ;
        RECT -26.005 -83.125 -25.675 -82.795 ;
        RECT -26.005 -84.485 -25.675 -84.155 ;
        RECT -26.005 -85.845 -25.675 -85.515 ;
        RECT -26.005 -87.205 -25.675 -86.875 ;
        RECT -26.005 -88.565 -25.675 -88.235 ;
        RECT -26.005 -89.925 -25.675 -89.595 ;
        RECT -26.005 -91.285 -25.675 -90.955 ;
        RECT -26.005 -92.645 -25.675 -92.315 ;
        RECT -26.005 -94.005 -25.675 -93.675 ;
        RECT -26.005 -95.365 -25.675 -95.035 ;
        RECT -26.005 -96.725 -25.675 -96.395 ;
        RECT -26.005 -98.085 -25.675 -97.755 ;
        RECT -26.005 -99.445 -25.675 -99.115 ;
        RECT -26.005 -100.805 -25.675 -100.475 ;
        RECT -26.005 -102.165 -25.675 -101.835 ;
        RECT -26.005 -103.525 -25.675 -103.195 ;
        RECT -26.005 -104.885 -25.675 -104.555 ;
        RECT -26.005 -106.245 -25.675 -105.915 ;
        RECT -26.005 -107.605 -25.675 -107.275 ;
        RECT -26.005 -108.965 -25.675 -108.635 ;
        RECT -26.005 -111.685 -25.675 -111.355 ;
        RECT -26.005 -113.045 -25.675 -112.715 ;
        RECT -26.005 -114.405 -25.675 -114.075 ;
        RECT -26.005 -115.765 -25.675 -115.435 ;
        RECT -26.005 -117.125 -25.675 -116.795 ;
        RECT -26.005 -118.485 -25.675 -118.155 ;
        RECT -26.005 -122.565 -25.675 -122.235 ;
        RECT -26.005 -123.925 -25.675 -123.595 ;
        RECT -26.005 -125.285 -25.675 -124.955 ;
        RECT -26.005 -126.645 -25.675 -126.315 ;
        RECT -26.005 -128.005 -25.675 -127.675 ;
        RECT -26.005 -129.365 -25.675 -129.035 ;
        RECT -26.005 -133.445 -25.675 -133.115 ;
        RECT -26.005 -134.805 -25.675 -134.475 ;
        RECT -26.005 -136.165 -25.675 -135.835 ;
        RECT -26.005 -138.885 -25.675 -138.555 ;
        RECT -26.005 -141.605 -25.675 -141.275 ;
        RECT -26.005 -142.965 -25.675 -142.635 ;
        RECT -26.005 -144.325 -25.675 -143.995 ;
        RECT -26.005 -145.685 -25.675 -145.355 ;
        RECT -26.005 -147.045 -25.675 -146.715 ;
        RECT -26.005 -148.405 -25.675 -148.075 ;
        RECT -26.005 -151.125 -25.675 -150.795 ;
        RECT -26.005 -152.485 -25.675 -152.155 ;
        RECT -26.005 -156.565 -25.675 -156.235 ;
        RECT -26.005 -157.925 -25.675 -157.595 ;
        RECT -26.005 -159.285 -25.675 -158.955 ;
        RECT -26.005 -160.645 -25.675 -160.315 ;
        RECT -26.005 -162.005 -25.675 -161.675 ;
        RECT -26.005 -163.365 -25.675 -163.035 ;
        RECT -26.005 -164.725 -25.675 -164.395 ;
        RECT -26.005 -166.085 -25.675 -165.755 ;
        RECT -26.005 -167.445 -25.675 -167.115 ;
        RECT -26.005 -170.165 -25.675 -169.835 ;
        RECT -26.005 -172.885 -25.675 -172.555 ;
        RECT -26.005 -174.245 -25.675 -173.915 ;
        RECT -26.005 -175.725 -25.675 -175.395 ;
        RECT -26.005 -176.965 -25.675 -176.635 ;
        RECT -26.005 -178.325 -25.675 -177.995 ;
        RECT -26.005 -180.57 -25.675 -179.44 ;
        RECT -26 -180.685 -25.68 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -24.645 172.555 -24.315 172.885 ;
        RECT -24.645 171.195 -24.315 171.525 ;
        RECT -24.645 169.835 -24.315 170.165 ;
        RECT -24.645 168.475 -24.315 168.805 ;
        RECT -24.645 167.115 -24.315 167.445 ;
        RECT -24.645 165.755 -24.315 166.085 ;
        RECT -24.645 164.395 -24.315 164.725 ;
        RECT -24.645 163.035 -24.315 163.365 ;
        RECT -24.645 161.675 -24.315 162.005 ;
        RECT -24.645 160.315 -24.315 160.645 ;
        RECT -24.645 158.955 -24.315 159.285 ;
        RECT -24.645 157.595 -24.315 157.925 ;
        RECT -24.645 156.235 -24.315 156.565 ;
        RECT -24.645 154.875 -24.315 155.205 ;
        RECT -24.645 153.515 -24.315 153.845 ;
        RECT -24.645 152.155 -24.315 152.485 ;
        RECT -24.645 150.795 -24.315 151.125 ;
        RECT -24.645 149.435 -24.315 149.765 ;
        RECT -24.645 148.075 -24.315 148.405 ;
        RECT -24.645 146.715 -24.315 147.045 ;
        RECT -24.645 145.355 -24.315 145.685 ;
        RECT -24.645 143.995 -24.315 144.325 ;
        RECT -24.645 142.635 -24.315 142.965 ;
        RECT -24.645 141.275 -24.315 141.605 ;
        RECT -24.645 139.915 -24.315 140.245 ;
        RECT -24.645 138.555 -24.315 138.885 ;
        RECT -24.645 137.195 -24.315 137.525 ;
        RECT -24.645 135.835 -24.315 136.165 ;
        RECT -24.645 134.475 -24.315 134.805 ;
        RECT -24.645 133.115 -24.315 133.445 ;
        RECT -24.645 131.755 -24.315 132.085 ;
        RECT -24.645 130.395 -24.315 130.725 ;
        RECT -24.645 129.035 -24.315 129.365 ;
        RECT -24.645 127.675 -24.315 128.005 ;
        RECT -24.645 126.315 -24.315 126.645 ;
        RECT -24.645 124.955 -24.315 125.285 ;
        RECT -24.645 123.595 -24.315 123.925 ;
        RECT -24.645 122.235 -24.315 122.565 ;
        RECT -24.645 120.875 -24.315 121.205 ;
        RECT -24.645 119.515 -24.315 119.845 ;
        RECT -24.645 118.155 -24.315 118.485 ;
        RECT -24.645 116.795 -24.315 117.125 ;
        RECT -24.645 115.435 -24.315 115.765 ;
        RECT -24.645 114.075 -24.315 114.405 ;
        RECT -24.645 112.715 -24.315 113.045 ;
        RECT -24.645 111.355 -24.315 111.685 ;
        RECT -24.645 109.995 -24.315 110.325 ;
        RECT -24.645 108.635 -24.315 108.965 ;
        RECT -24.645 107.275 -24.315 107.605 ;
        RECT -24.645 105.915 -24.315 106.245 ;
        RECT -24.645 104.555 -24.315 104.885 ;
        RECT -24.645 103.195 -24.315 103.525 ;
        RECT -24.645 101.835 -24.315 102.165 ;
        RECT -24.645 100.475 -24.315 100.805 ;
        RECT -24.645 99.115 -24.315 99.445 ;
        RECT -24.645 97.755 -24.315 98.085 ;
        RECT -24.645 96.395 -24.315 96.725 ;
        RECT -24.645 95.035 -24.315 95.365 ;
        RECT -24.645 93.675 -24.315 94.005 ;
        RECT -24.645 92.315 -24.315 92.645 ;
        RECT -24.645 90.955 -24.315 91.285 ;
        RECT -24.645 89.595 -24.315 89.925 ;
        RECT -24.645 88.235 -24.315 88.565 ;
        RECT -24.645 86.875 -24.315 87.205 ;
        RECT -24.645 85.515 -24.315 85.845 ;
        RECT -24.645 84.155 -24.315 84.485 ;
        RECT -24.645 82.795 -24.315 83.125 ;
        RECT -24.645 81.435 -24.315 81.765 ;
        RECT -24.645 80.075 -24.315 80.405 ;
        RECT -24.645 78.715 -24.315 79.045 ;
        RECT -24.645 77.355 -24.315 77.685 ;
        RECT -24.645 75.995 -24.315 76.325 ;
        RECT -24.645 74.635 -24.315 74.965 ;
        RECT -24.645 73.275 -24.315 73.605 ;
        RECT -24.645 71.915 -24.315 72.245 ;
        RECT -24.645 70.555 -24.315 70.885 ;
        RECT -24.645 69.195 -24.315 69.525 ;
        RECT -24.645 67.835 -24.315 68.165 ;
        RECT -24.645 66.475 -24.315 66.805 ;
        RECT -24.645 65.115 -24.315 65.445 ;
        RECT -24.645 63.755 -24.315 64.085 ;
        RECT -24.645 62.395 -24.315 62.725 ;
        RECT -24.645 61.035 -24.315 61.365 ;
        RECT -24.645 59.675 -24.315 60.005 ;
        RECT -24.645 58.315 -24.315 58.645 ;
        RECT -24.645 56.955 -24.315 57.285 ;
        RECT -24.645 55.595 -24.315 55.925 ;
        RECT -24.645 54.235 -24.315 54.565 ;
        RECT -24.645 52.875 -24.315 53.205 ;
        RECT -24.645 51.515 -24.315 51.845 ;
        RECT -24.645 50.155 -24.315 50.485 ;
        RECT -24.645 48.795 -24.315 49.125 ;
        RECT -24.645 47.435 -24.315 47.765 ;
        RECT -24.645 46.075 -24.315 46.405 ;
        RECT -24.645 44.715 -24.315 45.045 ;
        RECT -24.645 43.355 -24.315 43.685 ;
        RECT -24.645 41.995 -24.315 42.325 ;
        RECT -24.645 40.635 -24.315 40.965 ;
        RECT -24.645 39.275 -24.315 39.605 ;
        RECT -24.645 37.915 -24.315 38.245 ;
        RECT -24.645 36.555 -24.315 36.885 ;
        RECT -24.645 35.195 -24.315 35.525 ;
        RECT -24.645 33.835 -24.315 34.165 ;
        RECT -24.645 32.475 -24.315 32.805 ;
        RECT -24.645 31.115 -24.315 31.445 ;
        RECT -24.645 29.755 -24.315 30.085 ;
        RECT -24.645 28.395 -24.315 28.725 ;
        RECT -24.645 27.035 -24.315 27.365 ;
        RECT -24.645 25.675 -24.315 26.005 ;
        RECT -24.645 24.315 -24.315 24.645 ;
        RECT -24.645 22.955 -24.315 23.285 ;
        RECT -24.645 21.595 -24.315 21.925 ;
        RECT -24.645 20.235 -24.315 20.565 ;
        RECT -24.645 18.875 -24.315 19.205 ;
        RECT -24.645 17.515 -24.315 17.845 ;
        RECT -24.645 16.155 -24.315 16.485 ;
        RECT -24.645 14.795 -24.315 15.125 ;
        RECT -24.645 13.435 -24.315 13.765 ;
        RECT -24.645 12.075 -24.315 12.405 ;
        RECT -24.645 10.715 -24.315 11.045 ;
        RECT -24.645 9.355 -24.315 9.685 ;
        RECT -24.645 7.995 -24.315 8.325 ;
        RECT -24.645 6.635 -24.315 6.965 ;
        RECT -24.645 5.275 -24.315 5.605 ;
        RECT -24.645 3.915 -24.315 4.245 ;
        RECT -24.645 2.555 -24.315 2.885 ;
        RECT -24.645 1.195 -24.315 1.525 ;
        RECT -24.645 -0.165 -24.315 0.165 ;
        RECT -24.645 -2.885 -24.315 -2.555 ;
        RECT -24.645 -8.325 -24.315 -7.995 ;
        RECT -24.645 -9.685 -24.315 -9.355 ;
        RECT -24.645 -14.95 -24.315 -14.62 ;
        RECT -24.645 -17.845 -24.315 -17.515 ;
        RECT -24.645 -19.79 -24.315 -19.46 ;
        RECT -24.645 -20.565 -24.315 -20.235 ;
        RECT -24.645 -28.725 -24.315 -28.395 ;
        RECT -24.645 -31.445 -24.315 -31.115 ;
        RECT -24.645 -32.805 -24.315 -32.475 ;
        RECT -24.645 -35.525 -24.315 -35.195 ;
        RECT -24.645 -36.885 -24.315 -36.555 ;
        RECT -24.645 -37.93 -24.315 -37.6 ;
        RECT -24.645 -40.965 -24.315 -40.635 ;
        RECT -24.645 -42.77 -24.315 -42.44 ;
        RECT -24.645 -43.685 -24.315 -43.355 ;
        RECT -24.645 -50.485 -24.315 -50.155 ;
        RECT -24.645 -51.845 -24.315 -51.515 ;
        RECT -24.645 -54.565 -24.315 -54.235 ;
        RECT -24.645 -55.925 -24.315 -55.595 ;
        RECT -24.645 -60.005 -24.315 -59.675 ;
        RECT -24.645 -66.805 -24.315 -66.475 ;
        RECT -24.645 -68.165 -24.315 -67.835 ;
        RECT -24.645 -69.525 -24.315 -69.195 ;
        RECT -24.645 -70.885 -24.315 -70.555 ;
        RECT -24.645 -72.245 -24.315 -71.915 ;
        RECT -24.645 -73.605 -24.315 -73.275 ;
        RECT -24.645 -74.965 -24.315 -74.635 ;
        RECT -24.645 -76.325 -24.315 -75.995 ;
        RECT -24.645 -77.685 -24.315 -77.355 ;
        RECT -24.645 -79.045 -24.315 -78.715 ;
        RECT -24.645 -80.405 -24.315 -80.075 ;
        RECT -24.645 -81.765 -24.315 -81.435 ;
        RECT -24.645 -83.125 -24.315 -82.795 ;
        RECT -24.645 -84.485 -24.315 -84.155 ;
        RECT -24.645 -85.845 -24.315 -85.515 ;
        RECT -24.645 -87.205 -24.315 -86.875 ;
        RECT -24.645 -88.565 -24.315 -88.235 ;
        RECT -24.645 -89.925 -24.315 -89.595 ;
        RECT -24.645 -91.285 -24.315 -90.955 ;
        RECT -24.645 -92.645 -24.315 -92.315 ;
        RECT -24.645 -94.005 -24.315 -93.675 ;
        RECT -24.645 -95.365 -24.315 -95.035 ;
        RECT -24.645 -96.725 -24.315 -96.395 ;
        RECT -24.645 -98.085 -24.315 -97.755 ;
        RECT -24.645 -99.445 -24.315 -99.115 ;
        RECT -24.645 -100.805 -24.315 -100.475 ;
        RECT -24.645 -102.165 -24.315 -101.835 ;
        RECT -24.645 -103.525 -24.315 -103.195 ;
        RECT -24.645 -104.885 -24.315 -104.555 ;
        RECT -24.645 -106.245 -24.315 -105.915 ;
        RECT -24.645 -107.605 -24.315 -107.275 ;
        RECT -24.645 -108.965 -24.315 -108.635 ;
        RECT -24.645 -111.685 -24.315 -111.355 ;
        RECT -24.645 -113.045 -24.315 -112.715 ;
        RECT -24.645 -114.405 -24.315 -114.075 ;
        RECT -24.645 -115.765 -24.315 -115.435 ;
        RECT -24.645 -117.125 -24.315 -116.795 ;
        RECT -24.645 -118.485 -24.315 -118.155 ;
        RECT -24.645 -122.565 -24.315 -122.235 ;
        RECT -24.645 -123.925 -24.315 -123.595 ;
        RECT -24.645 -125.285 -24.315 -124.955 ;
        RECT -24.645 -126.645 -24.315 -126.315 ;
        RECT -24.645 -128.005 -24.315 -127.675 ;
        RECT -24.645 -133.445 -24.315 -133.115 ;
        RECT -24.645 -134.805 -24.315 -134.475 ;
        RECT -24.645 -136.165 -24.315 -135.835 ;
        RECT -24.645 -138.885 -24.315 -138.555 ;
        RECT -24.645 -141.605 -24.315 -141.275 ;
        RECT -24.645 -142.965 -24.315 -142.635 ;
        RECT -24.645 -145.685 -24.315 -145.355 ;
        RECT -24.645 -147.045 -24.315 -146.715 ;
        RECT -24.645 -148.405 -24.315 -148.075 ;
        RECT -24.645 -151.125 -24.315 -150.795 ;
        RECT -24.645 -152.485 -24.315 -152.155 ;
        RECT -24.645 -157.925 -24.315 -157.595 ;
        RECT -24.645 -159.285 -24.315 -158.955 ;
        RECT -24.645 -160.645 -24.315 -160.315 ;
        RECT -24.645 -162.005 -24.315 -161.675 ;
        RECT -24.645 -163.365 -24.315 -163.035 ;
        RECT -24.645 -164.725 -24.315 -164.395 ;
        RECT -24.645 -166.085 -24.315 -165.755 ;
        RECT -24.645 -167.445 -24.315 -167.115 ;
        RECT -24.645 -170.165 -24.315 -169.835 ;
        RECT -24.645 -172.885 -24.315 -172.555 ;
        RECT -24.645 -174.245 -24.315 -173.915 ;
        RECT -24.645 -175.725 -24.315 -175.395 ;
        RECT -24.645 -176.965 -24.315 -176.635 ;
        RECT -24.645 -178.325 -24.315 -177.995 ;
        RECT -24.645 -180.57 -24.315 -179.44 ;
        RECT -24.64 -180.685 -24.32 242.565 ;
        RECT -24.645 241.32 -24.315 242.45 ;
        RECT -24.645 239.195 -24.315 239.525 ;
        RECT -24.645 237.835 -24.315 238.165 ;
        RECT -24.645 236.475 -24.315 236.805 ;
        RECT -24.645 235.115 -24.315 235.445 ;
        RECT -24.645 233.755 -24.315 234.085 ;
        RECT -24.645 232.395 -24.315 232.725 ;
        RECT -24.645 231.035 -24.315 231.365 ;
        RECT -24.645 229.675 -24.315 230.005 ;
        RECT -24.645 228.315 -24.315 228.645 ;
        RECT -24.645 226.955 -24.315 227.285 ;
        RECT -24.645 225.595 -24.315 225.925 ;
        RECT -24.645 224.235 -24.315 224.565 ;
        RECT -24.645 222.875 -24.315 223.205 ;
        RECT -24.645 221.515 -24.315 221.845 ;
        RECT -24.645 220.155 -24.315 220.485 ;
        RECT -24.645 218.795 -24.315 219.125 ;
        RECT -24.645 217.435 -24.315 217.765 ;
        RECT -24.645 216.075 -24.315 216.405 ;
        RECT -24.645 214.715 -24.315 215.045 ;
        RECT -24.645 213.355 -24.315 213.685 ;
        RECT -24.645 211.995 -24.315 212.325 ;
        RECT -24.645 210.635 -24.315 210.965 ;
        RECT -24.645 209.275 -24.315 209.605 ;
        RECT -24.645 207.915 -24.315 208.245 ;
        RECT -24.645 206.555 -24.315 206.885 ;
        RECT -24.645 205.195 -24.315 205.525 ;
        RECT -24.645 203.835 -24.315 204.165 ;
        RECT -24.645 202.475 -24.315 202.805 ;
        RECT -24.645 201.115 -24.315 201.445 ;
        RECT -24.645 199.755 -24.315 200.085 ;
        RECT -24.645 198.395 -24.315 198.725 ;
        RECT -24.645 197.035 -24.315 197.365 ;
        RECT -24.645 195.675 -24.315 196.005 ;
        RECT -24.645 194.315 -24.315 194.645 ;
        RECT -24.645 192.955 -24.315 193.285 ;
        RECT -24.645 191.595 -24.315 191.925 ;
        RECT -24.645 190.235 -24.315 190.565 ;
        RECT -24.645 188.875 -24.315 189.205 ;
        RECT -24.645 187.515 -24.315 187.845 ;
        RECT -24.645 186.155 -24.315 186.485 ;
        RECT -24.645 184.795 -24.315 185.125 ;
        RECT -24.645 183.435 -24.315 183.765 ;
        RECT -24.645 182.075 -24.315 182.405 ;
        RECT -24.645 180.715 -24.315 181.045 ;
        RECT -24.645 179.355 -24.315 179.685 ;
        RECT -24.645 177.995 -24.315 178.325 ;
        RECT -24.645 176.635 -24.315 176.965 ;
        RECT -24.645 175.275 -24.315 175.605 ;
        RECT -24.645 173.915 -24.315 174.245 ;
    END
    PORT
      LAYER met3 ;
        RECT -32.805 241.32 -32.475 242.45 ;
        RECT -32.805 239.195 -32.475 239.525 ;
        RECT -32.805 237.835 -32.475 238.165 ;
        RECT -32.805 236.475 -32.475 236.805 ;
        RECT -32.805 235.115 -32.475 235.445 ;
        RECT -32.805 233.755 -32.475 234.085 ;
        RECT -32.805 232.395 -32.475 232.725 ;
        RECT -32.805 231.035 -32.475 231.365 ;
        RECT -32.805 229.675 -32.475 230.005 ;
        RECT -32.805 228.315 -32.475 228.645 ;
        RECT -32.805 226.955 -32.475 227.285 ;
        RECT -32.805 225.595 -32.475 225.925 ;
        RECT -32.805 224.235 -32.475 224.565 ;
        RECT -32.805 222.875 -32.475 223.205 ;
        RECT -32.805 221.515 -32.475 221.845 ;
        RECT -32.805 220.155 -32.475 220.485 ;
        RECT -32.805 218.795 -32.475 219.125 ;
        RECT -32.805 217.435 -32.475 217.765 ;
        RECT -32.805 216.075 -32.475 216.405 ;
        RECT -32.805 214.715 -32.475 215.045 ;
        RECT -32.805 213.355 -32.475 213.685 ;
        RECT -32.805 211.995 -32.475 212.325 ;
        RECT -32.805 210.635 -32.475 210.965 ;
        RECT -32.805 209.275 -32.475 209.605 ;
        RECT -32.805 207.915 -32.475 208.245 ;
        RECT -32.805 206.555 -32.475 206.885 ;
        RECT -32.805 205.195 -32.475 205.525 ;
        RECT -32.805 203.835 -32.475 204.165 ;
        RECT -32.805 202.475 -32.475 202.805 ;
        RECT -32.805 201.115 -32.475 201.445 ;
        RECT -32.805 199.755 -32.475 200.085 ;
        RECT -32.805 198.395 -32.475 198.725 ;
        RECT -32.805 197.035 -32.475 197.365 ;
        RECT -32.805 195.675 -32.475 196.005 ;
        RECT -32.805 194.315 -32.475 194.645 ;
        RECT -32.805 192.955 -32.475 193.285 ;
        RECT -32.805 191.595 -32.475 191.925 ;
        RECT -32.805 190.235 -32.475 190.565 ;
        RECT -32.805 188.875 -32.475 189.205 ;
        RECT -32.805 187.515 -32.475 187.845 ;
        RECT -32.805 186.155 -32.475 186.485 ;
        RECT -32.805 184.795 -32.475 185.125 ;
        RECT -32.805 183.435 -32.475 183.765 ;
        RECT -32.805 182.075 -32.475 182.405 ;
        RECT -32.805 180.715 -32.475 181.045 ;
        RECT -32.805 179.355 -32.475 179.685 ;
        RECT -32.805 177.995 -32.475 178.325 ;
        RECT -32.805 176.635 -32.475 176.965 ;
        RECT -32.805 175.275 -32.475 175.605 ;
        RECT -32.805 173.915 -32.475 174.245 ;
        RECT -32.805 172.555 -32.475 172.885 ;
        RECT -32.805 171.195 -32.475 171.525 ;
        RECT -32.805 169.835 -32.475 170.165 ;
        RECT -32.805 168.475 -32.475 168.805 ;
        RECT -32.805 167.115 -32.475 167.445 ;
        RECT -32.805 165.755 -32.475 166.085 ;
        RECT -32.805 164.395 -32.475 164.725 ;
        RECT -32.805 163.035 -32.475 163.365 ;
        RECT -32.805 161.675 -32.475 162.005 ;
        RECT -32.805 160.315 -32.475 160.645 ;
        RECT -32.805 158.955 -32.475 159.285 ;
        RECT -32.805 157.595 -32.475 157.925 ;
        RECT -32.805 156.235 -32.475 156.565 ;
        RECT -32.805 154.875 -32.475 155.205 ;
        RECT -32.805 153.515 -32.475 153.845 ;
        RECT -32.805 152.155 -32.475 152.485 ;
        RECT -32.805 150.795 -32.475 151.125 ;
        RECT -32.805 149.435 -32.475 149.765 ;
        RECT -32.805 148.075 -32.475 148.405 ;
        RECT -32.805 146.715 -32.475 147.045 ;
        RECT -32.805 145.355 -32.475 145.685 ;
        RECT -32.805 143.995 -32.475 144.325 ;
        RECT -32.805 142.635 -32.475 142.965 ;
        RECT -32.805 141.275 -32.475 141.605 ;
        RECT -32.805 139.915 -32.475 140.245 ;
        RECT -32.805 138.555 -32.475 138.885 ;
        RECT -32.805 137.195 -32.475 137.525 ;
        RECT -32.805 135.835 -32.475 136.165 ;
        RECT -32.805 134.475 -32.475 134.805 ;
        RECT -32.805 133.115 -32.475 133.445 ;
        RECT -32.805 131.755 -32.475 132.085 ;
        RECT -32.805 130.395 -32.475 130.725 ;
        RECT -32.805 129.035 -32.475 129.365 ;
        RECT -32.805 127.675 -32.475 128.005 ;
        RECT -32.805 126.315 -32.475 126.645 ;
        RECT -32.805 124.955 -32.475 125.285 ;
        RECT -32.805 123.595 -32.475 123.925 ;
        RECT -32.805 122.235 -32.475 122.565 ;
        RECT -32.805 120.875 -32.475 121.205 ;
        RECT -32.805 119.515 -32.475 119.845 ;
        RECT -32.805 118.155 -32.475 118.485 ;
        RECT -32.805 116.795 -32.475 117.125 ;
        RECT -32.805 115.435 -32.475 115.765 ;
        RECT -32.805 114.075 -32.475 114.405 ;
        RECT -32.805 112.715 -32.475 113.045 ;
        RECT -32.805 111.355 -32.475 111.685 ;
        RECT -32.805 109.995 -32.475 110.325 ;
        RECT -32.805 108.635 -32.475 108.965 ;
        RECT -32.805 107.275 -32.475 107.605 ;
        RECT -32.805 105.915 -32.475 106.245 ;
        RECT -32.805 104.555 -32.475 104.885 ;
        RECT -32.805 103.195 -32.475 103.525 ;
        RECT -32.805 101.835 -32.475 102.165 ;
        RECT -32.805 100.475 -32.475 100.805 ;
        RECT -32.805 99.115 -32.475 99.445 ;
        RECT -32.805 97.755 -32.475 98.085 ;
        RECT -32.805 96.395 -32.475 96.725 ;
        RECT -32.805 95.035 -32.475 95.365 ;
        RECT -32.805 93.675 -32.475 94.005 ;
        RECT -32.805 92.315 -32.475 92.645 ;
        RECT -32.805 90.955 -32.475 91.285 ;
        RECT -32.805 89.595 -32.475 89.925 ;
        RECT -32.805 88.235 -32.475 88.565 ;
        RECT -32.805 86.875 -32.475 87.205 ;
        RECT -32.805 85.515 -32.475 85.845 ;
        RECT -32.805 84.155 -32.475 84.485 ;
        RECT -32.805 82.795 -32.475 83.125 ;
        RECT -32.805 81.435 -32.475 81.765 ;
        RECT -32.805 80.075 -32.475 80.405 ;
        RECT -32.805 78.715 -32.475 79.045 ;
        RECT -32.805 77.355 -32.475 77.685 ;
        RECT -32.805 75.995 -32.475 76.325 ;
        RECT -32.805 74.635 -32.475 74.965 ;
        RECT -32.805 73.275 -32.475 73.605 ;
        RECT -32.805 71.915 -32.475 72.245 ;
        RECT -32.805 70.555 -32.475 70.885 ;
        RECT -32.805 69.195 -32.475 69.525 ;
        RECT -32.805 67.835 -32.475 68.165 ;
        RECT -32.805 66.475 -32.475 66.805 ;
        RECT -32.805 65.115 -32.475 65.445 ;
        RECT -32.805 63.755 -32.475 64.085 ;
        RECT -32.805 62.395 -32.475 62.725 ;
        RECT -32.805 61.035 -32.475 61.365 ;
        RECT -32.805 59.675 -32.475 60.005 ;
        RECT -32.805 58.315 -32.475 58.645 ;
        RECT -32.805 56.955 -32.475 57.285 ;
        RECT -32.805 55.595 -32.475 55.925 ;
        RECT -32.805 54.235 -32.475 54.565 ;
        RECT -32.805 52.875 -32.475 53.205 ;
        RECT -32.805 51.515 -32.475 51.845 ;
        RECT -32.805 50.155 -32.475 50.485 ;
        RECT -32.805 48.795 -32.475 49.125 ;
        RECT -32.805 47.435 -32.475 47.765 ;
        RECT -32.805 46.075 -32.475 46.405 ;
        RECT -32.805 44.715 -32.475 45.045 ;
        RECT -32.805 43.355 -32.475 43.685 ;
        RECT -32.805 41.995 -32.475 42.325 ;
        RECT -32.805 40.635 -32.475 40.965 ;
        RECT -32.805 39.275 -32.475 39.605 ;
        RECT -32.805 37.915 -32.475 38.245 ;
        RECT -32.805 36.555 -32.475 36.885 ;
        RECT -32.805 35.195 -32.475 35.525 ;
        RECT -32.805 33.835 -32.475 34.165 ;
        RECT -32.805 32.475 -32.475 32.805 ;
        RECT -32.805 31.115 -32.475 31.445 ;
        RECT -32.805 29.755 -32.475 30.085 ;
        RECT -32.805 28.395 -32.475 28.725 ;
        RECT -32.805 27.035 -32.475 27.365 ;
        RECT -32.805 25.675 -32.475 26.005 ;
        RECT -32.805 24.315 -32.475 24.645 ;
        RECT -32.805 22.955 -32.475 23.285 ;
        RECT -32.805 21.595 -32.475 21.925 ;
        RECT -32.805 20.235 -32.475 20.565 ;
        RECT -32.805 18.875 -32.475 19.205 ;
        RECT -32.805 17.515 -32.475 17.845 ;
        RECT -32.805 16.155 -32.475 16.485 ;
        RECT -32.805 14.795 -32.475 15.125 ;
        RECT -32.805 13.435 -32.475 13.765 ;
        RECT -32.805 12.075 -32.475 12.405 ;
        RECT -32.805 10.715 -32.475 11.045 ;
        RECT -32.805 9.355 -32.475 9.685 ;
        RECT -32.805 7.995 -32.475 8.325 ;
        RECT -32.805 6.635 -32.475 6.965 ;
        RECT -32.805 5.275 -32.475 5.605 ;
        RECT -32.805 3.915 -32.475 4.245 ;
        RECT -32.805 2.555 -32.475 2.885 ;
        RECT -32.805 1.195 -32.475 1.525 ;
        RECT -32.805 -0.165 -32.475 0.165 ;
        RECT -32.805 -8.325 -32.475 -7.995 ;
        RECT -32.805 -11.045 -32.475 -10.715 ;
        RECT -32.805 -15.125 -32.475 -14.795 ;
        RECT -32.805 -16.485 -32.475 -16.155 ;
        RECT -32.805 -17.845 -32.475 -17.515 ;
        RECT -32.805 -19.205 -32.475 -18.875 ;
        RECT -32.805 -20.565 -32.475 -20.235 ;
        RECT -32.805 -21.925 -32.475 -21.595 ;
        RECT -32.805 -23.285 -32.475 -22.955 ;
        RECT -32.805 -24.645 -32.475 -24.315 ;
        RECT -32.805 -31.445 -32.475 -31.115 ;
        RECT -32.805 -32.805 -32.475 -32.475 ;
        RECT -32.805 -35.525 -32.475 -35.195 ;
        RECT -32.805 -36.885 -32.475 -36.555 ;
        RECT -32.805 -37.93 -32.475 -37.6 ;
        RECT -32.805 -40.965 -32.475 -40.635 ;
        RECT -32.805 -42.77 -32.475 -42.44 ;
        RECT -32.805 -43.685 -32.475 -43.355 ;
        RECT -32.805 -50.485 -32.475 -50.155 ;
        RECT -32.805 -51.845 -32.475 -51.515 ;
        RECT -32.805 -54.565 -32.475 -54.235 ;
        RECT -32.805 -55.925 -32.475 -55.595 ;
        RECT -32.805 -60.005 -32.475 -59.675 ;
        RECT -32.805 -68.165 -32.475 -67.835 ;
        RECT -32.805 -69.525 -32.475 -69.195 ;
        RECT -32.805 -70.885 -32.475 -70.555 ;
        RECT -32.805 -72.245 -32.475 -71.915 ;
        RECT -32.805 -73.605 -32.475 -73.275 ;
        RECT -32.805 -74.965 -32.475 -74.635 ;
        RECT -32.805 -76.325 -32.475 -75.995 ;
        RECT -32.805 -77.685 -32.475 -77.355 ;
        RECT -32.805 -79.045 -32.475 -78.715 ;
        RECT -32.805 -80.405 -32.475 -80.075 ;
        RECT -32.805 -81.765 -32.475 -81.435 ;
        RECT -32.805 -83.125 -32.475 -82.795 ;
        RECT -32.805 -84.485 -32.475 -84.155 ;
        RECT -32.805 -85.845 -32.475 -85.515 ;
        RECT -32.805 -87.205 -32.475 -86.875 ;
        RECT -32.805 -88.565 -32.475 -88.235 ;
        RECT -32.805 -89.925 -32.475 -89.595 ;
        RECT -32.805 -92.645 -32.475 -92.315 ;
        RECT -32.805 -94.005 -32.475 -93.675 ;
        RECT -32.805 -95.365 -32.475 -95.035 ;
        RECT -32.805 -96.725 -32.475 -96.395 ;
        RECT -32.805 -98.73 -32.475 -98.4 ;
        RECT -32.805 -99.445 -32.475 -99.115 ;
        RECT -32.805 -102.165 -32.475 -101.835 ;
        RECT -32.805 -103.525 -32.475 -103.195 ;
        RECT -32.805 -104.885 -32.475 -104.555 ;
        RECT -32.805 -106.87 -32.475 -106.54 ;
        RECT -32.805 -107.605 -32.475 -107.275 ;
        RECT -32.805 -108.965 -32.475 -108.635 ;
        RECT -32.805 -113.045 -32.475 -112.715 ;
        RECT -32.805 -114.405 -32.475 -114.075 ;
        RECT -32.805 -115.765 -32.475 -115.435 ;
        RECT -32.805 -117.125 -32.475 -116.795 ;
        RECT -32.805 -118.485 -32.475 -118.155 ;
        RECT -32.805 -122.565 -32.475 -122.235 ;
        RECT -32.805 -125.285 -32.475 -124.955 ;
        RECT -32.805 -126.645 -32.475 -126.315 ;
        RECT -32.805 -128.005 -32.475 -127.675 ;
        RECT -32.805 -129.365 -32.475 -129.035 ;
        RECT -32.805 -133.445 -32.475 -133.115 ;
        RECT -32.805 -134.805 -32.475 -134.475 ;
        RECT -32.805 -136.165 -32.475 -135.835 ;
        RECT -32.805 -137.525 -32.475 -137.195 ;
        RECT -32.805 -138.885 -32.475 -138.555 ;
        RECT -32.805 -141.605 -32.475 -141.275 ;
        RECT -32.805 -142.965 -32.475 -142.635 ;
        RECT -32.805 -144.325 -32.475 -143.995 ;
        RECT -32.805 -145.685 -32.475 -145.355 ;
        RECT -32.805 -147.045 -32.475 -146.715 ;
        RECT -32.805 -148.405 -32.475 -148.075 ;
        RECT -32.805 -151.125 -32.475 -150.795 ;
        RECT -32.805 -152.485 -32.475 -152.155 ;
        RECT -32.805 -156.565 -32.475 -156.235 ;
        RECT -32.805 -157.925 -32.475 -157.595 ;
        RECT -32.805 -159.285 -32.475 -158.955 ;
        RECT -32.805 -160.645 -32.475 -160.315 ;
        RECT -32.805 -162.005 -32.475 -161.675 ;
        RECT -32.805 -163.365 -32.475 -163.035 ;
        RECT -32.805 -164.725 -32.475 -164.395 ;
        RECT -32.805 -166.085 -32.475 -165.755 ;
        RECT -32.805 -167.445 -32.475 -167.115 ;
        RECT -32.805 -170.165 -32.475 -169.835 ;
        RECT -32.805 -172.885 -32.475 -172.555 ;
        RECT -32.805 -174.245 -32.475 -173.915 ;
        RECT -32.805 -175.725 -32.475 -175.395 ;
        RECT -32.805 -176.965 -32.475 -176.635 ;
        RECT -32.805 -178.325 -32.475 -177.995 ;
        RECT -32.805 -180.57 -32.475 -179.44 ;
        RECT -32.8 -180.685 -32.48 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -31.445 241.32 -31.115 242.45 ;
        RECT -31.445 239.195 -31.115 239.525 ;
        RECT -31.445 237.835 -31.115 238.165 ;
        RECT -31.445 236.475 -31.115 236.805 ;
        RECT -31.445 235.115 -31.115 235.445 ;
        RECT -31.445 233.755 -31.115 234.085 ;
        RECT -31.445 232.395 -31.115 232.725 ;
        RECT -31.445 231.035 -31.115 231.365 ;
        RECT -31.445 229.675 -31.115 230.005 ;
        RECT -31.445 228.315 -31.115 228.645 ;
        RECT -31.445 226.955 -31.115 227.285 ;
        RECT -31.445 225.595 -31.115 225.925 ;
        RECT -31.445 224.235 -31.115 224.565 ;
        RECT -31.445 222.875 -31.115 223.205 ;
        RECT -31.445 221.515 -31.115 221.845 ;
        RECT -31.445 220.155 -31.115 220.485 ;
        RECT -31.445 218.795 -31.115 219.125 ;
        RECT -31.445 217.435 -31.115 217.765 ;
        RECT -31.445 216.075 -31.115 216.405 ;
        RECT -31.445 214.715 -31.115 215.045 ;
        RECT -31.445 213.355 -31.115 213.685 ;
        RECT -31.445 211.995 -31.115 212.325 ;
        RECT -31.445 210.635 -31.115 210.965 ;
        RECT -31.445 209.275 -31.115 209.605 ;
        RECT -31.445 207.915 -31.115 208.245 ;
        RECT -31.445 206.555 -31.115 206.885 ;
        RECT -31.445 205.195 -31.115 205.525 ;
        RECT -31.445 203.835 -31.115 204.165 ;
        RECT -31.445 202.475 -31.115 202.805 ;
        RECT -31.445 201.115 -31.115 201.445 ;
        RECT -31.445 199.755 -31.115 200.085 ;
        RECT -31.445 198.395 -31.115 198.725 ;
        RECT -31.445 197.035 -31.115 197.365 ;
        RECT -31.445 195.675 -31.115 196.005 ;
        RECT -31.445 194.315 -31.115 194.645 ;
        RECT -31.445 192.955 -31.115 193.285 ;
        RECT -31.445 191.595 -31.115 191.925 ;
        RECT -31.445 190.235 -31.115 190.565 ;
        RECT -31.445 188.875 -31.115 189.205 ;
        RECT -31.445 187.515 -31.115 187.845 ;
        RECT -31.445 186.155 -31.115 186.485 ;
        RECT -31.445 184.795 -31.115 185.125 ;
        RECT -31.445 183.435 -31.115 183.765 ;
        RECT -31.445 182.075 -31.115 182.405 ;
        RECT -31.445 180.715 -31.115 181.045 ;
        RECT -31.445 179.355 -31.115 179.685 ;
        RECT -31.445 177.995 -31.115 178.325 ;
        RECT -31.445 176.635 -31.115 176.965 ;
        RECT -31.445 175.275 -31.115 175.605 ;
        RECT -31.445 173.915 -31.115 174.245 ;
        RECT -31.445 172.555 -31.115 172.885 ;
        RECT -31.445 171.195 -31.115 171.525 ;
        RECT -31.445 169.835 -31.115 170.165 ;
        RECT -31.445 168.475 -31.115 168.805 ;
        RECT -31.445 167.115 -31.115 167.445 ;
        RECT -31.445 165.755 -31.115 166.085 ;
        RECT -31.445 164.395 -31.115 164.725 ;
        RECT -31.445 163.035 -31.115 163.365 ;
        RECT -31.445 161.675 -31.115 162.005 ;
        RECT -31.445 160.315 -31.115 160.645 ;
        RECT -31.445 158.955 -31.115 159.285 ;
        RECT -31.445 157.595 -31.115 157.925 ;
        RECT -31.445 156.235 -31.115 156.565 ;
        RECT -31.445 154.875 -31.115 155.205 ;
        RECT -31.445 153.515 -31.115 153.845 ;
        RECT -31.445 152.155 -31.115 152.485 ;
        RECT -31.445 150.795 -31.115 151.125 ;
        RECT -31.445 149.435 -31.115 149.765 ;
        RECT -31.445 148.075 -31.115 148.405 ;
        RECT -31.445 146.715 -31.115 147.045 ;
        RECT -31.445 145.355 -31.115 145.685 ;
        RECT -31.445 143.995 -31.115 144.325 ;
        RECT -31.445 142.635 -31.115 142.965 ;
        RECT -31.445 141.275 -31.115 141.605 ;
        RECT -31.445 139.915 -31.115 140.245 ;
        RECT -31.445 138.555 -31.115 138.885 ;
        RECT -31.445 137.195 -31.115 137.525 ;
        RECT -31.445 135.835 -31.115 136.165 ;
        RECT -31.445 134.475 -31.115 134.805 ;
        RECT -31.445 133.115 -31.115 133.445 ;
        RECT -31.445 131.755 -31.115 132.085 ;
        RECT -31.445 130.395 -31.115 130.725 ;
        RECT -31.445 129.035 -31.115 129.365 ;
        RECT -31.445 127.675 -31.115 128.005 ;
        RECT -31.445 126.315 -31.115 126.645 ;
        RECT -31.445 124.955 -31.115 125.285 ;
        RECT -31.445 123.595 -31.115 123.925 ;
        RECT -31.445 122.235 -31.115 122.565 ;
        RECT -31.445 120.875 -31.115 121.205 ;
        RECT -31.445 119.515 -31.115 119.845 ;
        RECT -31.445 118.155 -31.115 118.485 ;
        RECT -31.445 116.795 -31.115 117.125 ;
        RECT -31.445 115.435 -31.115 115.765 ;
        RECT -31.445 114.075 -31.115 114.405 ;
        RECT -31.445 112.715 -31.115 113.045 ;
        RECT -31.445 111.355 -31.115 111.685 ;
        RECT -31.445 109.995 -31.115 110.325 ;
        RECT -31.445 108.635 -31.115 108.965 ;
        RECT -31.445 107.275 -31.115 107.605 ;
        RECT -31.445 105.915 -31.115 106.245 ;
        RECT -31.445 104.555 -31.115 104.885 ;
        RECT -31.445 103.195 -31.115 103.525 ;
        RECT -31.445 101.835 -31.115 102.165 ;
        RECT -31.445 100.475 -31.115 100.805 ;
        RECT -31.445 99.115 -31.115 99.445 ;
        RECT -31.445 97.755 -31.115 98.085 ;
        RECT -31.445 96.395 -31.115 96.725 ;
        RECT -31.445 95.035 -31.115 95.365 ;
        RECT -31.445 93.675 -31.115 94.005 ;
        RECT -31.445 92.315 -31.115 92.645 ;
        RECT -31.445 90.955 -31.115 91.285 ;
        RECT -31.445 89.595 -31.115 89.925 ;
        RECT -31.445 88.235 -31.115 88.565 ;
        RECT -31.445 86.875 -31.115 87.205 ;
        RECT -31.445 85.515 -31.115 85.845 ;
        RECT -31.445 84.155 -31.115 84.485 ;
        RECT -31.445 82.795 -31.115 83.125 ;
        RECT -31.445 81.435 -31.115 81.765 ;
        RECT -31.445 80.075 -31.115 80.405 ;
        RECT -31.445 78.715 -31.115 79.045 ;
        RECT -31.445 77.355 -31.115 77.685 ;
        RECT -31.445 75.995 -31.115 76.325 ;
        RECT -31.445 74.635 -31.115 74.965 ;
        RECT -31.445 73.275 -31.115 73.605 ;
        RECT -31.445 71.915 -31.115 72.245 ;
        RECT -31.445 70.555 -31.115 70.885 ;
        RECT -31.445 69.195 -31.115 69.525 ;
        RECT -31.445 67.835 -31.115 68.165 ;
        RECT -31.445 66.475 -31.115 66.805 ;
        RECT -31.445 65.115 -31.115 65.445 ;
        RECT -31.445 63.755 -31.115 64.085 ;
        RECT -31.445 62.395 -31.115 62.725 ;
        RECT -31.445 61.035 -31.115 61.365 ;
        RECT -31.445 59.675 -31.115 60.005 ;
        RECT -31.445 58.315 -31.115 58.645 ;
        RECT -31.445 56.955 -31.115 57.285 ;
        RECT -31.445 55.595 -31.115 55.925 ;
        RECT -31.445 54.235 -31.115 54.565 ;
        RECT -31.445 52.875 -31.115 53.205 ;
        RECT -31.445 51.515 -31.115 51.845 ;
        RECT -31.445 50.155 -31.115 50.485 ;
        RECT -31.445 48.795 -31.115 49.125 ;
        RECT -31.445 47.435 -31.115 47.765 ;
        RECT -31.445 46.075 -31.115 46.405 ;
        RECT -31.445 44.715 -31.115 45.045 ;
        RECT -31.445 43.355 -31.115 43.685 ;
        RECT -31.445 41.995 -31.115 42.325 ;
        RECT -31.445 40.635 -31.115 40.965 ;
        RECT -31.445 39.275 -31.115 39.605 ;
        RECT -31.445 37.915 -31.115 38.245 ;
        RECT -31.445 36.555 -31.115 36.885 ;
        RECT -31.445 35.195 -31.115 35.525 ;
        RECT -31.445 33.835 -31.115 34.165 ;
        RECT -31.445 32.475 -31.115 32.805 ;
        RECT -31.445 31.115 -31.115 31.445 ;
        RECT -31.445 29.755 -31.115 30.085 ;
        RECT -31.445 28.395 -31.115 28.725 ;
        RECT -31.445 27.035 -31.115 27.365 ;
        RECT -31.445 25.675 -31.115 26.005 ;
        RECT -31.445 24.315 -31.115 24.645 ;
        RECT -31.445 22.955 -31.115 23.285 ;
        RECT -31.445 21.595 -31.115 21.925 ;
        RECT -31.445 20.235 -31.115 20.565 ;
        RECT -31.445 18.875 -31.115 19.205 ;
        RECT -31.445 17.515 -31.115 17.845 ;
        RECT -31.445 16.155 -31.115 16.485 ;
        RECT -31.445 14.795 -31.115 15.125 ;
        RECT -31.445 13.435 -31.115 13.765 ;
        RECT -31.445 12.075 -31.115 12.405 ;
        RECT -31.445 10.715 -31.115 11.045 ;
        RECT -31.445 9.355 -31.115 9.685 ;
        RECT -31.445 7.995 -31.115 8.325 ;
        RECT -31.445 6.635 -31.115 6.965 ;
        RECT -31.445 5.275 -31.115 5.605 ;
        RECT -31.445 3.915 -31.115 4.245 ;
        RECT -31.445 2.555 -31.115 2.885 ;
        RECT -31.445 1.195 -31.115 1.525 ;
        RECT -31.445 -0.165 -31.115 0.165 ;
        RECT -31.445 -8.325 -31.115 -7.995 ;
        RECT -31.445 -11.045 -31.115 -10.715 ;
        RECT -31.445 -15.125 -31.115 -14.795 ;
        RECT -31.445 -16.485 -31.115 -16.155 ;
        RECT -31.445 -17.845 -31.115 -17.515 ;
        RECT -31.445 -19.205 -31.115 -18.875 ;
        RECT -31.445 -20.565 -31.115 -20.235 ;
        RECT -31.445 -21.925 -31.115 -21.595 ;
        RECT -31.445 -23.285 -31.115 -22.955 ;
        RECT -31.445 -24.645 -31.115 -24.315 ;
        RECT -31.445 -31.445 -31.115 -31.115 ;
        RECT -31.445 -32.805 -31.115 -32.475 ;
        RECT -31.445 -35.525 -31.115 -35.195 ;
        RECT -31.445 -36.885 -31.115 -36.555 ;
        RECT -31.445 -37.93 -31.115 -37.6 ;
        RECT -31.445 -40.965 -31.115 -40.635 ;
        RECT -31.445 -42.77 -31.115 -42.44 ;
        RECT -31.445 -43.685 -31.115 -43.355 ;
        RECT -31.445 -50.485 -31.115 -50.155 ;
        RECT -31.445 -51.845 -31.115 -51.515 ;
        RECT -31.445 -54.565 -31.115 -54.235 ;
        RECT -31.445 -55.925 -31.115 -55.595 ;
        RECT -31.445 -60.005 -31.115 -59.675 ;
        RECT -31.445 -68.165 -31.115 -67.835 ;
        RECT -31.445 -69.525 -31.115 -69.195 ;
        RECT -31.445 -70.885 -31.115 -70.555 ;
        RECT -31.445 -72.245 -31.115 -71.915 ;
        RECT -31.445 -73.605 -31.115 -73.275 ;
        RECT -31.445 -74.965 -31.115 -74.635 ;
        RECT -31.445 -76.325 -31.115 -75.995 ;
        RECT -31.445 -77.685 -31.115 -77.355 ;
        RECT -31.445 -79.045 -31.115 -78.715 ;
        RECT -31.445 -80.405 -31.115 -80.075 ;
        RECT -31.445 -81.765 -31.115 -81.435 ;
        RECT -31.445 -83.125 -31.115 -82.795 ;
        RECT -31.445 -84.485 -31.115 -84.155 ;
        RECT -31.445 -85.845 -31.115 -85.515 ;
        RECT -31.445 -87.205 -31.115 -86.875 ;
        RECT -31.445 -88.565 -31.115 -88.235 ;
        RECT -31.445 -89.925 -31.115 -89.595 ;
        RECT -31.445 -92.645 -31.115 -92.315 ;
        RECT -31.445 -94.005 -31.115 -93.675 ;
        RECT -31.445 -95.365 -31.115 -95.035 ;
        RECT -31.445 -96.725 -31.115 -96.395 ;
        RECT -31.445 -98.73 -31.115 -98.4 ;
        RECT -31.445 -99.445 -31.115 -99.115 ;
        RECT -31.445 -102.165 -31.115 -101.835 ;
        RECT -31.445 -103.525 -31.115 -103.195 ;
        RECT -31.445 -104.885 -31.115 -104.555 ;
        RECT -31.445 -106.87 -31.115 -106.54 ;
        RECT -31.445 -107.605 -31.115 -107.275 ;
        RECT -31.445 -108.965 -31.115 -108.635 ;
        RECT -31.445 -113.045 -31.115 -112.715 ;
        RECT -31.445 -114.405 -31.115 -114.075 ;
        RECT -31.445 -115.765 -31.115 -115.435 ;
        RECT -31.445 -117.125 -31.115 -116.795 ;
        RECT -31.445 -118.485 -31.115 -118.155 ;
        RECT -31.445 -122.565 -31.115 -122.235 ;
        RECT -31.445 -123.925 -31.115 -123.595 ;
        RECT -31.445 -125.285 -31.115 -124.955 ;
        RECT -31.445 -126.645 -31.115 -126.315 ;
        RECT -31.445 -128.005 -31.115 -127.675 ;
        RECT -31.445 -129.365 -31.115 -129.035 ;
        RECT -31.445 -133.445 -31.115 -133.115 ;
        RECT -31.445 -134.805 -31.115 -134.475 ;
        RECT -31.445 -136.165 -31.115 -135.835 ;
        RECT -31.445 -138.885 -31.115 -138.555 ;
        RECT -31.445 -141.605 -31.115 -141.275 ;
        RECT -31.445 -142.965 -31.115 -142.635 ;
        RECT -31.445 -144.325 -31.115 -143.995 ;
        RECT -31.445 -145.685 -31.115 -145.355 ;
        RECT -31.445 -147.045 -31.115 -146.715 ;
        RECT -31.445 -148.405 -31.115 -148.075 ;
        RECT -31.445 -151.125 -31.115 -150.795 ;
        RECT -31.445 -152.485 -31.115 -152.155 ;
        RECT -31.445 -156.565 -31.115 -156.235 ;
        RECT -31.445 -157.925 -31.115 -157.595 ;
        RECT -31.445 -159.285 -31.115 -158.955 ;
        RECT -31.445 -160.645 -31.115 -160.315 ;
        RECT -31.445 -162.005 -31.115 -161.675 ;
        RECT -31.445 -163.365 -31.115 -163.035 ;
        RECT -31.445 -164.725 -31.115 -164.395 ;
        RECT -31.445 -166.085 -31.115 -165.755 ;
        RECT -31.445 -167.445 -31.115 -167.115 ;
        RECT -31.445 -170.165 -31.115 -169.835 ;
        RECT -31.445 -172.885 -31.115 -172.555 ;
        RECT -31.445 -174.245 -31.115 -173.915 ;
        RECT -31.445 -175.725 -31.115 -175.395 ;
        RECT -31.445 -176.965 -31.115 -176.635 ;
        RECT -31.445 -178.325 -31.115 -177.995 ;
        RECT -31.445 -180.57 -31.115 -179.44 ;
        RECT -31.44 -180.685 -31.12 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -30.085 241.32 -29.755 242.45 ;
        RECT -30.085 239.195 -29.755 239.525 ;
        RECT -30.085 237.835 -29.755 238.165 ;
        RECT -30.085 236.475 -29.755 236.805 ;
        RECT -30.085 235.115 -29.755 235.445 ;
        RECT -30.085 233.755 -29.755 234.085 ;
        RECT -30.085 232.395 -29.755 232.725 ;
        RECT -30.085 231.035 -29.755 231.365 ;
        RECT -30.085 229.675 -29.755 230.005 ;
        RECT -30.085 228.315 -29.755 228.645 ;
        RECT -30.085 226.955 -29.755 227.285 ;
        RECT -30.085 225.595 -29.755 225.925 ;
        RECT -30.085 224.235 -29.755 224.565 ;
        RECT -30.085 222.875 -29.755 223.205 ;
        RECT -30.085 221.515 -29.755 221.845 ;
        RECT -30.085 220.155 -29.755 220.485 ;
        RECT -30.085 218.795 -29.755 219.125 ;
        RECT -30.085 217.435 -29.755 217.765 ;
        RECT -30.085 216.075 -29.755 216.405 ;
        RECT -30.085 214.715 -29.755 215.045 ;
        RECT -30.085 213.355 -29.755 213.685 ;
        RECT -30.085 211.995 -29.755 212.325 ;
        RECT -30.085 210.635 -29.755 210.965 ;
        RECT -30.085 209.275 -29.755 209.605 ;
        RECT -30.085 207.915 -29.755 208.245 ;
        RECT -30.085 206.555 -29.755 206.885 ;
        RECT -30.085 205.195 -29.755 205.525 ;
        RECT -30.085 203.835 -29.755 204.165 ;
        RECT -30.085 202.475 -29.755 202.805 ;
        RECT -30.085 201.115 -29.755 201.445 ;
        RECT -30.085 199.755 -29.755 200.085 ;
        RECT -30.085 198.395 -29.755 198.725 ;
        RECT -30.085 197.035 -29.755 197.365 ;
        RECT -30.085 195.675 -29.755 196.005 ;
        RECT -30.085 194.315 -29.755 194.645 ;
        RECT -30.085 192.955 -29.755 193.285 ;
        RECT -30.085 191.595 -29.755 191.925 ;
        RECT -30.085 190.235 -29.755 190.565 ;
        RECT -30.085 188.875 -29.755 189.205 ;
        RECT -30.085 187.515 -29.755 187.845 ;
        RECT -30.085 186.155 -29.755 186.485 ;
        RECT -30.085 184.795 -29.755 185.125 ;
        RECT -30.085 183.435 -29.755 183.765 ;
        RECT -30.085 182.075 -29.755 182.405 ;
        RECT -30.085 180.715 -29.755 181.045 ;
        RECT -30.085 179.355 -29.755 179.685 ;
        RECT -30.085 177.995 -29.755 178.325 ;
        RECT -30.085 176.635 -29.755 176.965 ;
        RECT -30.085 175.275 -29.755 175.605 ;
        RECT -30.085 173.915 -29.755 174.245 ;
        RECT -30.085 172.555 -29.755 172.885 ;
        RECT -30.085 171.195 -29.755 171.525 ;
        RECT -30.085 169.835 -29.755 170.165 ;
        RECT -30.085 168.475 -29.755 168.805 ;
        RECT -30.085 167.115 -29.755 167.445 ;
        RECT -30.085 165.755 -29.755 166.085 ;
        RECT -30.085 164.395 -29.755 164.725 ;
        RECT -30.085 163.035 -29.755 163.365 ;
        RECT -30.085 161.675 -29.755 162.005 ;
        RECT -30.085 160.315 -29.755 160.645 ;
        RECT -30.085 158.955 -29.755 159.285 ;
        RECT -30.085 157.595 -29.755 157.925 ;
        RECT -30.085 156.235 -29.755 156.565 ;
        RECT -30.085 154.875 -29.755 155.205 ;
        RECT -30.085 153.515 -29.755 153.845 ;
        RECT -30.085 152.155 -29.755 152.485 ;
        RECT -30.085 150.795 -29.755 151.125 ;
        RECT -30.085 149.435 -29.755 149.765 ;
        RECT -30.085 148.075 -29.755 148.405 ;
        RECT -30.085 146.715 -29.755 147.045 ;
        RECT -30.085 145.355 -29.755 145.685 ;
        RECT -30.085 143.995 -29.755 144.325 ;
        RECT -30.085 142.635 -29.755 142.965 ;
        RECT -30.085 141.275 -29.755 141.605 ;
        RECT -30.085 139.915 -29.755 140.245 ;
        RECT -30.085 138.555 -29.755 138.885 ;
        RECT -30.085 137.195 -29.755 137.525 ;
        RECT -30.085 135.835 -29.755 136.165 ;
        RECT -30.085 134.475 -29.755 134.805 ;
        RECT -30.085 133.115 -29.755 133.445 ;
        RECT -30.085 131.755 -29.755 132.085 ;
        RECT -30.085 130.395 -29.755 130.725 ;
        RECT -30.085 129.035 -29.755 129.365 ;
        RECT -30.085 127.675 -29.755 128.005 ;
        RECT -30.085 126.315 -29.755 126.645 ;
        RECT -30.085 124.955 -29.755 125.285 ;
        RECT -30.085 123.595 -29.755 123.925 ;
        RECT -30.085 122.235 -29.755 122.565 ;
        RECT -30.085 120.875 -29.755 121.205 ;
        RECT -30.085 119.515 -29.755 119.845 ;
        RECT -30.085 118.155 -29.755 118.485 ;
        RECT -30.085 116.795 -29.755 117.125 ;
        RECT -30.085 115.435 -29.755 115.765 ;
        RECT -30.085 114.075 -29.755 114.405 ;
        RECT -30.085 112.715 -29.755 113.045 ;
        RECT -30.085 111.355 -29.755 111.685 ;
        RECT -30.085 109.995 -29.755 110.325 ;
        RECT -30.085 108.635 -29.755 108.965 ;
        RECT -30.085 107.275 -29.755 107.605 ;
        RECT -30.085 105.915 -29.755 106.245 ;
        RECT -30.085 104.555 -29.755 104.885 ;
        RECT -30.085 103.195 -29.755 103.525 ;
        RECT -30.085 101.835 -29.755 102.165 ;
        RECT -30.085 100.475 -29.755 100.805 ;
        RECT -30.085 99.115 -29.755 99.445 ;
        RECT -30.085 97.755 -29.755 98.085 ;
        RECT -30.085 96.395 -29.755 96.725 ;
        RECT -30.085 95.035 -29.755 95.365 ;
        RECT -30.085 93.675 -29.755 94.005 ;
        RECT -30.085 92.315 -29.755 92.645 ;
        RECT -30.085 90.955 -29.755 91.285 ;
        RECT -30.085 89.595 -29.755 89.925 ;
        RECT -30.085 88.235 -29.755 88.565 ;
        RECT -30.085 86.875 -29.755 87.205 ;
        RECT -30.085 85.515 -29.755 85.845 ;
        RECT -30.085 84.155 -29.755 84.485 ;
        RECT -30.085 82.795 -29.755 83.125 ;
        RECT -30.085 81.435 -29.755 81.765 ;
        RECT -30.085 80.075 -29.755 80.405 ;
        RECT -30.085 78.715 -29.755 79.045 ;
        RECT -30.085 77.355 -29.755 77.685 ;
        RECT -30.085 75.995 -29.755 76.325 ;
        RECT -30.085 74.635 -29.755 74.965 ;
        RECT -30.085 73.275 -29.755 73.605 ;
        RECT -30.085 71.915 -29.755 72.245 ;
        RECT -30.085 70.555 -29.755 70.885 ;
        RECT -30.085 69.195 -29.755 69.525 ;
        RECT -30.085 67.835 -29.755 68.165 ;
        RECT -30.085 66.475 -29.755 66.805 ;
        RECT -30.085 65.115 -29.755 65.445 ;
        RECT -30.085 63.755 -29.755 64.085 ;
        RECT -30.085 62.395 -29.755 62.725 ;
        RECT -30.085 61.035 -29.755 61.365 ;
        RECT -30.085 59.675 -29.755 60.005 ;
        RECT -30.085 58.315 -29.755 58.645 ;
        RECT -30.085 56.955 -29.755 57.285 ;
        RECT -30.085 55.595 -29.755 55.925 ;
        RECT -30.085 54.235 -29.755 54.565 ;
        RECT -30.085 52.875 -29.755 53.205 ;
        RECT -30.085 51.515 -29.755 51.845 ;
        RECT -30.085 50.155 -29.755 50.485 ;
        RECT -30.085 48.795 -29.755 49.125 ;
        RECT -30.085 47.435 -29.755 47.765 ;
        RECT -30.085 46.075 -29.755 46.405 ;
        RECT -30.085 44.715 -29.755 45.045 ;
        RECT -30.085 43.355 -29.755 43.685 ;
        RECT -30.085 41.995 -29.755 42.325 ;
        RECT -30.085 40.635 -29.755 40.965 ;
        RECT -30.085 39.275 -29.755 39.605 ;
        RECT -30.085 37.915 -29.755 38.245 ;
        RECT -30.085 36.555 -29.755 36.885 ;
        RECT -30.085 35.195 -29.755 35.525 ;
        RECT -30.085 33.835 -29.755 34.165 ;
        RECT -30.085 32.475 -29.755 32.805 ;
        RECT -30.085 31.115 -29.755 31.445 ;
        RECT -30.085 29.755 -29.755 30.085 ;
        RECT -30.085 28.395 -29.755 28.725 ;
        RECT -30.085 27.035 -29.755 27.365 ;
        RECT -30.085 25.675 -29.755 26.005 ;
        RECT -30.085 24.315 -29.755 24.645 ;
        RECT -30.085 22.955 -29.755 23.285 ;
        RECT -30.085 21.595 -29.755 21.925 ;
        RECT -30.085 20.235 -29.755 20.565 ;
        RECT -30.085 18.875 -29.755 19.205 ;
        RECT -30.085 17.515 -29.755 17.845 ;
        RECT -30.085 16.155 -29.755 16.485 ;
        RECT -30.085 14.795 -29.755 15.125 ;
        RECT -30.085 13.435 -29.755 13.765 ;
        RECT -30.085 12.075 -29.755 12.405 ;
        RECT -30.085 10.715 -29.755 11.045 ;
        RECT -30.085 9.355 -29.755 9.685 ;
        RECT -30.085 7.995 -29.755 8.325 ;
        RECT -30.085 6.635 -29.755 6.965 ;
        RECT -30.085 5.275 -29.755 5.605 ;
        RECT -30.085 3.915 -29.755 4.245 ;
        RECT -30.085 2.555 -29.755 2.885 ;
        RECT -30.085 1.195 -29.755 1.525 ;
        RECT -30.085 -0.165 -29.755 0.165 ;
        RECT -30.085 -8.325 -29.755 -7.995 ;
        RECT -30.085 -9.685 -29.755 -9.355 ;
        RECT -30.085 -17.845 -29.755 -17.515 ;
        RECT -30.085 -20.565 -29.755 -20.235 ;
        RECT -30.085 -31.445 -29.755 -31.115 ;
        RECT -30.085 -32.805 -29.755 -32.475 ;
        RECT -30.085 -35.525 -29.755 -35.195 ;
        RECT -30.085 -36.885 -29.755 -36.555 ;
        RECT -30.085 -37.93 -29.755 -37.6 ;
        RECT -30.085 -40.965 -29.755 -40.635 ;
        RECT -30.085 -42.77 -29.755 -42.44 ;
        RECT -30.085 -43.685 -29.755 -43.355 ;
        RECT -30.085 -50.485 -29.755 -50.155 ;
        RECT -30.085 -51.845 -29.755 -51.515 ;
        RECT -30.085 -54.565 -29.755 -54.235 ;
        RECT -30.085 -55.925 -29.755 -55.595 ;
        RECT -30.085 -60.005 -29.755 -59.675 ;
        RECT -30.08 -64.08 -29.76 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -30.085 -69.525 -29.755 -69.195 ;
        RECT -30.085 -70.885 -29.755 -70.555 ;
        RECT -30.085 -72.245 -29.755 -71.915 ;
        RECT -30.085 -73.605 -29.755 -73.275 ;
        RECT -30.085 -74.965 -29.755 -74.635 ;
        RECT -30.085 -76.325 -29.755 -75.995 ;
        RECT -30.085 -77.685 -29.755 -77.355 ;
        RECT -30.085 -79.045 -29.755 -78.715 ;
        RECT -30.085 -80.405 -29.755 -80.075 ;
        RECT -30.085 -81.765 -29.755 -81.435 ;
        RECT -30.085 -83.125 -29.755 -82.795 ;
        RECT -30.085 -84.485 -29.755 -84.155 ;
        RECT -30.085 -85.845 -29.755 -85.515 ;
        RECT -30.085 -87.205 -29.755 -86.875 ;
        RECT -30.085 -88.565 -29.755 -88.235 ;
        RECT -30.085 -89.925 -29.755 -89.595 ;
        RECT -30.085 -92.645 -29.755 -92.315 ;
        RECT -30.085 -94.005 -29.755 -93.675 ;
        RECT -30.085 -95.365 -29.755 -95.035 ;
        RECT -30.085 -96.725 -29.755 -96.395 ;
        RECT -30.085 -98.73 -29.755 -98.4 ;
        RECT -30.085 -99.445 -29.755 -99.115 ;
        RECT -30.085 -102.165 -29.755 -101.835 ;
        RECT -30.085 -103.525 -29.755 -103.195 ;
        RECT -30.085 -104.885 -29.755 -104.555 ;
        RECT -30.085 -106.87 -29.755 -106.54 ;
        RECT -30.085 -107.605 -29.755 -107.275 ;
        RECT -30.085 -108.965 -29.755 -108.635 ;
        RECT -30.08 -111.68 -29.76 -68.52 ;
    END
    PORT
      LAYER met3 ;
        RECT -30.085 -174.245 -29.755 -173.915 ;
        RECT -30.085 -175.725 -29.755 -175.395 ;
        RECT -30.085 -176.965 -29.755 -176.635 ;
        RECT -30.085 -178.325 -29.755 -177.995 ;
        RECT -30.085 -180.57 -29.755 -179.44 ;
        RECT -30.08 -180.685 -29.76 -172.56 ;
    END
    PORT
      LAYER met3 ;
        RECT -28.725 -0.165 -28.395 0.165 ;
        RECT -28.725 -8.325 -28.395 -7.995 ;
        RECT -28.725 -9.685 -28.395 -9.355 ;
        RECT -28.725 -14.95 -28.395 -14.62 ;
        RECT -28.725 -17.845 -28.395 -17.515 ;
        RECT -28.725 -19.79 -28.395 -19.46 ;
        RECT -28.725 -20.565 -28.395 -20.235 ;
        RECT -28.725 -31.445 -28.395 -31.115 ;
        RECT -28.725 -32.805 -28.395 -32.475 ;
        RECT -28.725 -35.525 -28.395 -35.195 ;
        RECT -28.725 -36.885 -28.395 -36.555 ;
        RECT -28.725 -37.93 -28.395 -37.6 ;
        RECT -28.725 -40.965 -28.395 -40.635 ;
        RECT -28.725 -42.77 -28.395 -42.44 ;
        RECT -28.725 -43.685 -28.395 -43.355 ;
        RECT -28.725 -50.485 -28.395 -50.155 ;
        RECT -28.725 -51.845 -28.395 -51.515 ;
        RECT -28.725 -54.565 -28.395 -54.235 ;
        RECT -28.725 -55.925 -28.395 -55.595 ;
        RECT -28.725 -60.005 -28.395 -59.675 ;
        RECT -28.72 -63.4 -28.4 242.565 ;
        RECT -28.725 241.32 -28.395 242.45 ;
        RECT -28.725 239.195 -28.395 239.525 ;
        RECT -28.725 237.835 -28.395 238.165 ;
        RECT -28.725 236.475 -28.395 236.805 ;
        RECT -28.725 235.115 -28.395 235.445 ;
        RECT -28.725 233.755 -28.395 234.085 ;
        RECT -28.725 232.395 -28.395 232.725 ;
        RECT -28.725 231.035 -28.395 231.365 ;
        RECT -28.725 229.675 -28.395 230.005 ;
        RECT -28.725 228.315 -28.395 228.645 ;
        RECT -28.725 226.955 -28.395 227.285 ;
        RECT -28.725 225.595 -28.395 225.925 ;
        RECT -28.725 224.235 -28.395 224.565 ;
        RECT -28.725 222.875 -28.395 223.205 ;
        RECT -28.725 221.515 -28.395 221.845 ;
        RECT -28.725 220.155 -28.395 220.485 ;
        RECT -28.725 218.795 -28.395 219.125 ;
        RECT -28.725 217.435 -28.395 217.765 ;
        RECT -28.725 216.075 -28.395 216.405 ;
        RECT -28.725 214.715 -28.395 215.045 ;
        RECT -28.725 213.355 -28.395 213.685 ;
        RECT -28.725 211.995 -28.395 212.325 ;
        RECT -28.725 210.635 -28.395 210.965 ;
        RECT -28.725 209.275 -28.395 209.605 ;
        RECT -28.725 207.915 -28.395 208.245 ;
        RECT -28.725 206.555 -28.395 206.885 ;
        RECT -28.725 205.195 -28.395 205.525 ;
        RECT -28.725 203.835 -28.395 204.165 ;
        RECT -28.725 202.475 -28.395 202.805 ;
        RECT -28.725 201.115 -28.395 201.445 ;
        RECT -28.725 199.755 -28.395 200.085 ;
        RECT -28.725 198.395 -28.395 198.725 ;
        RECT -28.725 197.035 -28.395 197.365 ;
        RECT -28.725 195.675 -28.395 196.005 ;
        RECT -28.725 194.315 -28.395 194.645 ;
        RECT -28.725 192.955 -28.395 193.285 ;
        RECT -28.725 191.595 -28.395 191.925 ;
        RECT -28.725 190.235 -28.395 190.565 ;
        RECT -28.725 188.875 -28.395 189.205 ;
        RECT -28.725 187.515 -28.395 187.845 ;
        RECT -28.725 186.155 -28.395 186.485 ;
        RECT -28.725 184.795 -28.395 185.125 ;
        RECT -28.725 183.435 -28.395 183.765 ;
        RECT -28.725 182.075 -28.395 182.405 ;
        RECT -28.725 180.715 -28.395 181.045 ;
        RECT -28.725 179.355 -28.395 179.685 ;
        RECT -28.725 177.995 -28.395 178.325 ;
        RECT -28.725 176.635 -28.395 176.965 ;
        RECT -28.725 175.275 -28.395 175.605 ;
        RECT -28.725 173.915 -28.395 174.245 ;
        RECT -28.725 172.555 -28.395 172.885 ;
        RECT -28.725 171.195 -28.395 171.525 ;
        RECT -28.725 169.835 -28.395 170.165 ;
        RECT -28.725 168.475 -28.395 168.805 ;
        RECT -28.725 167.115 -28.395 167.445 ;
        RECT -28.725 165.755 -28.395 166.085 ;
        RECT -28.725 164.395 -28.395 164.725 ;
        RECT -28.725 163.035 -28.395 163.365 ;
        RECT -28.725 161.675 -28.395 162.005 ;
        RECT -28.725 160.315 -28.395 160.645 ;
        RECT -28.725 158.955 -28.395 159.285 ;
        RECT -28.725 157.595 -28.395 157.925 ;
        RECT -28.725 156.235 -28.395 156.565 ;
        RECT -28.725 154.875 -28.395 155.205 ;
        RECT -28.725 153.515 -28.395 153.845 ;
        RECT -28.725 152.155 -28.395 152.485 ;
        RECT -28.725 150.795 -28.395 151.125 ;
        RECT -28.725 149.435 -28.395 149.765 ;
        RECT -28.725 148.075 -28.395 148.405 ;
        RECT -28.725 146.715 -28.395 147.045 ;
        RECT -28.725 145.355 -28.395 145.685 ;
        RECT -28.725 143.995 -28.395 144.325 ;
        RECT -28.725 142.635 -28.395 142.965 ;
        RECT -28.725 141.275 -28.395 141.605 ;
        RECT -28.725 139.915 -28.395 140.245 ;
        RECT -28.725 138.555 -28.395 138.885 ;
        RECT -28.725 137.195 -28.395 137.525 ;
        RECT -28.725 135.835 -28.395 136.165 ;
        RECT -28.725 134.475 -28.395 134.805 ;
        RECT -28.725 133.115 -28.395 133.445 ;
        RECT -28.725 131.755 -28.395 132.085 ;
        RECT -28.725 130.395 -28.395 130.725 ;
        RECT -28.725 129.035 -28.395 129.365 ;
        RECT -28.725 127.675 -28.395 128.005 ;
        RECT -28.725 126.315 -28.395 126.645 ;
        RECT -28.725 124.955 -28.395 125.285 ;
        RECT -28.725 123.595 -28.395 123.925 ;
        RECT -28.725 122.235 -28.395 122.565 ;
        RECT -28.725 120.875 -28.395 121.205 ;
        RECT -28.725 119.515 -28.395 119.845 ;
        RECT -28.725 118.155 -28.395 118.485 ;
        RECT -28.725 116.795 -28.395 117.125 ;
        RECT -28.725 115.435 -28.395 115.765 ;
        RECT -28.725 114.075 -28.395 114.405 ;
        RECT -28.725 112.715 -28.395 113.045 ;
        RECT -28.725 111.355 -28.395 111.685 ;
        RECT -28.725 109.995 -28.395 110.325 ;
        RECT -28.725 108.635 -28.395 108.965 ;
        RECT -28.725 107.275 -28.395 107.605 ;
        RECT -28.725 105.915 -28.395 106.245 ;
        RECT -28.725 104.555 -28.395 104.885 ;
        RECT -28.725 103.195 -28.395 103.525 ;
        RECT -28.725 101.835 -28.395 102.165 ;
        RECT -28.725 100.475 -28.395 100.805 ;
        RECT -28.725 99.115 -28.395 99.445 ;
        RECT -28.725 97.755 -28.395 98.085 ;
        RECT -28.725 96.395 -28.395 96.725 ;
        RECT -28.725 95.035 -28.395 95.365 ;
        RECT -28.725 93.675 -28.395 94.005 ;
        RECT -28.725 92.315 -28.395 92.645 ;
        RECT -28.725 90.955 -28.395 91.285 ;
        RECT -28.725 89.595 -28.395 89.925 ;
        RECT -28.725 88.235 -28.395 88.565 ;
        RECT -28.725 86.875 -28.395 87.205 ;
        RECT -28.725 85.515 -28.395 85.845 ;
        RECT -28.725 84.155 -28.395 84.485 ;
        RECT -28.725 82.795 -28.395 83.125 ;
        RECT -28.725 81.435 -28.395 81.765 ;
        RECT -28.725 80.075 -28.395 80.405 ;
        RECT -28.725 78.715 -28.395 79.045 ;
        RECT -28.725 77.355 -28.395 77.685 ;
        RECT -28.725 75.995 -28.395 76.325 ;
        RECT -28.725 74.635 -28.395 74.965 ;
        RECT -28.725 73.275 -28.395 73.605 ;
        RECT -28.725 71.915 -28.395 72.245 ;
        RECT -28.725 70.555 -28.395 70.885 ;
        RECT -28.725 69.195 -28.395 69.525 ;
        RECT -28.725 67.835 -28.395 68.165 ;
        RECT -28.725 66.475 -28.395 66.805 ;
        RECT -28.725 65.115 -28.395 65.445 ;
        RECT -28.725 63.755 -28.395 64.085 ;
        RECT -28.725 62.395 -28.395 62.725 ;
        RECT -28.725 61.035 -28.395 61.365 ;
        RECT -28.725 59.675 -28.395 60.005 ;
        RECT -28.725 58.315 -28.395 58.645 ;
        RECT -28.725 56.955 -28.395 57.285 ;
        RECT -28.725 55.595 -28.395 55.925 ;
        RECT -28.725 54.235 -28.395 54.565 ;
        RECT -28.725 52.875 -28.395 53.205 ;
        RECT -28.725 51.515 -28.395 51.845 ;
        RECT -28.725 50.155 -28.395 50.485 ;
        RECT -28.725 48.795 -28.395 49.125 ;
        RECT -28.725 47.435 -28.395 47.765 ;
        RECT -28.725 46.075 -28.395 46.405 ;
        RECT -28.725 44.715 -28.395 45.045 ;
        RECT -28.725 43.355 -28.395 43.685 ;
        RECT -28.725 41.995 -28.395 42.325 ;
        RECT -28.725 40.635 -28.395 40.965 ;
        RECT -28.725 39.275 -28.395 39.605 ;
        RECT -28.725 37.915 -28.395 38.245 ;
        RECT -28.725 36.555 -28.395 36.885 ;
        RECT -28.725 35.195 -28.395 35.525 ;
        RECT -28.725 33.835 -28.395 34.165 ;
        RECT -28.725 32.475 -28.395 32.805 ;
        RECT -28.725 31.115 -28.395 31.445 ;
        RECT -28.725 29.755 -28.395 30.085 ;
        RECT -28.725 28.395 -28.395 28.725 ;
        RECT -28.725 27.035 -28.395 27.365 ;
        RECT -28.725 25.675 -28.395 26.005 ;
        RECT -28.725 24.315 -28.395 24.645 ;
        RECT -28.725 22.955 -28.395 23.285 ;
        RECT -28.725 21.595 -28.395 21.925 ;
        RECT -28.725 20.235 -28.395 20.565 ;
        RECT -28.725 18.875 -28.395 19.205 ;
        RECT -28.725 17.515 -28.395 17.845 ;
        RECT -28.725 16.155 -28.395 16.485 ;
        RECT -28.725 14.795 -28.395 15.125 ;
        RECT -28.725 13.435 -28.395 13.765 ;
        RECT -28.725 12.075 -28.395 12.405 ;
        RECT -28.725 10.715 -28.395 11.045 ;
        RECT -28.725 9.355 -28.395 9.685 ;
        RECT -28.725 7.995 -28.395 8.325 ;
        RECT -28.725 6.635 -28.395 6.965 ;
        RECT -28.725 5.275 -28.395 5.605 ;
        RECT -28.725 3.915 -28.395 4.245 ;
        RECT -28.725 2.555 -28.395 2.885 ;
        RECT -28.725 1.195 -28.395 1.525 ;
    END
    PORT
      LAYER met3 ;
        RECT -38.245 241.32 -37.915 242.45 ;
        RECT -38.245 239.195 -37.915 239.525 ;
        RECT -38.245 237.835 -37.915 238.165 ;
        RECT -38.245 236.475 -37.915 236.805 ;
        RECT -38.245 235.115 -37.915 235.445 ;
        RECT -38.245 233.755 -37.915 234.085 ;
        RECT -38.245 232.395 -37.915 232.725 ;
        RECT -38.245 231.035 -37.915 231.365 ;
        RECT -38.245 229.675 -37.915 230.005 ;
        RECT -38.245 228.315 -37.915 228.645 ;
        RECT -38.245 226.955 -37.915 227.285 ;
        RECT -38.245 225.595 -37.915 225.925 ;
        RECT -38.245 224.235 -37.915 224.565 ;
        RECT -38.245 222.875 -37.915 223.205 ;
        RECT -38.245 221.515 -37.915 221.845 ;
        RECT -38.245 220.155 -37.915 220.485 ;
        RECT -38.245 218.795 -37.915 219.125 ;
        RECT -38.245 217.435 -37.915 217.765 ;
        RECT -38.245 216.075 -37.915 216.405 ;
        RECT -38.245 214.715 -37.915 215.045 ;
        RECT -38.245 213.355 -37.915 213.685 ;
        RECT -38.245 211.995 -37.915 212.325 ;
        RECT -38.245 210.635 -37.915 210.965 ;
        RECT -38.245 209.275 -37.915 209.605 ;
        RECT -38.245 207.915 -37.915 208.245 ;
        RECT -38.245 206.555 -37.915 206.885 ;
        RECT -38.245 205.195 -37.915 205.525 ;
        RECT -38.245 203.835 -37.915 204.165 ;
        RECT -38.245 202.475 -37.915 202.805 ;
        RECT -38.245 201.115 -37.915 201.445 ;
        RECT -38.245 199.755 -37.915 200.085 ;
        RECT -38.245 198.395 -37.915 198.725 ;
        RECT -38.245 197.035 -37.915 197.365 ;
        RECT -38.245 195.675 -37.915 196.005 ;
        RECT -38.245 194.315 -37.915 194.645 ;
        RECT -38.245 192.955 -37.915 193.285 ;
        RECT -38.245 191.595 -37.915 191.925 ;
        RECT -38.245 190.235 -37.915 190.565 ;
        RECT -38.245 188.875 -37.915 189.205 ;
        RECT -38.245 187.515 -37.915 187.845 ;
        RECT -38.245 186.155 -37.915 186.485 ;
        RECT -38.245 184.795 -37.915 185.125 ;
        RECT -38.245 183.435 -37.915 183.765 ;
        RECT -38.245 182.075 -37.915 182.405 ;
        RECT -38.245 180.715 -37.915 181.045 ;
        RECT -38.245 179.355 -37.915 179.685 ;
        RECT -38.245 177.995 -37.915 178.325 ;
        RECT -38.245 176.635 -37.915 176.965 ;
        RECT -38.245 175.275 -37.915 175.605 ;
        RECT -38.245 173.915 -37.915 174.245 ;
        RECT -38.245 172.555 -37.915 172.885 ;
        RECT -38.245 171.195 -37.915 171.525 ;
        RECT -38.245 169.835 -37.915 170.165 ;
        RECT -38.245 168.475 -37.915 168.805 ;
        RECT -38.245 167.115 -37.915 167.445 ;
        RECT -38.245 165.755 -37.915 166.085 ;
        RECT -38.245 164.395 -37.915 164.725 ;
        RECT -38.245 163.035 -37.915 163.365 ;
        RECT -38.245 161.675 -37.915 162.005 ;
        RECT -38.245 160.315 -37.915 160.645 ;
        RECT -38.245 158.955 -37.915 159.285 ;
        RECT -38.245 157.595 -37.915 157.925 ;
        RECT -38.245 156.235 -37.915 156.565 ;
        RECT -38.245 154.875 -37.915 155.205 ;
        RECT -38.245 153.515 -37.915 153.845 ;
        RECT -38.245 152.155 -37.915 152.485 ;
        RECT -38.245 150.795 -37.915 151.125 ;
        RECT -38.245 149.435 -37.915 149.765 ;
        RECT -38.245 148.075 -37.915 148.405 ;
        RECT -38.245 146.715 -37.915 147.045 ;
        RECT -38.245 145.355 -37.915 145.685 ;
        RECT -38.245 143.995 -37.915 144.325 ;
        RECT -38.245 142.635 -37.915 142.965 ;
        RECT -38.245 141.275 -37.915 141.605 ;
        RECT -38.245 139.915 -37.915 140.245 ;
        RECT -38.245 138.555 -37.915 138.885 ;
        RECT -38.245 137.195 -37.915 137.525 ;
        RECT -38.245 135.835 -37.915 136.165 ;
        RECT -38.245 134.475 -37.915 134.805 ;
        RECT -38.245 133.115 -37.915 133.445 ;
        RECT -38.245 131.755 -37.915 132.085 ;
        RECT -38.245 130.395 -37.915 130.725 ;
        RECT -38.245 129.035 -37.915 129.365 ;
        RECT -38.245 127.675 -37.915 128.005 ;
        RECT -38.245 126.315 -37.915 126.645 ;
        RECT -38.245 124.955 -37.915 125.285 ;
        RECT -38.245 123.595 -37.915 123.925 ;
        RECT -38.245 122.235 -37.915 122.565 ;
        RECT -38.245 120.875 -37.915 121.205 ;
        RECT -38.245 119.515 -37.915 119.845 ;
        RECT -38.245 118.155 -37.915 118.485 ;
        RECT -38.245 116.795 -37.915 117.125 ;
        RECT -38.245 115.435 -37.915 115.765 ;
        RECT -38.245 114.075 -37.915 114.405 ;
        RECT -38.245 112.715 -37.915 113.045 ;
        RECT -38.245 111.355 -37.915 111.685 ;
        RECT -38.245 109.995 -37.915 110.325 ;
        RECT -38.245 108.635 -37.915 108.965 ;
        RECT -38.245 107.275 -37.915 107.605 ;
        RECT -38.245 105.915 -37.915 106.245 ;
        RECT -38.245 104.555 -37.915 104.885 ;
        RECT -38.245 103.195 -37.915 103.525 ;
        RECT -38.245 101.835 -37.915 102.165 ;
        RECT -38.245 100.475 -37.915 100.805 ;
        RECT -38.245 99.115 -37.915 99.445 ;
        RECT -38.245 97.755 -37.915 98.085 ;
        RECT -38.245 96.395 -37.915 96.725 ;
        RECT -38.245 95.035 -37.915 95.365 ;
        RECT -38.245 93.675 -37.915 94.005 ;
        RECT -38.245 92.315 -37.915 92.645 ;
        RECT -38.245 90.955 -37.915 91.285 ;
        RECT -38.245 89.595 -37.915 89.925 ;
        RECT -38.245 88.235 -37.915 88.565 ;
        RECT -38.245 86.875 -37.915 87.205 ;
        RECT -38.245 85.515 -37.915 85.845 ;
        RECT -38.245 84.155 -37.915 84.485 ;
        RECT -38.245 82.795 -37.915 83.125 ;
        RECT -38.245 81.435 -37.915 81.765 ;
        RECT -38.245 80.075 -37.915 80.405 ;
        RECT -38.245 78.715 -37.915 79.045 ;
        RECT -38.245 77.355 -37.915 77.685 ;
        RECT -38.245 75.995 -37.915 76.325 ;
        RECT -38.245 74.635 -37.915 74.965 ;
        RECT -38.245 73.275 -37.915 73.605 ;
        RECT -38.245 71.915 -37.915 72.245 ;
        RECT -38.245 70.555 -37.915 70.885 ;
        RECT -38.245 69.195 -37.915 69.525 ;
        RECT -38.245 67.835 -37.915 68.165 ;
        RECT -38.245 66.475 -37.915 66.805 ;
        RECT -38.245 65.115 -37.915 65.445 ;
        RECT -38.245 63.755 -37.915 64.085 ;
        RECT -38.245 62.395 -37.915 62.725 ;
        RECT -38.245 61.035 -37.915 61.365 ;
        RECT -38.245 59.675 -37.915 60.005 ;
        RECT -38.245 58.315 -37.915 58.645 ;
        RECT -38.245 56.955 -37.915 57.285 ;
        RECT -38.245 55.595 -37.915 55.925 ;
        RECT -38.245 54.235 -37.915 54.565 ;
        RECT -38.245 52.875 -37.915 53.205 ;
        RECT -38.245 51.515 -37.915 51.845 ;
        RECT -38.245 50.155 -37.915 50.485 ;
        RECT -38.245 48.795 -37.915 49.125 ;
        RECT -38.245 47.435 -37.915 47.765 ;
        RECT -38.245 46.075 -37.915 46.405 ;
        RECT -38.245 44.715 -37.915 45.045 ;
        RECT -38.245 43.355 -37.915 43.685 ;
        RECT -38.245 41.995 -37.915 42.325 ;
        RECT -38.245 40.635 -37.915 40.965 ;
        RECT -38.245 39.275 -37.915 39.605 ;
        RECT -38.245 37.915 -37.915 38.245 ;
        RECT -38.245 36.555 -37.915 36.885 ;
        RECT -38.245 35.195 -37.915 35.525 ;
        RECT -38.245 33.835 -37.915 34.165 ;
        RECT -38.245 32.475 -37.915 32.805 ;
        RECT -38.245 31.115 -37.915 31.445 ;
        RECT -38.245 29.755 -37.915 30.085 ;
        RECT -38.245 28.395 -37.915 28.725 ;
        RECT -38.245 27.035 -37.915 27.365 ;
        RECT -38.245 25.675 -37.915 26.005 ;
        RECT -38.245 24.315 -37.915 24.645 ;
        RECT -38.245 22.955 -37.915 23.285 ;
        RECT -38.245 21.595 -37.915 21.925 ;
        RECT -38.245 20.235 -37.915 20.565 ;
        RECT -38.245 18.875 -37.915 19.205 ;
        RECT -38.245 17.515 -37.915 17.845 ;
        RECT -38.245 16.155 -37.915 16.485 ;
        RECT -38.245 14.795 -37.915 15.125 ;
        RECT -38.245 13.435 -37.915 13.765 ;
        RECT -38.245 12.075 -37.915 12.405 ;
        RECT -38.245 10.715 -37.915 11.045 ;
        RECT -38.245 9.355 -37.915 9.685 ;
        RECT -38.245 7.995 -37.915 8.325 ;
        RECT -38.245 6.635 -37.915 6.965 ;
        RECT -38.245 5.275 -37.915 5.605 ;
        RECT -38.245 3.915 -37.915 4.245 ;
        RECT -38.245 2.555 -37.915 2.885 ;
        RECT -38.245 1.195 -37.915 1.525 ;
        RECT -38.245 -0.165 -37.915 0.165 ;
        RECT -38.245 -2.885 -37.915 -2.555 ;
        RECT -38.245 -4.245 -37.915 -3.915 ;
        RECT -38.245 -11.045 -37.915 -10.715 ;
        RECT -38.245 -15.125 -37.915 -14.795 ;
        RECT -38.245 -16.485 -37.915 -16.155 ;
        RECT -38.245 -17.845 -37.915 -17.515 ;
        RECT -38.245 -19.205 -37.915 -18.875 ;
        RECT -38.245 -20.565 -37.915 -20.235 ;
        RECT -38.245 -21.925 -37.915 -21.595 ;
        RECT -38.245 -23.285 -37.915 -22.955 ;
        RECT -38.245 -24.645 -37.915 -24.315 ;
        RECT -38.245 -31.445 -37.915 -31.115 ;
        RECT -38.245 -32.805 -37.915 -32.475 ;
        RECT -38.245 -35.525 -37.915 -35.195 ;
        RECT -38.245 -36.885 -37.915 -36.555 ;
        RECT -38.245 -37.93 -37.915 -37.6 ;
        RECT -38.245 -40.965 -37.915 -40.635 ;
        RECT -38.245 -42.77 -37.915 -42.44 ;
        RECT -38.245 -43.685 -37.915 -43.355 ;
        RECT -38.245 -50.485 -37.915 -50.155 ;
        RECT -38.245 -51.845 -37.915 -51.515 ;
        RECT -38.245 -53.205 -37.915 -52.875 ;
        RECT -38.245 -54.565 -37.915 -54.235 ;
        RECT -38.245 -55.925 -37.915 -55.595 ;
        RECT -38.245 -57.285 -37.915 -56.955 ;
        RECT -38.245 -58.645 -37.915 -58.315 ;
        RECT -38.245 -60.005 -37.915 -59.675 ;
        RECT -38.245 -61.365 -37.915 -61.035 ;
        RECT -38.245 -64.085 -37.915 -63.755 ;
        RECT -38.245 -65.445 -37.915 -65.115 ;
        RECT -38.245 -66.805 -37.915 -66.475 ;
        RECT -38.245 -68.165 -37.915 -67.835 ;
        RECT -38.245 -69.525 -37.915 -69.195 ;
        RECT -38.245 -70.885 -37.915 -70.555 ;
        RECT -38.245 -72.245 -37.915 -71.915 ;
        RECT -38.245 -73.605 -37.915 -73.275 ;
        RECT -38.245 -74.965 -37.915 -74.635 ;
        RECT -38.245 -76.325 -37.915 -75.995 ;
        RECT -38.245 -77.685 -37.915 -77.355 ;
        RECT -38.245 -79.045 -37.915 -78.715 ;
        RECT -38.245 -80.405 -37.915 -80.075 ;
        RECT -38.245 -81.765 -37.915 -81.435 ;
        RECT -38.245 -83.125 -37.915 -82.795 ;
        RECT -38.245 -84.485 -37.915 -84.155 ;
        RECT -38.245 -85.845 -37.915 -85.515 ;
        RECT -38.245 -87.205 -37.915 -86.875 ;
        RECT -38.245 -88.565 -37.915 -88.235 ;
        RECT -38.245 -89.925 -37.915 -89.595 ;
        RECT -38.245 -92.645 -37.915 -92.315 ;
        RECT -38.245 -94.005 -37.915 -93.675 ;
        RECT -38.245 -95.365 -37.915 -95.035 ;
        RECT -38.245 -96.725 -37.915 -96.395 ;
        RECT -38.245 -98.73 -37.915 -98.4 ;
        RECT -38.245 -99.445 -37.915 -99.115 ;
        RECT -38.245 -102.165 -37.915 -101.835 ;
        RECT -38.245 -103.525 -37.915 -103.195 ;
        RECT -38.245 -104.885 -37.915 -104.555 ;
        RECT -38.245 -106.87 -37.915 -106.54 ;
        RECT -38.245 -107.605 -37.915 -107.275 ;
        RECT -38.245 -108.965 -37.915 -108.635 ;
        RECT -38.245 -113.045 -37.915 -112.715 ;
        RECT -38.245 -114.405 -37.915 -114.075 ;
        RECT -38.245 -115.765 -37.915 -115.435 ;
        RECT -38.245 -117.125 -37.915 -116.795 ;
        RECT -38.245 -118.485 -37.915 -118.155 ;
        RECT -38.245 -122.565 -37.915 -122.235 ;
        RECT -38.245 -123.925 -37.915 -123.595 ;
        RECT -38.245 -125.285 -37.915 -124.955 ;
        RECT -38.245 -126.645 -37.915 -126.315 ;
        RECT -38.245 -128.005 -37.915 -127.675 ;
        RECT -38.245 -129.365 -37.915 -129.035 ;
        RECT -38.245 -133.445 -37.915 -133.115 ;
        RECT -38.245 -134.805 -37.915 -134.475 ;
        RECT -38.245 -136.165 -37.915 -135.835 ;
        RECT -38.245 -137.525 -37.915 -137.195 ;
        RECT -38.245 -138.885 -37.915 -138.555 ;
        RECT -38.245 -140.245 -37.915 -139.915 ;
        RECT -38.245 -141.605 -37.915 -141.275 ;
        RECT -38.245 -142.965 -37.915 -142.635 ;
        RECT -38.245 -144.325 -37.915 -143.995 ;
        RECT -38.245 -145.685 -37.915 -145.355 ;
        RECT -38.245 -147.045 -37.915 -146.715 ;
        RECT -38.245 -148.405 -37.915 -148.075 ;
        RECT -38.245 -151.125 -37.915 -150.795 ;
        RECT -38.245 -152.485 -37.915 -152.155 ;
        RECT -38.245 -155.205 -37.915 -154.875 ;
        RECT -38.245 -156.565 -37.915 -156.235 ;
        RECT -38.245 -157.925 -37.915 -157.595 ;
        RECT -38.245 -159.285 -37.915 -158.955 ;
        RECT -38.245 -160.645 -37.915 -160.315 ;
        RECT -38.245 -162.005 -37.915 -161.675 ;
        RECT -38.245 -163.365 -37.915 -163.035 ;
        RECT -38.245 -164.725 -37.915 -164.395 ;
        RECT -38.245 -166.085 -37.915 -165.755 ;
        RECT -38.245 -167.445 -37.915 -167.115 ;
        RECT -38.245 -170.165 -37.915 -169.835 ;
        RECT -38.245 -172.885 -37.915 -172.555 ;
        RECT -38.245 -174.245 -37.915 -173.915 ;
        RECT -38.245 -175.725 -37.915 -175.395 ;
        RECT -38.245 -176.965 -37.915 -176.635 ;
        RECT -38.245 -178.325 -37.915 -177.995 ;
        RECT -38.245 -180.57 -37.915 -179.44 ;
        RECT -38.24 -180.685 -37.92 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -36.885 241.32 -36.555 242.45 ;
        RECT -36.885 239.195 -36.555 239.525 ;
        RECT -36.885 237.835 -36.555 238.165 ;
        RECT -36.885 236.475 -36.555 236.805 ;
        RECT -36.885 235.115 -36.555 235.445 ;
        RECT -36.885 233.755 -36.555 234.085 ;
        RECT -36.885 232.395 -36.555 232.725 ;
        RECT -36.885 231.035 -36.555 231.365 ;
        RECT -36.885 229.675 -36.555 230.005 ;
        RECT -36.885 228.315 -36.555 228.645 ;
        RECT -36.885 226.955 -36.555 227.285 ;
        RECT -36.885 225.595 -36.555 225.925 ;
        RECT -36.885 224.235 -36.555 224.565 ;
        RECT -36.885 222.875 -36.555 223.205 ;
        RECT -36.885 221.515 -36.555 221.845 ;
        RECT -36.885 220.155 -36.555 220.485 ;
        RECT -36.885 218.795 -36.555 219.125 ;
        RECT -36.885 217.435 -36.555 217.765 ;
        RECT -36.885 216.075 -36.555 216.405 ;
        RECT -36.885 214.715 -36.555 215.045 ;
        RECT -36.885 213.355 -36.555 213.685 ;
        RECT -36.885 211.995 -36.555 212.325 ;
        RECT -36.885 210.635 -36.555 210.965 ;
        RECT -36.885 209.275 -36.555 209.605 ;
        RECT -36.885 207.915 -36.555 208.245 ;
        RECT -36.885 206.555 -36.555 206.885 ;
        RECT -36.885 205.195 -36.555 205.525 ;
        RECT -36.885 203.835 -36.555 204.165 ;
        RECT -36.885 202.475 -36.555 202.805 ;
        RECT -36.885 201.115 -36.555 201.445 ;
        RECT -36.885 199.755 -36.555 200.085 ;
        RECT -36.885 198.395 -36.555 198.725 ;
        RECT -36.885 197.035 -36.555 197.365 ;
        RECT -36.885 195.675 -36.555 196.005 ;
        RECT -36.885 194.315 -36.555 194.645 ;
        RECT -36.885 192.955 -36.555 193.285 ;
        RECT -36.885 191.595 -36.555 191.925 ;
        RECT -36.885 190.235 -36.555 190.565 ;
        RECT -36.885 188.875 -36.555 189.205 ;
        RECT -36.885 187.515 -36.555 187.845 ;
        RECT -36.885 186.155 -36.555 186.485 ;
        RECT -36.885 184.795 -36.555 185.125 ;
        RECT -36.885 183.435 -36.555 183.765 ;
        RECT -36.885 182.075 -36.555 182.405 ;
        RECT -36.885 180.715 -36.555 181.045 ;
        RECT -36.885 179.355 -36.555 179.685 ;
        RECT -36.885 177.995 -36.555 178.325 ;
        RECT -36.885 176.635 -36.555 176.965 ;
        RECT -36.885 175.275 -36.555 175.605 ;
        RECT -36.885 173.915 -36.555 174.245 ;
        RECT -36.885 172.555 -36.555 172.885 ;
        RECT -36.885 171.195 -36.555 171.525 ;
        RECT -36.885 169.835 -36.555 170.165 ;
        RECT -36.885 168.475 -36.555 168.805 ;
        RECT -36.885 167.115 -36.555 167.445 ;
        RECT -36.885 165.755 -36.555 166.085 ;
        RECT -36.885 164.395 -36.555 164.725 ;
        RECT -36.885 163.035 -36.555 163.365 ;
        RECT -36.885 161.675 -36.555 162.005 ;
        RECT -36.885 160.315 -36.555 160.645 ;
        RECT -36.885 158.955 -36.555 159.285 ;
        RECT -36.885 157.595 -36.555 157.925 ;
        RECT -36.885 156.235 -36.555 156.565 ;
        RECT -36.885 154.875 -36.555 155.205 ;
        RECT -36.885 153.515 -36.555 153.845 ;
        RECT -36.885 152.155 -36.555 152.485 ;
        RECT -36.885 150.795 -36.555 151.125 ;
        RECT -36.885 149.435 -36.555 149.765 ;
        RECT -36.885 148.075 -36.555 148.405 ;
        RECT -36.885 146.715 -36.555 147.045 ;
        RECT -36.885 145.355 -36.555 145.685 ;
        RECT -36.885 143.995 -36.555 144.325 ;
        RECT -36.885 142.635 -36.555 142.965 ;
        RECT -36.885 141.275 -36.555 141.605 ;
        RECT -36.885 139.915 -36.555 140.245 ;
        RECT -36.885 138.555 -36.555 138.885 ;
        RECT -36.885 137.195 -36.555 137.525 ;
        RECT -36.885 135.835 -36.555 136.165 ;
        RECT -36.885 134.475 -36.555 134.805 ;
        RECT -36.885 133.115 -36.555 133.445 ;
        RECT -36.885 131.755 -36.555 132.085 ;
        RECT -36.885 130.395 -36.555 130.725 ;
        RECT -36.885 129.035 -36.555 129.365 ;
        RECT -36.885 127.675 -36.555 128.005 ;
        RECT -36.885 126.315 -36.555 126.645 ;
        RECT -36.885 124.955 -36.555 125.285 ;
        RECT -36.885 123.595 -36.555 123.925 ;
        RECT -36.885 122.235 -36.555 122.565 ;
        RECT -36.885 120.875 -36.555 121.205 ;
        RECT -36.885 119.515 -36.555 119.845 ;
        RECT -36.885 118.155 -36.555 118.485 ;
        RECT -36.885 116.795 -36.555 117.125 ;
        RECT -36.885 115.435 -36.555 115.765 ;
        RECT -36.885 114.075 -36.555 114.405 ;
        RECT -36.885 112.715 -36.555 113.045 ;
        RECT -36.885 111.355 -36.555 111.685 ;
        RECT -36.885 109.995 -36.555 110.325 ;
        RECT -36.885 108.635 -36.555 108.965 ;
        RECT -36.885 107.275 -36.555 107.605 ;
        RECT -36.885 105.915 -36.555 106.245 ;
        RECT -36.885 104.555 -36.555 104.885 ;
        RECT -36.885 103.195 -36.555 103.525 ;
        RECT -36.885 101.835 -36.555 102.165 ;
        RECT -36.885 100.475 -36.555 100.805 ;
        RECT -36.885 99.115 -36.555 99.445 ;
        RECT -36.885 97.755 -36.555 98.085 ;
        RECT -36.885 96.395 -36.555 96.725 ;
        RECT -36.885 95.035 -36.555 95.365 ;
        RECT -36.885 93.675 -36.555 94.005 ;
        RECT -36.885 92.315 -36.555 92.645 ;
        RECT -36.885 90.955 -36.555 91.285 ;
        RECT -36.885 89.595 -36.555 89.925 ;
        RECT -36.885 88.235 -36.555 88.565 ;
        RECT -36.885 86.875 -36.555 87.205 ;
        RECT -36.885 85.515 -36.555 85.845 ;
        RECT -36.885 84.155 -36.555 84.485 ;
        RECT -36.885 82.795 -36.555 83.125 ;
        RECT -36.885 81.435 -36.555 81.765 ;
        RECT -36.885 80.075 -36.555 80.405 ;
        RECT -36.885 78.715 -36.555 79.045 ;
        RECT -36.885 77.355 -36.555 77.685 ;
        RECT -36.885 75.995 -36.555 76.325 ;
        RECT -36.885 74.635 -36.555 74.965 ;
        RECT -36.885 73.275 -36.555 73.605 ;
        RECT -36.885 71.915 -36.555 72.245 ;
        RECT -36.885 70.555 -36.555 70.885 ;
        RECT -36.885 69.195 -36.555 69.525 ;
        RECT -36.885 67.835 -36.555 68.165 ;
        RECT -36.885 66.475 -36.555 66.805 ;
        RECT -36.885 65.115 -36.555 65.445 ;
        RECT -36.885 63.755 -36.555 64.085 ;
        RECT -36.885 62.395 -36.555 62.725 ;
        RECT -36.885 61.035 -36.555 61.365 ;
        RECT -36.885 59.675 -36.555 60.005 ;
        RECT -36.885 58.315 -36.555 58.645 ;
        RECT -36.885 56.955 -36.555 57.285 ;
        RECT -36.885 55.595 -36.555 55.925 ;
        RECT -36.885 54.235 -36.555 54.565 ;
        RECT -36.885 52.875 -36.555 53.205 ;
        RECT -36.885 51.515 -36.555 51.845 ;
        RECT -36.885 50.155 -36.555 50.485 ;
        RECT -36.885 48.795 -36.555 49.125 ;
        RECT -36.885 47.435 -36.555 47.765 ;
        RECT -36.885 46.075 -36.555 46.405 ;
        RECT -36.885 44.715 -36.555 45.045 ;
        RECT -36.885 43.355 -36.555 43.685 ;
        RECT -36.885 41.995 -36.555 42.325 ;
        RECT -36.885 40.635 -36.555 40.965 ;
        RECT -36.885 39.275 -36.555 39.605 ;
        RECT -36.885 37.915 -36.555 38.245 ;
        RECT -36.885 36.555 -36.555 36.885 ;
        RECT -36.885 35.195 -36.555 35.525 ;
        RECT -36.885 33.835 -36.555 34.165 ;
        RECT -36.885 32.475 -36.555 32.805 ;
        RECT -36.885 31.115 -36.555 31.445 ;
        RECT -36.885 29.755 -36.555 30.085 ;
        RECT -36.885 28.395 -36.555 28.725 ;
        RECT -36.885 27.035 -36.555 27.365 ;
        RECT -36.885 25.675 -36.555 26.005 ;
        RECT -36.885 24.315 -36.555 24.645 ;
        RECT -36.885 22.955 -36.555 23.285 ;
        RECT -36.885 21.595 -36.555 21.925 ;
        RECT -36.885 20.235 -36.555 20.565 ;
        RECT -36.885 18.875 -36.555 19.205 ;
        RECT -36.885 17.515 -36.555 17.845 ;
        RECT -36.885 16.155 -36.555 16.485 ;
        RECT -36.885 14.795 -36.555 15.125 ;
        RECT -36.885 13.435 -36.555 13.765 ;
        RECT -36.885 12.075 -36.555 12.405 ;
        RECT -36.885 10.715 -36.555 11.045 ;
        RECT -36.885 9.355 -36.555 9.685 ;
        RECT -36.885 7.995 -36.555 8.325 ;
        RECT -36.885 6.635 -36.555 6.965 ;
        RECT -36.885 5.275 -36.555 5.605 ;
        RECT -36.885 3.915 -36.555 4.245 ;
        RECT -36.885 2.555 -36.555 2.885 ;
        RECT -36.885 1.195 -36.555 1.525 ;
        RECT -36.885 -0.165 -36.555 0.165 ;
        RECT -36.885 -2.885 -36.555 -2.555 ;
        RECT -36.885 -11.045 -36.555 -10.715 ;
        RECT -36.885 -15.125 -36.555 -14.795 ;
        RECT -36.885 -16.485 -36.555 -16.155 ;
        RECT -36.885 -17.845 -36.555 -17.515 ;
        RECT -36.885 -19.205 -36.555 -18.875 ;
        RECT -36.885 -20.565 -36.555 -20.235 ;
        RECT -36.885 -21.925 -36.555 -21.595 ;
        RECT -36.885 -23.285 -36.555 -22.955 ;
        RECT -36.885 -24.645 -36.555 -24.315 ;
        RECT -36.885 -31.445 -36.555 -31.115 ;
        RECT -36.885 -32.805 -36.555 -32.475 ;
        RECT -36.885 -35.525 -36.555 -35.195 ;
        RECT -36.885 -36.885 -36.555 -36.555 ;
        RECT -36.885 -37.93 -36.555 -37.6 ;
        RECT -36.885 -40.965 -36.555 -40.635 ;
        RECT -36.885 -42.77 -36.555 -42.44 ;
        RECT -36.885 -43.685 -36.555 -43.355 ;
        RECT -36.885 -50.485 -36.555 -50.155 ;
        RECT -36.885 -51.845 -36.555 -51.515 ;
        RECT -36.885 -53.205 -36.555 -52.875 ;
        RECT -36.885 -54.565 -36.555 -54.235 ;
        RECT -36.885 -55.925 -36.555 -55.595 ;
        RECT -36.885 -57.285 -36.555 -56.955 ;
        RECT -36.885 -58.645 -36.555 -58.315 ;
        RECT -36.885 -60.005 -36.555 -59.675 ;
        RECT -36.885 -61.365 -36.555 -61.035 ;
        RECT -36.885 -64.085 -36.555 -63.755 ;
        RECT -36.885 -65.445 -36.555 -65.115 ;
        RECT -36.885 -66.805 -36.555 -66.475 ;
        RECT -36.885 -68.165 -36.555 -67.835 ;
        RECT -36.885 -69.525 -36.555 -69.195 ;
        RECT -36.885 -70.885 -36.555 -70.555 ;
        RECT -36.885 -72.245 -36.555 -71.915 ;
        RECT -36.885 -73.605 -36.555 -73.275 ;
        RECT -36.885 -74.965 -36.555 -74.635 ;
        RECT -36.885 -76.325 -36.555 -75.995 ;
        RECT -36.885 -77.685 -36.555 -77.355 ;
        RECT -36.885 -79.045 -36.555 -78.715 ;
        RECT -36.885 -80.405 -36.555 -80.075 ;
        RECT -36.885 -81.765 -36.555 -81.435 ;
        RECT -36.885 -83.125 -36.555 -82.795 ;
        RECT -36.885 -84.485 -36.555 -84.155 ;
        RECT -36.885 -85.845 -36.555 -85.515 ;
        RECT -36.885 -87.205 -36.555 -86.875 ;
        RECT -36.885 -88.565 -36.555 -88.235 ;
        RECT -36.885 -89.925 -36.555 -89.595 ;
        RECT -36.885 -92.645 -36.555 -92.315 ;
        RECT -36.885 -94.005 -36.555 -93.675 ;
        RECT -36.885 -95.365 -36.555 -95.035 ;
        RECT -36.885 -96.725 -36.555 -96.395 ;
        RECT -36.885 -98.73 -36.555 -98.4 ;
        RECT -36.885 -99.445 -36.555 -99.115 ;
        RECT -36.885 -102.165 -36.555 -101.835 ;
        RECT -36.885 -103.525 -36.555 -103.195 ;
        RECT -36.885 -104.885 -36.555 -104.555 ;
        RECT -36.885 -106.87 -36.555 -106.54 ;
        RECT -36.885 -107.605 -36.555 -107.275 ;
        RECT -36.885 -108.965 -36.555 -108.635 ;
        RECT -36.885 -113.045 -36.555 -112.715 ;
        RECT -36.885 -114.405 -36.555 -114.075 ;
        RECT -36.885 -115.765 -36.555 -115.435 ;
        RECT -36.885 -117.125 -36.555 -116.795 ;
        RECT -36.885 -118.485 -36.555 -118.155 ;
        RECT -36.885 -122.565 -36.555 -122.235 ;
        RECT -36.885 -123.925 -36.555 -123.595 ;
        RECT -36.885 -125.285 -36.555 -124.955 ;
        RECT -36.885 -126.645 -36.555 -126.315 ;
        RECT -36.885 -128.005 -36.555 -127.675 ;
        RECT -36.885 -129.365 -36.555 -129.035 ;
        RECT -36.885 -133.445 -36.555 -133.115 ;
        RECT -36.885 -134.805 -36.555 -134.475 ;
        RECT -36.885 -136.165 -36.555 -135.835 ;
        RECT -36.885 -137.525 -36.555 -137.195 ;
        RECT -36.885 -138.885 -36.555 -138.555 ;
        RECT -36.885 -140.245 -36.555 -139.915 ;
        RECT -36.885 -141.605 -36.555 -141.275 ;
        RECT -36.885 -142.965 -36.555 -142.635 ;
        RECT -36.885 -144.325 -36.555 -143.995 ;
        RECT -36.885 -145.685 -36.555 -145.355 ;
        RECT -36.885 -147.045 -36.555 -146.715 ;
        RECT -36.885 -148.405 -36.555 -148.075 ;
        RECT -36.885 -151.125 -36.555 -150.795 ;
        RECT -36.885 -152.485 -36.555 -152.155 ;
        RECT -36.885 -156.565 -36.555 -156.235 ;
        RECT -36.885 -157.925 -36.555 -157.595 ;
        RECT -36.885 -159.285 -36.555 -158.955 ;
        RECT -36.885 -160.645 -36.555 -160.315 ;
        RECT -36.885 -162.005 -36.555 -161.675 ;
        RECT -36.885 -163.365 -36.555 -163.035 ;
        RECT -36.885 -164.725 -36.555 -164.395 ;
        RECT -36.885 -166.085 -36.555 -165.755 ;
        RECT -36.885 -167.445 -36.555 -167.115 ;
        RECT -36.885 -170.165 -36.555 -169.835 ;
        RECT -36.885 -172.885 -36.555 -172.555 ;
        RECT -36.885 -174.245 -36.555 -173.915 ;
        RECT -36.885 -175.725 -36.555 -175.395 ;
        RECT -36.885 -176.965 -36.555 -176.635 ;
        RECT -36.885 -178.325 -36.555 -177.995 ;
        RECT -36.885 -180.57 -36.555 -179.44 ;
        RECT -36.88 -180.685 -36.56 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -35.525 241.32 -35.195 242.45 ;
        RECT -35.525 239.195 -35.195 239.525 ;
        RECT -35.525 237.835 -35.195 238.165 ;
        RECT -35.525 236.475 -35.195 236.805 ;
        RECT -35.525 235.115 -35.195 235.445 ;
        RECT -35.525 233.755 -35.195 234.085 ;
        RECT -35.525 232.395 -35.195 232.725 ;
        RECT -35.525 231.035 -35.195 231.365 ;
        RECT -35.525 229.675 -35.195 230.005 ;
        RECT -35.525 228.315 -35.195 228.645 ;
        RECT -35.525 226.955 -35.195 227.285 ;
        RECT -35.525 225.595 -35.195 225.925 ;
        RECT -35.525 224.235 -35.195 224.565 ;
        RECT -35.525 222.875 -35.195 223.205 ;
        RECT -35.525 221.515 -35.195 221.845 ;
        RECT -35.525 220.155 -35.195 220.485 ;
        RECT -35.525 218.795 -35.195 219.125 ;
        RECT -35.525 217.435 -35.195 217.765 ;
        RECT -35.525 216.075 -35.195 216.405 ;
        RECT -35.525 214.715 -35.195 215.045 ;
        RECT -35.525 213.355 -35.195 213.685 ;
        RECT -35.525 211.995 -35.195 212.325 ;
        RECT -35.525 210.635 -35.195 210.965 ;
        RECT -35.525 209.275 -35.195 209.605 ;
        RECT -35.525 207.915 -35.195 208.245 ;
        RECT -35.525 206.555 -35.195 206.885 ;
        RECT -35.525 205.195 -35.195 205.525 ;
        RECT -35.525 203.835 -35.195 204.165 ;
        RECT -35.525 202.475 -35.195 202.805 ;
        RECT -35.525 201.115 -35.195 201.445 ;
        RECT -35.525 199.755 -35.195 200.085 ;
        RECT -35.525 198.395 -35.195 198.725 ;
        RECT -35.525 197.035 -35.195 197.365 ;
        RECT -35.525 195.675 -35.195 196.005 ;
        RECT -35.525 194.315 -35.195 194.645 ;
        RECT -35.525 192.955 -35.195 193.285 ;
        RECT -35.525 191.595 -35.195 191.925 ;
        RECT -35.525 190.235 -35.195 190.565 ;
        RECT -35.525 188.875 -35.195 189.205 ;
        RECT -35.525 187.515 -35.195 187.845 ;
        RECT -35.525 186.155 -35.195 186.485 ;
        RECT -35.525 184.795 -35.195 185.125 ;
        RECT -35.525 183.435 -35.195 183.765 ;
        RECT -35.525 182.075 -35.195 182.405 ;
        RECT -35.525 180.715 -35.195 181.045 ;
        RECT -35.525 179.355 -35.195 179.685 ;
        RECT -35.525 177.995 -35.195 178.325 ;
        RECT -35.525 176.635 -35.195 176.965 ;
        RECT -35.525 175.275 -35.195 175.605 ;
        RECT -35.525 173.915 -35.195 174.245 ;
        RECT -35.525 172.555 -35.195 172.885 ;
        RECT -35.525 171.195 -35.195 171.525 ;
        RECT -35.525 169.835 -35.195 170.165 ;
        RECT -35.525 168.475 -35.195 168.805 ;
        RECT -35.525 167.115 -35.195 167.445 ;
        RECT -35.525 165.755 -35.195 166.085 ;
        RECT -35.525 164.395 -35.195 164.725 ;
        RECT -35.525 163.035 -35.195 163.365 ;
        RECT -35.525 161.675 -35.195 162.005 ;
        RECT -35.525 160.315 -35.195 160.645 ;
        RECT -35.525 158.955 -35.195 159.285 ;
        RECT -35.525 157.595 -35.195 157.925 ;
        RECT -35.525 156.235 -35.195 156.565 ;
        RECT -35.525 154.875 -35.195 155.205 ;
        RECT -35.525 153.515 -35.195 153.845 ;
        RECT -35.525 152.155 -35.195 152.485 ;
        RECT -35.525 150.795 -35.195 151.125 ;
        RECT -35.525 149.435 -35.195 149.765 ;
        RECT -35.525 148.075 -35.195 148.405 ;
        RECT -35.525 146.715 -35.195 147.045 ;
        RECT -35.525 145.355 -35.195 145.685 ;
        RECT -35.525 143.995 -35.195 144.325 ;
        RECT -35.525 142.635 -35.195 142.965 ;
        RECT -35.525 141.275 -35.195 141.605 ;
        RECT -35.525 139.915 -35.195 140.245 ;
        RECT -35.525 138.555 -35.195 138.885 ;
        RECT -35.525 137.195 -35.195 137.525 ;
        RECT -35.525 135.835 -35.195 136.165 ;
        RECT -35.525 134.475 -35.195 134.805 ;
        RECT -35.525 133.115 -35.195 133.445 ;
        RECT -35.525 131.755 -35.195 132.085 ;
        RECT -35.525 130.395 -35.195 130.725 ;
        RECT -35.525 129.035 -35.195 129.365 ;
        RECT -35.525 127.675 -35.195 128.005 ;
        RECT -35.525 126.315 -35.195 126.645 ;
        RECT -35.525 124.955 -35.195 125.285 ;
        RECT -35.525 123.595 -35.195 123.925 ;
        RECT -35.525 122.235 -35.195 122.565 ;
        RECT -35.525 120.875 -35.195 121.205 ;
        RECT -35.525 119.515 -35.195 119.845 ;
        RECT -35.525 118.155 -35.195 118.485 ;
        RECT -35.525 116.795 -35.195 117.125 ;
        RECT -35.525 115.435 -35.195 115.765 ;
        RECT -35.525 114.075 -35.195 114.405 ;
        RECT -35.525 112.715 -35.195 113.045 ;
        RECT -35.525 111.355 -35.195 111.685 ;
        RECT -35.525 109.995 -35.195 110.325 ;
        RECT -35.525 108.635 -35.195 108.965 ;
        RECT -35.525 107.275 -35.195 107.605 ;
        RECT -35.525 105.915 -35.195 106.245 ;
        RECT -35.525 104.555 -35.195 104.885 ;
        RECT -35.525 103.195 -35.195 103.525 ;
        RECT -35.525 101.835 -35.195 102.165 ;
        RECT -35.525 100.475 -35.195 100.805 ;
        RECT -35.525 99.115 -35.195 99.445 ;
        RECT -35.525 97.755 -35.195 98.085 ;
        RECT -35.525 96.395 -35.195 96.725 ;
        RECT -35.525 95.035 -35.195 95.365 ;
        RECT -35.525 93.675 -35.195 94.005 ;
        RECT -35.525 92.315 -35.195 92.645 ;
        RECT -35.525 90.955 -35.195 91.285 ;
        RECT -35.525 89.595 -35.195 89.925 ;
        RECT -35.525 88.235 -35.195 88.565 ;
        RECT -35.525 86.875 -35.195 87.205 ;
        RECT -35.525 85.515 -35.195 85.845 ;
        RECT -35.525 84.155 -35.195 84.485 ;
        RECT -35.525 82.795 -35.195 83.125 ;
        RECT -35.525 81.435 -35.195 81.765 ;
        RECT -35.525 80.075 -35.195 80.405 ;
        RECT -35.525 78.715 -35.195 79.045 ;
        RECT -35.525 77.355 -35.195 77.685 ;
        RECT -35.525 75.995 -35.195 76.325 ;
        RECT -35.525 74.635 -35.195 74.965 ;
        RECT -35.525 73.275 -35.195 73.605 ;
        RECT -35.525 71.915 -35.195 72.245 ;
        RECT -35.525 70.555 -35.195 70.885 ;
        RECT -35.525 69.195 -35.195 69.525 ;
        RECT -35.525 67.835 -35.195 68.165 ;
        RECT -35.525 66.475 -35.195 66.805 ;
        RECT -35.525 65.115 -35.195 65.445 ;
        RECT -35.525 63.755 -35.195 64.085 ;
        RECT -35.525 62.395 -35.195 62.725 ;
        RECT -35.525 61.035 -35.195 61.365 ;
        RECT -35.525 59.675 -35.195 60.005 ;
        RECT -35.525 58.315 -35.195 58.645 ;
        RECT -35.525 56.955 -35.195 57.285 ;
        RECT -35.525 55.595 -35.195 55.925 ;
        RECT -35.525 54.235 -35.195 54.565 ;
        RECT -35.525 52.875 -35.195 53.205 ;
        RECT -35.525 51.515 -35.195 51.845 ;
        RECT -35.525 50.155 -35.195 50.485 ;
        RECT -35.525 48.795 -35.195 49.125 ;
        RECT -35.525 47.435 -35.195 47.765 ;
        RECT -35.525 46.075 -35.195 46.405 ;
        RECT -35.525 44.715 -35.195 45.045 ;
        RECT -35.525 43.355 -35.195 43.685 ;
        RECT -35.525 41.995 -35.195 42.325 ;
        RECT -35.525 40.635 -35.195 40.965 ;
        RECT -35.525 39.275 -35.195 39.605 ;
        RECT -35.525 37.915 -35.195 38.245 ;
        RECT -35.525 36.555 -35.195 36.885 ;
        RECT -35.525 35.195 -35.195 35.525 ;
        RECT -35.525 33.835 -35.195 34.165 ;
        RECT -35.525 32.475 -35.195 32.805 ;
        RECT -35.525 31.115 -35.195 31.445 ;
        RECT -35.525 29.755 -35.195 30.085 ;
        RECT -35.525 28.395 -35.195 28.725 ;
        RECT -35.525 27.035 -35.195 27.365 ;
        RECT -35.525 25.675 -35.195 26.005 ;
        RECT -35.525 24.315 -35.195 24.645 ;
        RECT -35.525 22.955 -35.195 23.285 ;
        RECT -35.525 21.595 -35.195 21.925 ;
        RECT -35.525 20.235 -35.195 20.565 ;
        RECT -35.525 18.875 -35.195 19.205 ;
        RECT -35.525 17.515 -35.195 17.845 ;
        RECT -35.525 16.155 -35.195 16.485 ;
        RECT -35.525 14.795 -35.195 15.125 ;
        RECT -35.525 13.435 -35.195 13.765 ;
        RECT -35.525 12.075 -35.195 12.405 ;
        RECT -35.525 10.715 -35.195 11.045 ;
        RECT -35.525 9.355 -35.195 9.685 ;
        RECT -35.525 7.995 -35.195 8.325 ;
        RECT -35.525 6.635 -35.195 6.965 ;
        RECT -35.525 5.275 -35.195 5.605 ;
        RECT -35.525 3.915 -35.195 4.245 ;
        RECT -35.525 2.555 -35.195 2.885 ;
        RECT -35.525 1.195 -35.195 1.525 ;
        RECT -35.525 -0.165 -35.195 0.165 ;
        RECT -35.525 -8.325 -35.195 -7.995 ;
        RECT -35.525 -11.045 -35.195 -10.715 ;
        RECT -35.525 -15.125 -35.195 -14.795 ;
        RECT -35.525 -16.485 -35.195 -16.155 ;
        RECT -35.525 -17.845 -35.195 -17.515 ;
        RECT -35.525 -19.205 -35.195 -18.875 ;
        RECT -35.525 -20.565 -35.195 -20.235 ;
        RECT -35.525 -21.925 -35.195 -21.595 ;
        RECT -35.525 -23.285 -35.195 -22.955 ;
        RECT -35.525 -24.645 -35.195 -24.315 ;
        RECT -35.525 -31.445 -35.195 -31.115 ;
        RECT -35.525 -32.805 -35.195 -32.475 ;
        RECT -35.525 -35.525 -35.195 -35.195 ;
        RECT -35.525 -36.885 -35.195 -36.555 ;
        RECT -35.525 -37.93 -35.195 -37.6 ;
        RECT -35.525 -40.965 -35.195 -40.635 ;
        RECT -35.525 -42.77 -35.195 -42.44 ;
        RECT -35.525 -43.685 -35.195 -43.355 ;
        RECT -35.525 -50.485 -35.195 -50.155 ;
        RECT -35.525 -51.845 -35.195 -51.515 ;
        RECT -35.525 -53.205 -35.195 -52.875 ;
        RECT -35.525 -54.565 -35.195 -54.235 ;
        RECT -35.525 -55.925 -35.195 -55.595 ;
        RECT -35.525 -57.285 -35.195 -56.955 ;
        RECT -35.525 -58.645 -35.195 -58.315 ;
        RECT -35.525 -60.005 -35.195 -59.675 ;
        RECT -35.525 -61.365 -35.195 -61.035 ;
        RECT -35.525 -64.085 -35.195 -63.755 ;
        RECT -35.525 -65.445 -35.195 -65.115 ;
        RECT -35.525 -66.805 -35.195 -66.475 ;
        RECT -35.525 -68.165 -35.195 -67.835 ;
        RECT -35.525 -69.525 -35.195 -69.195 ;
        RECT -35.525 -70.885 -35.195 -70.555 ;
        RECT -35.525 -72.245 -35.195 -71.915 ;
        RECT -35.525 -73.605 -35.195 -73.275 ;
        RECT -35.525 -74.965 -35.195 -74.635 ;
        RECT -35.525 -76.325 -35.195 -75.995 ;
        RECT -35.525 -77.685 -35.195 -77.355 ;
        RECT -35.525 -79.045 -35.195 -78.715 ;
        RECT -35.525 -80.405 -35.195 -80.075 ;
        RECT -35.525 -81.765 -35.195 -81.435 ;
        RECT -35.525 -83.125 -35.195 -82.795 ;
        RECT -35.525 -84.485 -35.195 -84.155 ;
        RECT -35.525 -85.845 -35.195 -85.515 ;
        RECT -35.525 -87.205 -35.195 -86.875 ;
        RECT -35.525 -88.565 -35.195 -88.235 ;
        RECT -35.525 -89.925 -35.195 -89.595 ;
        RECT -35.525 -92.645 -35.195 -92.315 ;
        RECT -35.525 -94.005 -35.195 -93.675 ;
        RECT -35.525 -95.365 -35.195 -95.035 ;
        RECT -35.525 -96.725 -35.195 -96.395 ;
        RECT -35.525 -98.73 -35.195 -98.4 ;
        RECT -35.525 -99.445 -35.195 -99.115 ;
        RECT -35.525 -102.165 -35.195 -101.835 ;
        RECT -35.525 -103.525 -35.195 -103.195 ;
        RECT -35.525 -104.885 -35.195 -104.555 ;
        RECT -35.525 -106.87 -35.195 -106.54 ;
        RECT -35.525 -107.605 -35.195 -107.275 ;
        RECT -35.525 -108.965 -35.195 -108.635 ;
        RECT -35.52 -111.68 -35.2 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -35.525 -174.245 -35.195 -173.915 ;
        RECT -35.525 -175.725 -35.195 -175.395 ;
        RECT -35.525 -176.965 -35.195 -176.635 ;
        RECT -35.525 -178.325 -35.195 -177.995 ;
        RECT -35.525 -180.57 -35.195 -179.44 ;
        RECT -35.52 -180.685 -35.2 -172.56 ;
    END
    PORT
      LAYER met3 ;
        RECT -34.165 -77.685 -33.835 -77.355 ;
        RECT -34.165 -79.045 -33.835 -78.715 ;
        RECT -34.165 -80.405 -33.835 -80.075 ;
        RECT -34.165 -81.765 -33.835 -81.435 ;
        RECT -34.165 -83.125 -33.835 -82.795 ;
        RECT -34.165 -84.485 -33.835 -84.155 ;
        RECT -34.165 -85.845 -33.835 -85.515 ;
        RECT -34.165 -87.205 -33.835 -86.875 ;
        RECT -34.165 -88.565 -33.835 -88.235 ;
        RECT -34.165 -89.925 -33.835 -89.595 ;
        RECT -34.165 -92.645 -33.835 -92.315 ;
        RECT -34.165 -94.005 -33.835 -93.675 ;
        RECT -34.165 -95.365 -33.835 -95.035 ;
        RECT -34.165 -96.725 -33.835 -96.395 ;
        RECT -34.165 -98.73 -33.835 -98.4 ;
        RECT -34.165 -99.445 -33.835 -99.115 ;
        RECT -34.165 -102.165 -33.835 -101.835 ;
        RECT -34.165 -103.525 -33.835 -103.195 ;
        RECT -34.165 -104.885 -33.835 -104.555 ;
        RECT -34.165 -106.87 -33.835 -106.54 ;
        RECT -34.165 -107.605 -33.835 -107.275 ;
        RECT -34.165 -108.965 -33.835 -108.635 ;
        RECT -34.165 -114.405 -33.835 -114.075 ;
        RECT -34.165 -115.765 -33.835 -115.435 ;
        RECT -34.165 -117.125 -33.835 -116.795 ;
        RECT -34.165 -118.485 -33.835 -118.155 ;
        RECT -34.165 -122.565 -33.835 -122.235 ;
        RECT -34.165 -125.285 -33.835 -124.955 ;
        RECT -34.165 -126.645 -33.835 -126.315 ;
        RECT -34.165 -128.005 -33.835 -127.675 ;
        RECT -34.165 -129.365 -33.835 -129.035 ;
        RECT -34.165 -133.445 -33.835 -133.115 ;
        RECT -34.165 -134.805 -33.835 -134.475 ;
        RECT -34.165 -136.165 -33.835 -135.835 ;
        RECT -34.165 -137.525 -33.835 -137.195 ;
        RECT -34.165 -138.885 -33.835 -138.555 ;
        RECT -34.165 -141.605 -33.835 -141.275 ;
        RECT -34.165 -142.965 -33.835 -142.635 ;
        RECT -34.165 -144.325 -33.835 -143.995 ;
        RECT -34.165 -145.685 -33.835 -145.355 ;
        RECT -34.165 -147.045 -33.835 -146.715 ;
        RECT -34.165 -148.405 -33.835 -148.075 ;
        RECT -34.165 -151.125 -33.835 -150.795 ;
        RECT -34.165 -152.485 -33.835 -152.155 ;
        RECT -34.165 -156.565 -33.835 -156.235 ;
        RECT -34.165 -157.925 -33.835 -157.595 ;
        RECT -34.165 -159.285 -33.835 -158.955 ;
        RECT -34.165 -160.645 -33.835 -160.315 ;
        RECT -34.165 -162.005 -33.835 -161.675 ;
        RECT -34.165 -163.365 -33.835 -163.035 ;
        RECT -34.165 -164.725 -33.835 -164.395 ;
        RECT -34.165 -166.085 -33.835 -165.755 ;
        RECT -34.165 -167.445 -33.835 -167.115 ;
        RECT -34.165 -170.165 -33.835 -169.835 ;
        RECT -34.16 -172.2 -33.84 242.565 ;
        RECT -34.165 241.32 -33.835 242.45 ;
        RECT -34.165 239.195 -33.835 239.525 ;
        RECT -34.165 237.835 -33.835 238.165 ;
        RECT -34.165 236.475 -33.835 236.805 ;
        RECT -34.165 235.115 -33.835 235.445 ;
        RECT -34.165 233.755 -33.835 234.085 ;
        RECT -34.165 232.395 -33.835 232.725 ;
        RECT -34.165 231.035 -33.835 231.365 ;
        RECT -34.165 229.675 -33.835 230.005 ;
        RECT -34.165 228.315 -33.835 228.645 ;
        RECT -34.165 226.955 -33.835 227.285 ;
        RECT -34.165 225.595 -33.835 225.925 ;
        RECT -34.165 224.235 -33.835 224.565 ;
        RECT -34.165 222.875 -33.835 223.205 ;
        RECT -34.165 221.515 -33.835 221.845 ;
        RECT -34.165 220.155 -33.835 220.485 ;
        RECT -34.165 218.795 -33.835 219.125 ;
        RECT -34.165 217.435 -33.835 217.765 ;
        RECT -34.165 216.075 -33.835 216.405 ;
        RECT -34.165 214.715 -33.835 215.045 ;
        RECT -34.165 213.355 -33.835 213.685 ;
        RECT -34.165 211.995 -33.835 212.325 ;
        RECT -34.165 210.635 -33.835 210.965 ;
        RECT -34.165 209.275 -33.835 209.605 ;
        RECT -34.165 207.915 -33.835 208.245 ;
        RECT -34.165 206.555 -33.835 206.885 ;
        RECT -34.165 205.195 -33.835 205.525 ;
        RECT -34.165 203.835 -33.835 204.165 ;
        RECT -34.165 202.475 -33.835 202.805 ;
        RECT -34.165 201.115 -33.835 201.445 ;
        RECT -34.165 199.755 -33.835 200.085 ;
        RECT -34.165 198.395 -33.835 198.725 ;
        RECT -34.165 197.035 -33.835 197.365 ;
        RECT -34.165 195.675 -33.835 196.005 ;
        RECT -34.165 194.315 -33.835 194.645 ;
        RECT -34.165 192.955 -33.835 193.285 ;
        RECT -34.165 191.595 -33.835 191.925 ;
        RECT -34.165 190.235 -33.835 190.565 ;
        RECT -34.165 188.875 -33.835 189.205 ;
        RECT -34.165 187.515 -33.835 187.845 ;
        RECT -34.165 186.155 -33.835 186.485 ;
        RECT -34.165 184.795 -33.835 185.125 ;
        RECT -34.165 183.435 -33.835 183.765 ;
        RECT -34.165 182.075 -33.835 182.405 ;
        RECT -34.165 180.715 -33.835 181.045 ;
        RECT -34.165 179.355 -33.835 179.685 ;
        RECT -34.165 177.995 -33.835 178.325 ;
        RECT -34.165 176.635 -33.835 176.965 ;
        RECT -34.165 175.275 -33.835 175.605 ;
        RECT -34.165 173.915 -33.835 174.245 ;
        RECT -34.165 172.555 -33.835 172.885 ;
        RECT -34.165 171.195 -33.835 171.525 ;
        RECT -34.165 169.835 -33.835 170.165 ;
        RECT -34.165 168.475 -33.835 168.805 ;
        RECT -34.165 167.115 -33.835 167.445 ;
        RECT -34.165 165.755 -33.835 166.085 ;
        RECT -34.165 164.395 -33.835 164.725 ;
        RECT -34.165 163.035 -33.835 163.365 ;
        RECT -34.165 161.675 -33.835 162.005 ;
        RECT -34.165 160.315 -33.835 160.645 ;
        RECT -34.165 158.955 -33.835 159.285 ;
        RECT -34.165 157.595 -33.835 157.925 ;
        RECT -34.165 156.235 -33.835 156.565 ;
        RECT -34.165 154.875 -33.835 155.205 ;
        RECT -34.165 153.515 -33.835 153.845 ;
        RECT -34.165 152.155 -33.835 152.485 ;
        RECT -34.165 150.795 -33.835 151.125 ;
        RECT -34.165 149.435 -33.835 149.765 ;
        RECT -34.165 148.075 -33.835 148.405 ;
        RECT -34.165 146.715 -33.835 147.045 ;
        RECT -34.165 145.355 -33.835 145.685 ;
        RECT -34.165 143.995 -33.835 144.325 ;
        RECT -34.165 142.635 -33.835 142.965 ;
        RECT -34.165 141.275 -33.835 141.605 ;
        RECT -34.165 139.915 -33.835 140.245 ;
        RECT -34.165 138.555 -33.835 138.885 ;
        RECT -34.165 137.195 -33.835 137.525 ;
        RECT -34.165 135.835 -33.835 136.165 ;
        RECT -34.165 134.475 -33.835 134.805 ;
        RECT -34.165 133.115 -33.835 133.445 ;
        RECT -34.165 131.755 -33.835 132.085 ;
        RECT -34.165 130.395 -33.835 130.725 ;
        RECT -34.165 129.035 -33.835 129.365 ;
        RECT -34.165 127.675 -33.835 128.005 ;
        RECT -34.165 126.315 -33.835 126.645 ;
        RECT -34.165 124.955 -33.835 125.285 ;
        RECT -34.165 123.595 -33.835 123.925 ;
        RECT -34.165 122.235 -33.835 122.565 ;
        RECT -34.165 120.875 -33.835 121.205 ;
        RECT -34.165 119.515 -33.835 119.845 ;
        RECT -34.165 118.155 -33.835 118.485 ;
        RECT -34.165 116.795 -33.835 117.125 ;
        RECT -34.165 115.435 -33.835 115.765 ;
        RECT -34.165 114.075 -33.835 114.405 ;
        RECT -34.165 112.715 -33.835 113.045 ;
        RECT -34.165 111.355 -33.835 111.685 ;
        RECT -34.165 109.995 -33.835 110.325 ;
        RECT -34.165 108.635 -33.835 108.965 ;
        RECT -34.165 107.275 -33.835 107.605 ;
        RECT -34.165 105.915 -33.835 106.245 ;
        RECT -34.165 104.555 -33.835 104.885 ;
        RECT -34.165 103.195 -33.835 103.525 ;
        RECT -34.165 101.835 -33.835 102.165 ;
        RECT -34.165 100.475 -33.835 100.805 ;
        RECT -34.165 99.115 -33.835 99.445 ;
        RECT -34.165 97.755 -33.835 98.085 ;
        RECT -34.165 96.395 -33.835 96.725 ;
        RECT -34.165 95.035 -33.835 95.365 ;
        RECT -34.165 93.675 -33.835 94.005 ;
        RECT -34.165 92.315 -33.835 92.645 ;
        RECT -34.165 90.955 -33.835 91.285 ;
        RECT -34.165 89.595 -33.835 89.925 ;
        RECT -34.165 88.235 -33.835 88.565 ;
        RECT -34.165 86.875 -33.835 87.205 ;
        RECT -34.165 85.515 -33.835 85.845 ;
        RECT -34.165 84.155 -33.835 84.485 ;
        RECT -34.165 82.795 -33.835 83.125 ;
        RECT -34.165 81.435 -33.835 81.765 ;
        RECT -34.165 80.075 -33.835 80.405 ;
        RECT -34.165 78.715 -33.835 79.045 ;
        RECT -34.165 77.355 -33.835 77.685 ;
        RECT -34.165 75.995 -33.835 76.325 ;
        RECT -34.165 74.635 -33.835 74.965 ;
        RECT -34.165 73.275 -33.835 73.605 ;
        RECT -34.165 71.915 -33.835 72.245 ;
        RECT -34.165 70.555 -33.835 70.885 ;
        RECT -34.165 69.195 -33.835 69.525 ;
        RECT -34.165 67.835 -33.835 68.165 ;
        RECT -34.165 66.475 -33.835 66.805 ;
        RECT -34.165 65.115 -33.835 65.445 ;
        RECT -34.165 63.755 -33.835 64.085 ;
        RECT -34.165 62.395 -33.835 62.725 ;
        RECT -34.165 61.035 -33.835 61.365 ;
        RECT -34.165 59.675 -33.835 60.005 ;
        RECT -34.165 58.315 -33.835 58.645 ;
        RECT -34.165 56.955 -33.835 57.285 ;
        RECT -34.165 55.595 -33.835 55.925 ;
        RECT -34.165 54.235 -33.835 54.565 ;
        RECT -34.165 52.875 -33.835 53.205 ;
        RECT -34.165 51.515 -33.835 51.845 ;
        RECT -34.165 50.155 -33.835 50.485 ;
        RECT -34.165 48.795 -33.835 49.125 ;
        RECT -34.165 47.435 -33.835 47.765 ;
        RECT -34.165 46.075 -33.835 46.405 ;
        RECT -34.165 44.715 -33.835 45.045 ;
        RECT -34.165 43.355 -33.835 43.685 ;
        RECT -34.165 41.995 -33.835 42.325 ;
        RECT -34.165 40.635 -33.835 40.965 ;
        RECT -34.165 39.275 -33.835 39.605 ;
        RECT -34.165 37.915 -33.835 38.245 ;
        RECT -34.165 36.555 -33.835 36.885 ;
        RECT -34.165 35.195 -33.835 35.525 ;
        RECT -34.165 33.835 -33.835 34.165 ;
        RECT -34.165 32.475 -33.835 32.805 ;
        RECT -34.165 31.115 -33.835 31.445 ;
        RECT -34.165 29.755 -33.835 30.085 ;
        RECT -34.165 28.395 -33.835 28.725 ;
        RECT -34.165 27.035 -33.835 27.365 ;
        RECT -34.165 25.675 -33.835 26.005 ;
        RECT -34.165 24.315 -33.835 24.645 ;
        RECT -34.165 22.955 -33.835 23.285 ;
        RECT -34.165 21.595 -33.835 21.925 ;
        RECT -34.165 20.235 -33.835 20.565 ;
        RECT -34.165 18.875 -33.835 19.205 ;
        RECT -34.165 17.515 -33.835 17.845 ;
        RECT -34.165 16.155 -33.835 16.485 ;
        RECT -34.165 14.795 -33.835 15.125 ;
        RECT -34.165 13.435 -33.835 13.765 ;
        RECT -34.165 12.075 -33.835 12.405 ;
        RECT -34.165 10.715 -33.835 11.045 ;
        RECT -34.165 9.355 -33.835 9.685 ;
        RECT -34.165 7.995 -33.835 8.325 ;
        RECT -34.165 6.635 -33.835 6.965 ;
        RECT -34.165 5.275 -33.835 5.605 ;
        RECT -34.165 3.915 -33.835 4.245 ;
        RECT -34.165 2.555 -33.835 2.885 ;
        RECT -34.165 1.195 -33.835 1.525 ;
        RECT -34.165 -0.165 -33.835 0.165 ;
        RECT -34.165 -8.325 -33.835 -7.995 ;
        RECT -34.165 -11.045 -33.835 -10.715 ;
        RECT -34.165 -15.125 -33.835 -14.795 ;
        RECT -34.165 -16.485 -33.835 -16.155 ;
        RECT -34.165 -17.845 -33.835 -17.515 ;
        RECT -34.165 -19.205 -33.835 -18.875 ;
        RECT -34.165 -20.565 -33.835 -20.235 ;
        RECT -34.165 -21.925 -33.835 -21.595 ;
        RECT -34.165 -23.285 -33.835 -22.955 ;
        RECT -34.165 -24.645 -33.835 -24.315 ;
        RECT -34.165 -31.445 -33.835 -31.115 ;
        RECT -34.165 -32.805 -33.835 -32.475 ;
        RECT -34.165 -35.525 -33.835 -35.195 ;
        RECT -34.165 -36.885 -33.835 -36.555 ;
        RECT -34.165 -37.93 -33.835 -37.6 ;
        RECT -34.165 -40.965 -33.835 -40.635 ;
        RECT -34.165 -42.77 -33.835 -42.44 ;
        RECT -34.165 -43.685 -33.835 -43.355 ;
        RECT -34.165 -50.485 -33.835 -50.155 ;
        RECT -34.165 -51.845 -33.835 -51.515 ;
        RECT -34.165 -54.565 -33.835 -54.235 ;
        RECT -34.165 -55.925 -33.835 -55.595 ;
        RECT -34.165 -60.005 -33.835 -59.675 ;
        RECT -34.165 -68.165 -33.835 -67.835 ;
        RECT -34.165 -69.525 -33.835 -69.195 ;
        RECT -34.165 -70.885 -33.835 -70.555 ;
        RECT -34.165 -72.245 -33.835 -71.915 ;
        RECT -34.165 -73.605 -33.835 -73.275 ;
        RECT -34.165 -74.965 -33.835 -74.635 ;
        RECT -34.165 -76.325 -33.835 -75.995 ;
    END
    PORT
      LAYER met3 ;
        RECT -45.045 -69.525 -44.715 -69.195 ;
        RECT -45.045 -70.885 -44.715 -70.555 ;
        RECT -45.045 -72.245 -44.715 -71.915 ;
        RECT -45.045 -73.605 -44.715 -73.275 ;
        RECT -45.045 -74.965 -44.715 -74.635 ;
        RECT -45.045 -76.325 -44.715 -75.995 ;
        RECT -45.045 -77.685 -44.715 -77.355 ;
        RECT -45.045 -79.045 -44.715 -78.715 ;
        RECT -45.045 -80.405 -44.715 -80.075 ;
        RECT -45.045 -81.765 -44.715 -81.435 ;
        RECT -45.045 -83.125 -44.715 -82.795 ;
        RECT -45.045 -84.485 -44.715 -84.155 ;
        RECT -45.045 -85.845 -44.715 -85.515 ;
        RECT -45.045 -87.205 -44.715 -86.875 ;
        RECT -45.045 -88.565 -44.715 -88.235 ;
        RECT -45.045 -89.925 -44.715 -89.595 ;
        RECT -45.045 -92.645 -44.715 -92.315 ;
        RECT -45.045 -94.005 -44.715 -93.675 ;
        RECT -45.045 -95.365 -44.715 -95.035 ;
        RECT -45.045 -96.725 -44.715 -96.395 ;
        RECT -45.045 -98.73 -44.715 -98.4 ;
        RECT -45.045 -99.445 -44.715 -99.115 ;
        RECT -45.045 -102.165 -44.715 -101.835 ;
        RECT -45.045 -103.525 -44.715 -103.195 ;
        RECT -45.045 -104.885 -44.715 -104.555 ;
        RECT -45.045 -106.87 -44.715 -106.54 ;
        RECT -45.045 -107.605 -44.715 -107.275 ;
        RECT -45.045 -108.965 -44.715 -108.635 ;
        RECT -45.045 -113.045 -44.715 -112.715 ;
        RECT -45.045 -114.405 -44.715 -114.075 ;
        RECT -45.045 -115.765 -44.715 -115.435 ;
        RECT -45.045 -117.125 -44.715 -116.795 ;
        RECT -45.045 -118.485 -44.715 -118.155 ;
        RECT -45.045 -122.565 -44.715 -122.235 ;
        RECT -45.045 -123.925 -44.715 -123.595 ;
        RECT -45.045 -125.285 -44.715 -124.955 ;
        RECT -45.045 -126.645 -44.715 -126.315 ;
        RECT -45.045 -128.005 -44.715 -127.675 ;
        RECT -45.045 -129.365 -44.715 -129.035 ;
        RECT -45.045 -130.725 -44.715 -130.395 ;
        RECT -45.045 -132.085 -44.715 -131.755 ;
        RECT -45.045 -133.445 -44.715 -133.115 ;
        RECT -45.045 -134.805 -44.715 -134.475 ;
        RECT -45.045 -136.165 -44.715 -135.835 ;
        RECT -45.045 -137.525 -44.715 -137.195 ;
        RECT -45.045 -138.885 -44.715 -138.555 ;
        RECT -45.045 -140.245 -44.715 -139.915 ;
        RECT -45.045 -141.605 -44.715 -141.275 ;
        RECT -45.045 -142.965 -44.715 -142.635 ;
        RECT -45.045 -144.325 -44.715 -143.995 ;
        RECT -45.045 -145.685 -44.715 -145.355 ;
        RECT -45.045 -147.045 -44.715 -146.715 ;
        RECT -45.045 -148.405 -44.715 -148.075 ;
        RECT -45.045 -149.765 -44.715 -149.435 ;
        RECT -45.045 -151.125 -44.715 -150.795 ;
        RECT -45.045 -152.485 -44.715 -152.155 ;
        RECT -45.045 -153.845 -44.715 -153.515 ;
        RECT -45.045 -155.205 -44.715 -154.875 ;
        RECT -45.045 -156.565 -44.715 -156.235 ;
        RECT -45.045 -157.925 -44.715 -157.595 ;
        RECT -45.045 -159.285 -44.715 -158.955 ;
        RECT -45.045 -160.645 -44.715 -160.315 ;
        RECT -45.045 -162.005 -44.715 -161.675 ;
        RECT -45.045 -163.365 -44.715 -163.035 ;
        RECT -45.045 -164.725 -44.715 -164.395 ;
        RECT -45.045 -166.085 -44.715 -165.755 ;
        RECT -45.045 -167.445 -44.715 -167.115 ;
        RECT -45.045 -170.165 -44.715 -169.835 ;
        RECT -45.045 -172.885 -44.715 -172.555 ;
        RECT -45.045 -174.245 -44.715 -173.915 ;
        RECT -45.045 -175.725 -44.715 -175.395 ;
        RECT -45.045 -176.965 -44.715 -176.635 ;
        RECT -45.045 -178.325 -44.715 -177.995 ;
        RECT -45.045 -180.57 -44.715 -179.44 ;
        RECT -45.04 -180.685 -44.72 -69.195 ;
    END
    PORT
      LAYER met3 ;
        RECT -43.685 241.32 -43.355 242.45 ;
        RECT -43.685 239.195 -43.355 239.525 ;
        RECT -43.685 237.835 -43.355 238.165 ;
        RECT -43.685 236.475 -43.355 236.805 ;
        RECT -43.685 235.115 -43.355 235.445 ;
        RECT -43.685 233.755 -43.355 234.085 ;
        RECT -43.685 232.395 -43.355 232.725 ;
        RECT -43.685 231.035 -43.355 231.365 ;
        RECT -43.685 229.675 -43.355 230.005 ;
        RECT -43.685 228.315 -43.355 228.645 ;
        RECT -43.685 226.955 -43.355 227.285 ;
        RECT -43.685 225.595 -43.355 225.925 ;
        RECT -43.685 224.235 -43.355 224.565 ;
        RECT -43.685 222.875 -43.355 223.205 ;
        RECT -43.685 221.515 -43.355 221.845 ;
        RECT -43.685 220.155 -43.355 220.485 ;
        RECT -43.685 218.795 -43.355 219.125 ;
        RECT -43.685 217.435 -43.355 217.765 ;
        RECT -43.685 216.075 -43.355 216.405 ;
        RECT -43.685 214.715 -43.355 215.045 ;
        RECT -43.685 213.355 -43.355 213.685 ;
        RECT -43.685 211.995 -43.355 212.325 ;
        RECT -43.685 210.635 -43.355 210.965 ;
        RECT -43.685 209.275 -43.355 209.605 ;
        RECT -43.685 207.915 -43.355 208.245 ;
        RECT -43.685 206.555 -43.355 206.885 ;
        RECT -43.685 205.195 -43.355 205.525 ;
        RECT -43.685 203.835 -43.355 204.165 ;
        RECT -43.685 202.475 -43.355 202.805 ;
        RECT -43.685 201.115 -43.355 201.445 ;
        RECT -43.685 199.755 -43.355 200.085 ;
        RECT -43.685 198.395 -43.355 198.725 ;
        RECT -43.685 197.035 -43.355 197.365 ;
        RECT -43.685 195.675 -43.355 196.005 ;
        RECT -43.685 194.315 -43.355 194.645 ;
        RECT -43.685 192.955 -43.355 193.285 ;
        RECT -43.685 191.595 -43.355 191.925 ;
        RECT -43.685 190.235 -43.355 190.565 ;
        RECT -43.685 188.875 -43.355 189.205 ;
        RECT -43.685 187.515 -43.355 187.845 ;
        RECT -43.685 186.155 -43.355 186.485 ;
        RECT -43.685 184.795 -43.355 185.125 ;
        RECT -43.685 183.435 -43.355 183.765 ;
        RECT -43.685 182.075 -43.355 182.405 ;
        RECT -43.685 180.715 -43.355 181.045 ;
        RECT -43.685 179.355 -43.355 179.685 ;
        RECT -43.685 177.995 -43.355 178.325 ;
        RECT -43.685 176.635 -43.355 176.965 ;
        RECT -43.685 175.275 -43.355 175.605 ;
        RECT -43.685 173.915 -43.355 174.245 ;
        RECT -43.685 172.555 -43.355 172.885 ;
        RECT -43.685 171.195 -43.355 171.525 ;
        RECT -43.685 169.835 -43.355 170.165 ;
        RECT -43.685 168.475 -43.355 168.805 ;
        RECT -43.685 167.115 -43.355 167.445 ;
        RECT -43.685 165.755 -43.355 166.085 ;
        RECT -43.685 164.395 -43.355 164.725 ;
        RECT -43.685 163.035 -43.355 163.365 ;
        RECT -43.685 161.675 -43.355 162.005 ;
        RECT -43.685 160.315 -43.355 160.645 ;
        RECT -43.685 158.955 -43.355 159.285 ;
        RECT -43.685 157.595 -43.355 157.925 ;
        RECT -43.685 156.235 -43.355 156.565 ;
        RECT -43.685 154.875 -43.355 155.205 ;
        RECT -43.685 153.515 -43.355 153.845 ;
        RECT -43.685 152.155 -43.355 152.485 ;
        RECT -43.685 150.795 -43.355 151.125 ;
        RECT -43.685 149.435 -43.355 149.765 ;
        RECT -43.685 148.075 -43.355 148.405 ;
        RECT -43.685 146.715 -43.355 147.045 ;
        RECT -43.685 145.355 -43.355 145.685 ;
        RECT -43.685 143.995 -43.355 144.325 ;
        RECT -43.685 142.635 -43.355 142.965 ;
        RECT -43.685 141.275 -43.355 141.605 ;
        RECT -43.685 139.915 -43.355 140.245 ;
        RECT -43.685 138.555 -43.355 138.885 ;
        RECT -43.685 137.195 -43.355 137.525 ;
        RECT -43.685 135.835 -43.355 136.165 ;
        RECT -43.685 134.475 -43.355 134.805 ;
        RECT -43.685 133.115 -43.355 133.445 ;
        RECT -43.685 131.755 -43.355 132.085 ;
        RECT -43.685 130.395 -43.355 130.725 ;
        RECT -43.685 129.035 -43.355 129.365 ;
        RECT -43.685 127.675 -43.355 128.005 ;
        RECT -43.685 126.315 -43.355 126.645 ;
        RECT -43.685 124.955 -43.355 125.285 ;
        RECT -43.685 123.595 -43.355 123.925 ;
        RECT -43.685 122.235 -43.355 122.565 ;
        RECT -43.685 120.875 -43.355 121.205 ;
        RECT -43.685 119.515 -43.355 119.845 ;
        RECT -43.685 118.155 -43.355 118.485 ;
        RECT -43.685 116.795 -43.355 117.125 ;
        RECT -43.685 115.435 -43.355 115.765 ;
        RECT -43.685 114.075 -43.355 114.405 ;
        RECT -43.685 112.715 -43.355 113.045 ;
        RECT -43.685 111.355 -43.355 111.685 ;
        RECT -43.685 109.995 -43.355 110.325 ;
        RECT -43.685 108.635 -43.355 108.965 ;
        RECT -43.685 107.275 -43.355 107.605 ;
        RECT -43.685 105.915 -43.355 106.245 ;
        RECT -43.685 104.555 -43.355 104.885 ;
        RECT -43.685 103.195 -43.355 103.525 ;
        RECT -43.685 101.835 -43.355 102.165 ;
        RECT -43.685 100.475 -43.355 100.805 ;
        RECT -43.685 99.115 -43.355 99.445 ;
        RECT -43.685 97.755 -43.355 98.085 ;
        RECT -43.685 96.395 -43.355 96.725 ;
        RECT -43.685 95.035 -43.355 95.365 ;
        RECT -43.685 93.675 -43.355 94.005 ;
        RECT -43.685 92.315 -43.355 92.645 ;
        RECT -43.685 90.955 -43.355 91.285 ;
        RECT -43.685 89.595 -43.355 89.925 ;
        RECT -43.685 88.235 -43.355 88.565 ;
        RECT -43.685 86.875 -43.355 87.205 ;
        RECT -43.685 85.515 -43.355 85.845 ;
        RECT -43.685 84.155 -43.355 84.485 ;
        RECT -43.685 82.795 -43.355 83.125 ;
        RECT -43.685 81.435 -43.355 81.765 ;
        RECT -43.685 80.075 -43.355 80.405 ;
        RECT -43.685 78.715 -43.355 79.045 ;
        RECT -43.685 77.355 -43.355 77.685 ;
        RECT -43.685 75.995 -43.355 76.325 ;
        RECT -43.685 74.635 -43.355 74.965 ;
        RECT -43.685 73.275 -43.355 73.605 ;
        RECT -43.685 71.915 -43.355 72.245 ;
        RECT -43.685 70.555 -43.355 70.885 ;
        RECT -43.685 69.195 -43.355 69.525 ;
        RECT -43.685 67.835 -43.355 68.165 ;
        RECT -43.685 66.475 -43.355 66.805 ;
        RECT -43.685 65.115 -43.355 65.445 ;
        RECT -43.685 63.755 -43.355 64.085 ;
        RECT -43.685 62.395 -43.355 62.725 ;
        RECT -43.685 61.035 -43.355 61.365 ;
        RECT -43.685 59.675 -43.355 60.005 ;
        RECT -43.685 58.315 -43.355 58.645 ;
        RECT -43.685 56.955 -43.355 57.285 ;
        RECT -43.685 55.595 -43.355 55.925 ;
        RECT -43.685 54.235 -43.355 54.565 ;
        RECT -43.685 52.875 -43.355 53.205 ;
        RECT -43.685 51.515 -43.355 51.845 ;
        RECT -43.685 50.155 -43.355 50.485 ;
        RECT -43.685 48.795 -43.355 49.125 ;
        RECT -43.685 47.435 -43.355 47.765 ;
        RECT -43.685 46.075 -43.355 46.405 ;
        RECT -43.685 44.715 -43.355 45.045 ;
        RECT -43.685 43.355 -43.355 43.685 ;
        RECT -43.685 41.995 -43.355 42.325 ;
        RECT -43.685 40.635 -43.355 40.965 ;
        RECT -43.685 39.275 -43.355 39.605 ;
        RECT -43.685 37.915 -43.355 38.245 ;
        RECT -43.685 36.555 -43.355 36.885 ;
        RECT -43.685 35.195 -43.355 35.525 ;
        RECT -43.685 33.835 -43.355 34.165 ;
        RECT -43.685 32.475 -43.355 32.805 ;
        RECT -43.685 31.115 -43.355 31.445 ;
        RECT -43.685 29.755 -43.355 30.085 ;
        RECT -43.685 28.395 -43.355 28.725 ;
        RECT -43.685 27.035 -43.355 27.365 ;
        RECT -43.685 25.675 -43.355 26.005 ;
        RECT -43.685 24.315 -43.355 24.645 ;
        RECT -43.685 22.955 -43.355 23.285 ;
        RECT -43.685 21.595 -43.355 21.925 ;
        RECT -43.685 20.235 -43.355 20.565 ;
        RECT -43.685 18.875 -43.355 19.205 ;
        RECT -43.685 17.515 -43.355 17.845 ;
        RECT -43.685 16.155 -43.355 16.485 ;
        RECT -43.685 14.795 -43.355 15.125 ;
        RECT -43.685 13.435 -43.355 13.765 ;
        RECT -43.685 12.075 -43.355 12.405 ;
        RECT -43.685 10.715 -43.355 11.045 ;
        RECT -43.685 9.355 -43.355 9.685 ;
        RECT -43.685 7.995 -43.355 8.325 ;
        RECT -43.685 6.635 -43.355 6.965 ;
        RECT -43.685 5.275 -43.355 5.605 ;
        RECT -43.685 3.915 -43.355 4.245 ;
        RECT -43.685 2.555 -43.355 2.885 ;
        RECT -43.685 1.195 -43.355 1.525 ;
        RECT -43.685 -0.165 -43.355 0.165 ;
        RECT -43.685 -4.245 -43.355 -3.915 ;
        RECT -43.685 -5.605 -43.355 -5.275 ;
        RECT -43.685 -6.965 -43.355 -6.635 ;
        RECT -43.685 -11.045 -43.355 -10.715 ;
        RECT -43.685 -15.125 -43.355 -14.795 ;
        RECT -43.685 -16.485 -43.355 -16.155 ;
        RECT -43.685 -17.845 -43.355 -17.515 ;
        RECT -43.685 -19.205 -43.355 -18.875 ;
        RECT -43.685 -20.565 -43.355 -20.235 ;
        RECT -43.685 -21.925 -43.355 -21.595 ;
        RECT -43.685 -23.285 -43.355 -22.955 ;
        RECT -43.685 -24.645 -43.355 -24.315 ;
        RECT -43.685 -31.445 -43.355 -31.115 ;
        RECT -43.685 -32.805 -43.355 -32.475 ;
        RECT -43.685 -35.525 -43.355 -35.195 ;
        RECT -43.685 -36.885 -43.355 -36.555 ;
        RECT -43.685 -37.93 -43.355 -37.6 ;
        RECT -43.685 -40.965 -43.355 -40.635 ;
        RECT -43.685 -42.77 -43.355 -42.44 ;
        RECT -43.685 -43.685 -43.355 -43.355 ;
        RECT -43.685 -50.485 -43.355 -50.155 ;
        RECT -43.685 -51.845 -43.355 -51.515 ;
        RECT -43.685 -54.565 -43.355 -54.235 ;
        RECT -43.685 -55.925 -43.355 -55.595 ;
        RECT -43.685 -60.005 -43.355 -59.675 ;
        RECT -43.68 -64.08 -43.36 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -43.685 -69.525 -43.355 -69.195 ;
        RECT -43.685 -70.885 -43.355 -70.555 ;
        RECT -43.685 -72.245 -43.355 -71.915 ;
        RECT -43.685 -73.605 -43.355 -73.275 ;
        RECT -43.685 -74.965 -43.355 -74.635 ;
        RECT -43.685 -76.325 -43.355 -75.995 ;
        RECT -43.685 -77.685 -43.355 -77.355 ;
        RECT -43.685 -79.045 -43.355 -78.715 ;
        RECT -43.685 -80.405 -43.355 -80.075 ;
        RECT -43.685 -81.765 -43.355 -81.435 ;
        RECT -43.685 -83.125 -43.355 -82.795 ;
        RECT -43.685 -84.485 -43.355 -84.155 ;
        RECT -43.685 -85.845 -43.355 -85.515 ;
        RECT -43.685 -87.205 -43.355 -86.875 ;
        RECT -43.685 -88.565 -43.355 -88.235 ;
        RECT -43.685 -89.925 -43.355 -89.595 ;
        RECT -43.685 -92.645 -43.355 -92.315 ;
        RECT -43.685 -94.005 -43.355 -93.675 ;
        RECT -43.685 -95.365 -43.355 -95.035 ;
        RECT -43.685 -96.725 -43.355 -96.395 ;
        RECT -43.685 -98.73 -43.355 -98.4 ;
        RECT -43.685 -99.445 -43.355 -99.115 ;
        RECT -43.685 -102.165 -43.355 -101.835 ;
        RECT -43.685 -103.525 -43.355 -103.195 ;
        RECT -43.685 -104.885 -43.355 -104.555 ;
        RECT -43.685 -106.87 -43.355 -106.54 ;
        RECT -43.685 -107.605 -43.355 -107.275 ;
        RECT -43.685 -108.965 -43.355 -108.635 ;
        RECT -43.685 -113.045 -43.355 -112.715 ;
        RECT -43.685 -114.405 -43.355 -114.075 ;
        RECT -43.685 -115.765 -43.355 -115.435 ;
        RECT -43.685 -117.125 -43.355 -116.795 ;
        RECT -43.685 -118.485 -43.355 -118.155 ;
        RECT -43.685 -122.565 -43.355 -122.235 ;
        RECT -43.685 -123.925 -43.355 -123.595 ;
        RECT -43.685 -125.285 -43.355 -124.955 ;
        RECT -43.685 -126.645 -43.355 -126.315 ;
        RECT -43.685 -128.005 -43.355 -127.675 ;
        RECT -43.685 -129.365 -43.355 -129.035 ;
        RECT -43.685 -130.725 -43.355 -130.395 ;
        RECT -43.685 -132.085 -43.355 -131.755 ;
        RECT -43.685 -133.445 -43.355 -133.115 ;
        RECT -43.685 -134.805 -43.355 -134.475 ;
        RECT -43.685 -136.165 -43.355 -135.835 ;
        RECT -43.685 -137.525 -43.355 -137.195 ;
        RECT -43.685 -138.885 -43.355 -138.555 ;
        RECT -43.685 -140.245 -43.355 -139.915 ;
        RECT -43.685 -141.605 -43.355 -141.275 ;
        RECT -43.685 -142.965 -43.355 -142.635 ;
        RECT -43.685 -144.325 -43.355 -143.995 ;
        RECT -43.685 -145.685 -43.355 -145.355 ;
        RECT -43.685 -147.045 -43.355 -146.715 ;
        RECT -43.685 -148.405 -43.355 -148.075 ;
        RECT -43.685 -149.765 -43.355 -149.435 ;
        RECT -43.685 -151.125 -43.355 -150.795 ;
        RECT -43.685 -152.485 -43.355 -152.155 ;
        RECT -43.685 -153.845 -43.355 -153.515 ;
        RECT -43.685 -155.205 -43.355 -154.875 ;
        RECT -43.685 -156.565 -43.355 -156.235 ;
        RECT -43.685 -157.925 -43.355 -157.595 ;
        RECT -43.685 -159.285 -43.355 -158.955 ;
        RECT -43.685 -160.645 -43.355 -160.315 ;
        RECT -43.685 -162.005 -43.355 -161.675 ;
        RECT -43.685 -163.365 -43.355 -163.035 ;
        RECT -43.685 -164.725 -43.355 -164.395 ;
        RECT -43.685 -166.085 -43.355 -165.755 ;
        RECT -43.685 -167.445 -43.355 -167.115 ;
        RECT -43.685 -170.165 -43.355 -169.835 ;
        RECT -43.685 -172.885 -43.355 -172.555 ;
        RECT -43.685 -174.245 -43.355 -173.915 ;
        RECT -43.685 -175.725 -43.355 -175.395 ;
        RECT -43.685 -176.965 -43.355 -176.635 ;
        RECT -43.685 -178.325 -43.355 -177.995 ;
        RECT -43.685 -180.57 -43.355 -179.44 ;
        RECT -43.68 -180.685 -43.36 -67.84 ;
    END
    PORT
      LAYER met3 ;
        RECT -42.325 241.32 -41.995 242.45 ;
        RECT -42.325 239.195 -41.995 239.525 ;
        RECT -42.325 237.835 -41.995 238.165 ;
        RECT -42.325 236.475 -41.995 236.805 ;
        RECT -42.325 235.115 -41.995 235.445 ;
        RECT -42.325 233.755 -41.995 234.085 ;
        RECT -42.325 232.395 -41.995 232.725 ;
        RECT -42.325 231.035 -41.995 231.365 ;
        RECT -42.325 229.675 -41.995 230.005 ;
        RECT -42.325 228.315 -41.995 228.645 ;
        RECT -42.325 226.955 -41.995 227.285 ;
        RECT -42.325 225.595 -41.995 225.925 ;
        RECT -42.325 224.235 -41.995 224.565 ;
        RECT -42.325 222.875 -41.995 223.205 ;
        RECT -42.325 221.515 -41.995 221.845 ;
        RECT -42.325 220.155 -41.995 220.485 ;
        RECT -42.325 218.795 -41.995 219.125 ;
        RECT -42.325 217.435 -41.995 217.765 ;
        RECT -42.325 216.075 -41.995 216.405 ;
        RECT -42.325 214.715 -41.995 215.045 ;
        RECT -42.325 213.355 -41.995 213.685 ;
        RECT -42.325 211.995 -41.995 212.325 ;
        RECT -42.325 210.635 -41.995 210.965 ;
        RECT -42.325 209.275 -41.995 209.605 ;
        RECT -42.325 207.915 -41.995 208.245 ;
        RECT -42.325 206.555 -41.995 206.885 ;
        RECT -42.325 205.195 -41.995 205.525 ;
        RECT -42.325 203.835 -41.995 204.165 ;
        RECT -42.325 202.475 -41.995 202.805 ;
        RECT -42.325 201.115 -41.995 201.445 ;
        RECT -42.325 199.755 -41.995 200.085 ;
        RECT -42.325 198.395 -41.995 198.725 ;
        RECT -42.325 197.035 -41.995 197.365 ;
        RECT -42.325 195.675 -41.995 196.005 ;
        RECT -42.325 194.315 -41.995 194.645 ;
        RECT -42.325 192.955 -41.995 193.285 ;
        RECT -42.325 191.595 -41.995 191.925 ;
        RECT -42.325 190.235 -41.995 190.565 ;
        RECT -42.325 188.875 -41.995 189.205 ;
        RECT -42.325 187.515 -41.995 187.845 ;
        RECT -42.325 186.155 -41.995 186.485 ;
        RECT -42.325 184.795 -41.995 185.125 ;
        RECT -42.325 183.435 -41.995 183.765 ;
        RECT -42.325 182.075 -41.995 182.405 ;
        RECT -42.325 180.715 -41.995 181.045 ;
        RECT -42.325 179.355 -41.995 179.685 ;
        RECT -42.325 177.995 -41.995 178.325 ;
        RECT -42.325 176.635 -41.995 176.965 ;
        RECT -42.325 175.275 -41.995 175.605 ;
        RECT -42.325 173.915 -41.995 174.245 ;
        RECT -42.325 172.555 -41.995 172.885 ;
        RECT -42.325 171.195 -41.995 171.525 ;
        RECT -42.325 169.835 -41.995 170.165 ;
        RECT -42.325 168.475 -41.995 168.805 ;
        RECT -42.325 167.115 -41.995 167.445 ;
        RECT -42.325 165.755 -41.995 166.085 ;
        RECT -42.325 164.395 -41.995 164.725 ;
        RECT -42.325 163.035 -41.995 163.365 ;
        RECT -42.325 161.675 -41.995 162.005 ;
        RECT -42.325 160.315 -41.995 160.645 ;
        RECT -42.325 158.955 -41.995 159.285 ;
        RECT -42.325 157.595 -41.995 157.925 ;
        RECT -42.325 156.235 -41.995 156.565 ;
        RECT -42.325 154.875 -41.995 155.205 ;
        RECT -42.325 153.515 -41.995 153.845 ;
        RECT -42.325 152.155 -41.995 152.485 ;
        RECT -42.325 150.795 -41.995 151.125 ;
        RECT -42.325 149.435 -41.995 149.765 ;
        RECT -42.325 148.075 -41.995 148.405 ;
        RECT -42.325 146.715 -41.995 147.045 ;
        RECT -42.325 145.355 -41.995 145.685 ;
        RECT -42.325 143.995 -41.995 144.325 ;
        RECT -42.325 142.635 -41.995 142.965 ;
        RECT -42.325 141.275 -41.995 141.605 ;
        RECT -42.325 139.915 -41.995 140.245 ;
        RECT -42.325 138.555 -41.995 138.885 ;
        RECT -42.325 137.195 -41.995 137.525 ;
        RECT -42.325 135.835 -41.995 136.165 ;
        RECT -42.325 134.475 -41.995 134.805 ;
        RECT -42.325 133.115 -41.995 133.445 ;
        RECT -42.325 131.755 -41.995 132.085 ;
        RECT -42.325 130.395 -41.995 130.725 ;
        RECT -42.325 129.035 -41.995 129.365 ;
        RECT -42.325 127.675 -41.995 128.005 ;
        RECT -42.325 126.315 -41.995 126.645 ;
        RECT -42.325 124.955 -41.995 125.285 ;
        RECT -42.325 123.595 -41.995 123.925 ;
        RECT -42.325 122.235 -41.995 122.565 ;
        RECT -42.325 120.875 -41.995 121.205 ;
        RECT -42.325 119.515 -41.995 119.845 ;
        RECT -42.325 118.155 -41.995 118.485 ;
        RECT -42.325 116.795 -41.995 117.125 ;
        RECT -42.325 115.435 -41.995 115.765 ;
        RECT -42.325 114.075 -41.995 114.405 ;
        RECT -42.325 112.715 -41.995 113.045 ;
        RECT -42.325 111.355 -41.995 111.685 ;
        RECT -42.325 109.995 -41.995 110.325 ;
        RECT -42.325 108.635 -41.995 108.965 ;
        RECT -42.325 107.275 -41.995 107.605 ;
        RECT -42.325 105.915 -41.995 106.245 ;
        RECT -42.325 104.555 -41.995 104.885 ;
        RECT -42.325 103.195 -41.995 103.525 ;
        RECT -42.325 101.835 -41.995 102.165 ;
        RECT -42.325 100.475 -41.995 100.805 ;
        RECT -42.325 99.115 -41.995 99.445 ;
        RECT -42.325 97.755 -41.995 98.085 ;
        RECT -42.325 96.395 -41.995 96.725 ;
        RECT -42.325 95.035 -41.995 95.365 ;
        RECT -42.325 93.675 -41.995 94.005 ;
        RECT -42.325 92.315 -41.995 92.645 ;
        RECT -42.325 90.955 -41.995 91.285 ;
        RECT -42.325 89.595 -41.995 89.925 ;
        RECT -42.325 88.235 -41.995 88.565 ;
        RECT -42.325 86.875 -41.995 87.205 ;
        RECT -42.325 85.515 -41.995 85.845 ;
        RECT -42.325 84.155 -41.995 84.485 ;
        RECT -42.325 82.795 -41.995 83.125 ;
        RECT -42.325 81.435 -41.995 81.765 ;
        RECT -42.325 80.075 -41.995 80.405 ;
        RECT -42.325 78.715 -41.995 79.045 ;
        RECT -42.325 77.355 -41.995 77.685 ;
        RECT -42.325 75.995 -41.995 76.325 ;
        RECT -42.325 74.635 -41.995 74.965 ;
        RECT -42.325 73.275 -41.995 73.605 ;
        RECT -42.325 71.915 -41.995 72.245 ;
        RECT -42.325 70.555 -41.995 70.885 ;
        RECT -42.325 69.195 -41.995 69.525 ;
        RECT -42.325 67.835 -41.995 68.165 ;
        RECT -42.325 66.475 -41.995 66.805 ;
        RECT -42.325 65.115 -41.995 65.445 ;
        RECT -42.325 63.755 -41.995 64.085 ;
        RECT -42.325 62.395 -41.995 62.725 ;
        RECT -42.325 61.035 -41.995 61.365 ;
        RECT -42.325 59.675 -41.995 60.005 ;
        RECT -42.325 58.315 -41.995 58.645 ;
        RECT -42.325 56.955 -41.995 57.285 ;
        RECT -42.325 55.595 -41.995 55.925 ;
        RECT -42.325 54.235 -41.995 54.565 ;
        RECT -42.325 52.875 -41.995 53.205 ;
        RECT -42.325 51.515 -41.995 51.845 ;
        RECT -42.325 50.155 -41.995 50.485 ;
        RECT -42.325 48.795 -41.995 49.125 ;
        RECT -42.325 47.435 -41.995 47.765 ;
        RECT -42.325 46.075 -41.995 46.405 ;
        RECT -42.325 44.715 -41.995 45.045 ;
        RECT -42.325 43.355 -41.995 43.685 ;
        RECT -42.325 41.995 -41.995 42.325 ;
        RECT -42.325 40.635 -41.995 40.965 ;
        RECT -42.325 39.275 -41.995 39.605 ;
        RECT -42.325 37.915 -41.995 38.245 ;
        RECT -42.325 36.555 -41.995 36.885 ;
        RECT -42.325 35.195 -41.995 35.525 ;
        RECT -42.325 33.835 -41.995 34.165 ;
        RECT -42.325 32.475 -41.995 32.805 ;
        RECT -42.325 31.115 -41.995 31.445 ;
        RECT -42.325 29.755 -41.995 30.085 ;
        RECT -42.325 28.395 -41.995 28.725 ;
        RECT -42.325 27.035 -41.995 27.365 ;
        RECT -42.325 25.675 -41.995 26.005 ;
        RECT -42.325 24.315 -41.995 24.645 ;
        RECT -42.325 22.955 -41.995 23.285 ;
        RECT -42.325 21.595 -41.995 21.925 ;
        RECT -42.325 20.235 -41.995 20.565 ;
        RECT -42.325 18.875 -41.995 19.205 ;
        RECT -42.325 17.515 -41.995 17.845 ;
        RECT -42.325 16.155 -41.995 16.485 ;
        RECT -42.325 14.795 -41.995 15.125 ;
        RECT -42.325 13.435 -41.995 13.765 ;
        RECT -42.325 12.075 -41.995 12.405 ;
        RECT -42.325 10.715 -41.995 11.045 ;
        RECT -42.325 9.355 -41.995 9.685 ;
        RECT -42.325 7.995 -41.995 8.325 ;
        RECT -42.325 6.635 -41.995 6.965 ;
        RECT -42.325 5.275 -41.995 5.605 ;
        RECT -42.325 3.915 -41.995 4.245 ;
        RECT -42.325 2.555 -41.995 2.885 ;
        RECT -42.325 1.195 -41.995 1.525 ;
        RECT -42.325 -0.165 -41.995 0.165 ;
        RECT -42.325 -5.605 -41.995 -5.275 ;
        RECT -42.325 -6.965 -41.995 -6.635 ;
        RECT -42.325 -11.045 -41.995 -10.715 ;
        RECT -42.325 -15.125 -41.995 -14.795 ;
        RECT -42.325 -16.485 -41.995 -16.155 ;
        RECT -42.325 -17.845 -41.995 -17.515 ;
        RECT -42.325 -19.205 -41.995 -18.875 ;
        RECT -42.325 -20.565 -41.995 -20.235 ;
        RECT -42.325 -21.925 -41.995 -21.595 ;
        RECT -42.325 -23.285 -41.995 -22.955 ;
        RECT -42.325 -24.645 -41.995 -24.315 ;
        RECT -42.325 -31.445 -41.995 -31.115 ;
        RECT -42.325 -32.805 -41.995 -32.475 ;
        RECT -42.325 -35.525 -41.995 -35.195 ;
        RECT -42.325 -36.885 -41.995 -36.555 ;
        RECT -42.325 -37.93 -41.995 -37.6 ;
        RECT -42.325 -40.965 -41.995 -40.635 ;
        RECT -42.325 -42.77 -41.995 -42.44 ;
        RECT -42.325 -43.685 -41.995 -43.355 ;
        RECT -42.325 -50.485 -41.995 -50.155 ;
        RECT -42.325 -51.845 -41.995 -51.515 ;
        RECT -42.325 -54.565 -41.995 -54.235 ;
        RECT -42.325 -55.925 -41.995 -55.595 ;
        RECT -42.325 -60.005 -41.995 -59.675 ;
        RECT -42.325 -66.805 -41.995 -66.475 ;
        RECT -42.325 -69.525 -41.995 -69.195 ;
        RECT -42.325 -70.885 -41.995 -70.555 ;
        RECT -42.325 -72.245 -41.995 -71.915 ;
        RECT -42.325 -73.605 -41.995 -73.275 ;
        RECT -42.325 -74.965 -41.995 -74.635 ;
        RECT -42.325 -76.325 -41.995 -75.995 ;
        RECT -42.325 -77.685 -41.995 -77.355 ;
        RECT -42.325 -79.045 -41.995 -78.715 ;
        RECT -42.325 -80.405 -41.995 -80.075 ;
        RECT -42.325 -81.765 -41.995 -81.435 ;
        RECT -42.325 -83.125 -41.995 -82.795 ;
        RECT -42.325 -84.485 -41.995 -84.155 ;
        RECT -42.325 -85.845 -41.995 -85.515 ;
        RECT -42.325 -87.205 -41.995 -86.875 ;
        RECT -42.325 -88.565 -41.995 -88.235 ;
        RECT -42.325 -89.925 -41.995 -89.595 ;
        RECT -42.325 -92.645 -41.995 -92.315 ;
        RECT -42.325 -94.005 -41.995 -93.675 ;
        RECT -42.325 -95.365 -41.995 -95.035 ;
        RECT -42.325 -96.725 -41.995 -96.395 ;
        RECT -42.325 -98.73 -41.995 -98.4 ;
        RECT -42.325 -99.445 -41.995 -99.115 ;
        RECT -42.325 -102.165 -41.995 -101.835 ;
        RECT -42.325 -103.525 -41.995 -103.195 ;
        RECT -42.325 -104.885 -41.995 -104.555 ;
        RECT -42.325 -106.87 -41.995 -106.54 ;
        RECT -42.325 -107.605 -41.995 -107.275 ;
        RECT -42.325 -108.965 -41.995 -108.635 ;
        RECT -42.32 -112.36 -42 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -42.325 -174.245 -41.995 -173.915 ;
        RECT -42.325 -175.725 -41.995 -175.395 ;
        RECT -42.325 -176.965 -41.995 -176.635 ;
        RECT -42.325 -178.325 -41.995 -177.995 ;
        RECT -42.325 -180.57 -41.995 -179.44 ;
        RECT -42.32 -180.685 -42 -173.915 ;
    END
    PORT
      LAYER met3 ;
        RECT -40.965 241.32 -40.635 242.45 ;
        RECT -40.965 239.195 -40.635 239.525 ;
        RECT -40.965 237.835 -40.635 238.165 ;
        RECT -40.965 236.475 -40.635 236.805 ;
        RECT -40.965 235.115 -40.635 235.445 ;
        RECT -40.965 233.755 -40.635 234.085 ;
        RECT -40.965 232.395 -40.635 232.725 ;
        RECT -40.965 231.035 -40.635 231.365 ;
        RECT -40.965 229.675 -40.635 230.005 ;
        RECT -40.965 228.315 -40.635 228.645 ;
        RECT -40.965 226.955 -40.635 227.285 ;
        RECT -40.965 225.595 -40.635 225.925 ;
        RECT -40.965 224.235 -40.635 224.565 ;
        RECT -40.965 222.875 -40.635 223.205 ;
        RECT -40.965 221.515 -40.635 221.845 ;
        RECT -40.965 220.155 -40.635 220.485 ;
        RECT -40.965 218.795 -40.635 219.125 ;
        RECT -40.965 217.435 -40.635 217.765 ;
        RECT -40.965 216.075 -40.635 216.405 ;
        RECT -40.965 214.715 -40.635 215.045 ;
        RECT -40.965 213.355 -40.635 213.685 ;
        RECT -40.965 211.995 -40.635 212.325 ;
        RECT -40.965 210.635 -40.635 210.965 ;
        RECT -40.965 209.275 -40.635 209.605 ;
        RECT -40.965 207.915 -40.635 208.245 ;
        RECT -40.965 206.555 -40.635 206.885 ;
        RECT -40.965 205.195 -40.635 205.525 ;
        RECT -40.965 203.835 -40.635 204.165 ;
        RECT -40.965 202.475 -40.635 202.805 ;
        RECT -40.965 201.115 -40.635 201.445 ;
        RECT -40.965 199.755 -40.635 200.085 ;
        RECT -40.965 198.395 -40.635 198.725 ;
        RECT -40.965 197.035 -40.635 197.365 ;
        RECT -40.965 195.675 -40.635 196.005 ;
        RECT -40.965 194.315 -40.635 194.645 ;
        RECT -40.965 192.955 -40.635 193.285 ;
        RECT -40.965 191.595 -40.635 191.925 ;
        RECT -40.965 190.235 -40.635 190.565 ;
        RECT -40.965 188.875 -40.635 189.205 ;
        RECT -40.965 187.515 -40.635 187.845 ;
        RECT -40.965 186.155 -40.635 186.485 ;
        RECT -40.965 184.795 -40.635 185.125 ;
        RECT -40.965 183.435 -40.635 183.765 ;
        RECT -40.965 182.075 -40.635 182.405 ;
        RECT -40.965 180.715 -40.635 181.045 ;
        RECT -40.965 179.355 -40.635 179.685 ;
        RECT -40.965 177.995 -40.635 178.325 ;
        RECT -40.965 176.635 -40.635 176.965 ;
        RECT -40.965 175.275 -40.635 175.605 ;
        RECT -40.965 173.915 -40.635 174.245 ;
        RECT -40.965 172.555 -40.635 172.885 ;
        RECT -40.965 171.195 -40.635 171.525 ;
        RECT -40.965 169.835 -40.635 170.165 ;
        RECT -40.965 168.475 -40.635 168.805 ;
        RECT -40.965 167.115 -40.635 167.445 ;
        RECT -40.965 165.755 -40.635 166.085 ;
        RECT -40.965 164.395 -40.635 164.725 ;
        RECT -40.965 163.035 -40.635 163.365 ;
        RECT -40.965 161.675 -40.635 162.005 ;
        RECT -40.965 160.315 -40.635 160.645 ;
        RECT -40.965 158.955 -40.635 159.285 ;
        RECT -40.965 157.595 -40.635 157.925 ;
        RECT -40.965 156.235 -40.635 156.565 ;
        RECT -40.965 154.875 -40.635 155.205 ;
        RECT -40.965 153.515 -40.635 153.845 ;
        RECT -40.965 152.155 -40.635 152.485 ;
        RECT -40.965 150.795 -40.635 151.125 ;
        RECT -40.965 149.435 -40.635 149.765 ;
        RECT -40.965 148.075 -40.635 148.405 ;
        RECT -40.965 146.715 -40.635 147.045 ;
        RECT -40.965 145.355 -40.635 145.685 ;
        RECT -40.965 143.995 -40.635 144.325 ;
        RECT -40.965 142.635 -40.635 142.965 ;
        RECT -40.965 141.275 -40.635 141.605 ;
        RECT -40.965 139.915 -40.635 140.245 ;
        RECT -40.965 138.555 -40.635 138.885 ;
        RECT -40.965 137.195 -40.635 137.525 ;
        RECT -40.965 135.835 -40.635 136.165 ;
        RECT -40.965 134.475 -40.635 134.805 ;
        RECT -40.965 133.115 -40.635 133.445 ;
        RECT -40.965 131.755 -40.635 132.085 ;
        RECT -40.965 130.395 -40.635 130.725 ;
        RECT -40.965 129.035 -40.635 129.365 ;
        RECT -40.965 127.675 -40.635 128.005 ;
        RECT -40.965 126.315 -40.635 126.645 ;
        RECT -40.965 124.955 -40.635 125.285 ;
        RECT -40.965 123.595 -40.635 123.925 ;
        RECT -40.965 122.235 -40.635 122.565 ;
        RECT -40.965 120.875 -40.635 121.205 ;
        RECT -40.965 119.515 -40.635 119.845 ;
        RECT -40.965 118.155 -40.635 118.485 ;
        RECT -40.965 116.795 -40.635 117.125 ;
        RECT -40.965 115.435 -40.635 115.765 ;
        RECT -40.965 114.075 -40.635 114.405 ;
        RECT -40.965 112.715 -40.635 113.045 ;
        RECT -40.965 111.355 -40.635 111.685 ;
        RECT -40.965 109.995 -40.635 110.325 ;
        RECT -40.965 108.635 -40.635 108.965 ;
        RECT -40.965 107.275 -40.635 107.605 ;
        RECT -40.965 105.915 -40.635 106.245 ;
        RECT -40.965 104.555 -40.635 104.885 ;
        RECT -40.965 103.195 -40.635 103.525 ;
        RECT -40.965 101.835 -40.635 102.165 ;
        RECT -40.965 100.475 -40.635 100.805 ;
        RECT -40.965 99.115 -40.635 99.445 ;
        RECT -40.965 97.755 -40.635 98.085 ;
        RECT -40.965 96.395 -40.635 96.725 ;
        RECT -40.965 95.035 -40.635 95.365 ;
        RECT -40.965 93.675 -40.635 94.005 ;
        RECT -40.965 92.315 -40.635 92.645 ;
        RECT -40.965 90.955 -40.635 91.285 ;
        RECT -40.965 89.595 -40.635 89.925 ;
        RECT -40.965 88.235 -40.635 88.565 ;
        RECT -40.965 86.875 -40.635 87.205 ;
        RECT -40.965 85.515 -40.635 85.845 ;
        RECT -40.965 84.155 -40.635 84.485 ;
        RECT -40.965 82.795 -40.635 83.125 ;
        RECT -40.965 81.435 -40.635 81.765 ;
        RECT -40.965 80.075 -40.635 80.405 ;
        RECT -40.965 78.715 -40.635 79.045 ;
        RECT -40.965 77.355 -40.635 77.685 ;
        RECT -40.965 75.995 -40.635 76.325 ;
        RECT -40.965 74.635 -40.635 74.965 ;
        RECT -40.965 73.275 -40.635 73.605 ;
        RECT -40.965 71.915 -40.635 72.245 ;
        RECT -40.965 70.555 -40.635 70.885 ;
        RECT -40.965 69.195 -40.635 69.525 ;
        RECT -40.965 67.835 -40.635 68.165 ;
        RECT -40.965 66.475 -40.635 66.805 ;
        RECT -40.965 65.115 -40.635 65.445 ;
        RECT -40.965 63.755 -40.635 64.085 ;
        RECT -40.965 62.395 -40.635 62.725 ;
        RECT -40.965 61.035 -40.635 61.365 ;
        RECT -40.965 59.675 -40.635 60.005 ;
        RECT -40.965 58.315 -40.635 58.645 ;
        RECT -40.965 56.955 -40.635 57.285 ;
        RECT -40.965 55.595 -40.635 55.925 ;
        RECT -40.965 54.235 -40.635 54.565 ;
        RECT -40.965 52.875 -40.635 53.205 ;
        RECT -40.965 51.515 -40.635 51.845 ;
        RECT -40.965 50.155 -40.635 50.485 ;
        RECT -40.965 48.795 -40.635 49.125 ;
        RECT -40.965 47.435 -40.635 47.765 ;
        RECT -40.965 46.075 -40.635 46.405 ;
        RECT -40.965 44.715 -40.635 45.045 ;
        RECT -40.965 43.355 -40.635 43.685 ;
        RECT -40.965 41.995 -40.635 42.325 ;
        RECT -40.965 40.635 -40.635 40.965 ;
        RECT -40.965 39.275 -40.635 39.605 ;
        RECT -40.965 37.915 -40.635 38.245 ;
        RECT -40.965 36.555 -40.635 36.885 ;
        RECT -40.965 35.195 -40.635 35.525 ;
        RECT -40.965 33.835 -40.635 34.165 ;
        RECT -40.965 32.475 -40.635 32.805 ;
        RECT -40.965 31.115 -40.635 31.445 ;
        RECT -40.965 29.755 -40.635 30.085 ;
        RECT -40.965 28.395 -40.635 28.725 ;
        RECT -40.965 27.035 -40.635 27.365 ;
        RECT -40.965 25.675 -40.635 26.005 ;
        RECT -40.965 24.315 -40.635 24.645 ;
        RECT -40.965 22.955 -40.635 23.285 ;
        RECT -40.965 21.595 -40.635 21.925 ;
        RECT -40.965 20.235 -40.635 20.565 ;
        RECT -40.965 18.875 -40.635 19.205 ;
        RECT -40.965 17.515 -40.635 17.845 ;
        RECT -40.965 16.155 -40.635 16.485 ;
        RECT -40.965 14.795 -40.635 15.125 ;
        RECT -40.965 13.435 -40.635 13.765 ;
        RECT -40.965 12.075 -40.635 12.405 ;
        RECT -40.965 10.715 -40.635 11.045 ;
        RECT -40.965 9.355 -40.635 9.685 ;
        RECT -40.965 7.995 -40.635 8.325 ;
        RECT -40.965 6.635 -40.635 6.965 ;
        RECT -40.965 5.275 -40.635 5.605 ;
        RECT -40.965 3.915 -40.635 4.245 ;
        RECT -40.965 2.555 -40.635 2.885 ;
        RECT -40.965 1.195 -40.635 1.525 ;
        RECT -40.965 -0.165 -40.635 0.165 ;
        RECT -40.965 -4.245 -40.635 -3.915 ;
        RECT -40.965 -5.605 -40.635 -5.275 ;
        RECT -40.965 -6.965 -40.635 -6.635 ;
        RECT -40.965 -11.045 -40.635 -10.715 ;
        RECT -40.965 -15.125 -40.635 -14.795 ;
        RECT -40.965 -16.485 -40.635 -16.155 ;
        RECT -40.965 -17.845 -40.635 -17.515 ;
        RECT -40.965 -19.205 -40.635 -18.875 ;
        RECT -40.965 -20.565 -40.635 -20.235 ;
        RECT -40.965 -21.925 -40.635 -21.595 ;
        RECT -40.965 -23.285 -40.635 -22.955 ;
        RECT -40.965 -24.645 -40.635 -24.315 ;
        RECT -40.965 -31.445 -40.635 -31.115 ;
        RECT -40.965 -32.805 -40.635 -32.475 ;
        RECT -40.965 -35.525 -40.635 -35.195 ;
        RECT -40.965 -36.885 -40.635 -36.555 ;
        RECT -40.965 -37.93 -40.635 -37.6 ;
        RECT -40.965 -40.965 -40.635 -40.635 ;
        RECT -40.965 -42.77 -40.635 -42.44 ;
        RECT -40.965 -43.685 -40.635 -43.355 ;
        RECT -40.965 -50.485 -40.635 -50.155 ;
        RECT -40.965 -51.845 -40.635 -51.515 ;
        RECT -40.965 -54.565 -40.635 -54.235 ;
        RECT -40.965 -55.925 -40.635 -55.595 ;
        RECT -40.965 -60.005 -40.635 -59.675 ;
        RECT -40.965 -66.805 -40.635 -66.475 ;
        RECT -40.965 -69.525 -40.635 -69.195 ;
        RECT -40.965 -70.885 -40.635 -70.555 ;
        RECT -40.965 -72.245 -40.635 -71.915 ;
        RECT -40.965 -73.605 -40.635 -73.275 ;
        RECT -40.965 -74.965 -40.635 -74.635 ;
        RECT -40.965 -76.325 -40.635 -75.995 ;
        RECT -40.965 -77.685 -40.635 -77.355 ;
        RECT -40.965 -79.045 -40.635 -78.715 ;
        RECT -40.965 -80.405 -40.635 -80.075 ;
        RECT -40.965 -81.765 -40.635 -81.435 ;
        RECT -40.965 -83.125 -40.635 -82.795 ;
        RECT -40.965 -84.485 -40.635 -84.155 ;
        RECT -40.965 -85.845 -40.635 -85.515 ;
        RECT -40.965 -87.205 -40.635 -86.875 ;
        RECT -40.965 -88.565 -40.635 -88.235 ;
        RECT -40.965 -89.925 -40.635 -89.595 ;
        RECT -40.965 -92.645 -40.635 -92.315 ;
        RECT -40.965 -94.005 -40.635 -93.675 ;
        RECT -40.965 -95.365 -40.635 -95.035 ;
        RECT -40.965 -96.725 -40.635 -96.395 ;
        RECT -40.965 -98.73 -40.635 -98.4 ;
        RECT -40.965 -99.445 -40.635 -99.115 ;
        RECT -40.965 -102.165 -40.635 -101.835 ;
        RECT -40.965 -103.525 -40.635 -103.195 ;
        RECT -40.965 -104.885 -40.635 -104.555 ;
        RECT -40.965 -106.87 -40.635 -106.54 ;
        RECT -40.965 -107.605 -40.635 -107.275 ;
        RECT -40.965 -108.965 -40.635 -108.635 ;
        RECT -40.965 -114.405 -40.635 -114.075 ;
        RECT -40.965 -115.765 -40.635 -115.435 ;
        RECT -40.965 -117.125 -40.635 -116.795 ;
        RECT -40.965 -118.485 -40.635 -118.155 ;
        RECT -40.965 -122.565 -40.635 -122.235 ;
        RECT -40.965 -123.925 -40.635 -123.595 ;
        RECT -40.965 -125.285 -40.635 -124.955 ;
        RECT -40.965 -126.645 -40.635 -126.315 ;
        RECT -40.965 -128.005 -40.635 -127.675 ;
        RECT -40.965 -129.365 -40.635 -129.035 ;
        RECT -40.965 -130.725 -40.635 -130.395 ;
        RECT -40.965 -132.085 -40.635 -131.755 ;
        RECT -40.965 -133.445 -40.635 -133.115 ;
        RECT -40.965 -134.805 -40.635 -134.475 ;
        RECT -40.965 -136.165 -40.635 -135.835 ;
        RECT -40.965 -137.525 -40.635 -137.195 ;
        RECT -40.965 -138.885 -40.635 -138.555 ;
        RECT -40.965 -140.245 -40.635 -139.915 ;
        RECT -40.965 -141.605 -40.635 -141.275 ;
        RECT -40.965 -142.965 -40.635 -142.635 ;
        RECT -40.965 -144.325 -40.635 -143.995 ;
        RECT -40.965 -145.685 -40.635 -145.355 ;
        RECT -40.965 -147.045 -40.635 -146.715 ;
        RECT -40.965 -148.405 -40.635 -148.075 ;
        RECT -40.965 -151.125 -40.635 -150.795 ;
        RECT -40.965 -152.485 -40.635 -152.155 ;
        RECT -40.965 -153.845 -40.635 -153.515 ;
        RECT -40.965 -155.205 -40.635 -154.875 ;
        RECT -40.965 -157.925 -40.635 -157.595 ;
        RECT -40.965 -159.285 -40.635 -158.955 ;
        RECT -40.965 -160.645 -40.635 -160.315 ;
        RECT -40.965 -162.005 -40.635 -161.675 ;
        RECT -40.965 -163.365 -40.635 -163.035 ;
        RECT -40.965 -164.725 -40.635 -164.395 ;
        RECT -40.965 -166.085 -40.635 -165.755 ;
        RECT -40.965 -167.445 -40.635 -167.115 ;
        RECT -40.965 -170.165 -40.635 -169.835 ;
        RECT -40.965 -174.245 -40.635 -173.915 ;
        RECT -40.965 -176.965 -40.635 -176.635 ;
        RECT -40.965 -178.325 -40.635 -177.995 ;
        RECT -40.965 -180.57 -40.635 -179.44 ;
        RECT -40.96 -180.685 -40.64 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -39.605 48.795 -39.275 49.125 ;
        RECT -39.605 47.435 -39.275 47.765 ;
        RECT -39.605 46.075 -39.275 46.405 ;
        RECT -39.605 44.715 -39.275 45.045 ;
        RECT -39.605 43.355 -39.275 43.685 ;
        RECT -39.605 41.995 -39.275 42.325 ;
        RECT -39.605 40.635 -39.275 40.965 ;
        RECT -39.605 39.275 -39.275 39.605 ;
        RECT -39.605 37.915 -39.275 38.245 ;
        RECT -39.605 36.555 -39.275 36.885 ;
        RECT -39.605 35.195 -39.275 35.525 ;
        RECT -39.605 33.835 -39.275 34.165 ;
        RECT -39.605 32.475 -39.275 32.805 ;
        RECT -39.605 31.115 -39.275 31.445 ;
        RECT -39.605 29.755 -39.275 30.085 ;
        RECT -39.605 28.395 -39.275 28.725 ;
        RECT -39.605 27.035 -39.275 27.365 ;
        RECT -39.605 25.675 -39.275 26.005 ;
        RECT -39.605 24.315 -39.275 24.645 ;
        RECT -39.605 22.955 -39.275 23.285 ;
        RECT -39.605 21.595 -39.275 21.925 ;
        RECT -39.605 20.235 -39.275 20.565 ;
        RECT -39.605 18.875 -39.275 19.205 ;
        RECT -39.605 17.515 -39.275 17.845 ;
        RECT -39.605 16.155 -39.275 16.485 ;
        RECT -39.605 14.795 -39.275 15.125 ;
        RECT -39.605 13.435 -39.275 13.765 ;
        RECT -39.605 12.075 -39.275 12.405 ;
        RECT -39.605 10.715 -39.275 11.045 ;
        RECT -39.605 9.355 -39.275 9.685 ;
        RECT -39.605 7.995 -39.275 8.325 ;
        RECT -39.605 6.635 -39.275 6.965 ;
        RECT -39.605 5.275 -39.275 5.605 ;
        RECT -39.605 3.915 -39.275 4.245 ;
        RECT -39.605 2.555 -39.275 2.885 ;
        RECT -39.605 1.195 -39.275 1.525 ;
        RECT -39.605 -0.165 -39.275 0.165 ;
        RECT -39.605 -2.885 -39.275 -2.555 ;
        RECT -39.605 -4.245 -39.275 -3.915 ;
        RECT -39.605 -5.605 -39.275 -5.275 ;
        RECT -39.605 -11.045 -39.275 -10.715 ;
        RECT -39.605 -15.125 -39.275 -14.795 ;
        RECT -39.605 -16.485 -39.275 -16.155 ;
        RECT -39.605 -17.845 -39.275 -17.515 ;
        RECT -39.605 -19.205 -39.275 -18.875 ;
        RECT -39.605 -20.565 -39.275 -20.235 ;
        RECT -39.605 -21.925 -39.275 -21.595 ;
        RECT -39.605 -23.285 -39.275 -22.955 ;
        RECT -39.605 -24.645 -39.275 -24.315 ;
        RECT -39.605 -31.445 -39.275 -31.115 ;
        RECT -39.605 -32.805 -39.275 -32.475 ;
        RECT -39.605 -35.525 -39.275 -35.195 ;
        RECT -39.605 -36.885 -39.275 -36.555 ;
        RECT -39.605 -37.93 -39.275 -37.6 ;
        RECT -39.605 -40.965 -39.275 -40.635 ;
        RECT -39.605 -42.77 -39.275 -42.44 ;
        RECT -39.605 -43.685 -39.275 -43.355 ;
        RECT -39.605 -50.485 -39.275 -50.155 ;
        RECT -39.605 -51.845 -39.275 -51.515 ;
        RECT -39.605 -54.565 -39.275 -54.235 ;
        RECT -39.605 -55.925 -39.275 -55.595 ;
        RECT -39.605 -60.005 -39.275 -59.675 ;
        RECT -39.605 -66.805 -39.275 -66.475 ;
        RECT -39.605 -69.525 -39.275 -69.195 ;
        RECT -39.605 -70.885 -39.275 -70.555 ;
        RECT -39.605 -72.245 -39.275 -71.915 ;
        RECT -39.605 -73.605 -39.275 -73.275 ;
        RECT -39.605 -74.965 -39.275 -74.635 ;
        RECT -39.605 -76.325 -39.275 -75.995 ;
        RECT -39.605 -77.685 -39.275 -77.355 ;
        RECT -39.605 -79.045 -39.275 -78.715 ;
        RECT -39.605 -80.405 -39.275 -80.075 ;
        RECT -39.605 -81.765 -39.275 -81.435 ;
        RECT -39.605 -83.125 -39.275 -82.795 ;
        RECT -39.605 -84.485 -39.275 -84.155 ;
        RECT -39.605 -85.845 -39.275 -85.515 ;
        RECT -39.605 -87.205 -39.275 -86.875 ;
        RECT -39.605 -88.565 -39.275 -88.235 ;
        RECT -39.605 -89.925 -39.275 -89.595 ;
        RECT -39.605 -92.645 -39.275 -92.315 ;
        RECT -39.605 -94.005 -39.275 -93.675 ;
        RECT -39.605 -95.365 -39.275 -95.035 ;
        RECT -39.605 -96.725 -39.275 -96.395 ;
        RECT -39.605 -98.73 -39.275 -98.4 ;
        RECT -39.605 -99.445 -39.275 -99.115 ;
        RECT -39.605 -102.165 -39.275 -101.835 ;
        RECT -39.605 -103.525 -39.275 -103.195 ;
        RECT -39.605 -104.885 -39.275 -104.555 ;
        RECT -39.605 -106.87 -39.275 -106.54 ;
        RECT -39.605 -107.605 -39.275 -107.275 ;
        RECT -39.605 -108.965 -39.275 -108.635 ;
        RECT -39.605 -114.405 -39.275 -114.075 ;
        RECT -39.605 -115.765 -39.275 -115.435 ;
        RECT -39.605 -117.125 -39.275 -116.795 ;
        RECT -39.605 -118.485 -39.275 -118.155 ;
        RECT -39.605 -122.565 -39.275 -122.235 ;
        RECT -39.605 -123.925 -39.275 -123.595 ;
        RECT -39.605 -125.285 -39.275 -124.955 ;
        RECT -39.605 -126.645 -39.275 -126.315 ;
        RECT -39.605 -128.005 -39.275 -127.675 ;
        RECT -39.605 -129.365 -39.275 -129.035 ;
        RECT -39.605 -130.725 -39.275 -130.395 ;
        RECT -39.605 -133.445 -39.275 -133.115 ;
        RECT -39.605 -134.805 -39.275 -134.475 ;
        RECT -39.605 -136.165 -39.275 -135.835 ;
        RECT -39.605 -137.525 -39.275 -137.195 ;
        RECT -39.605 -138.885 -39.275 -138.555 ;
        RECT -39.605 -140.245 -39.275 -139.915 ;
        RECT -39.605 -141.605 -39.275 -141.275 ;
        RECT -39.605 -142.965 -39.275 -142.635 ;
        RECT -39.605 -144.325 -39.275 -143.995 ;
        RECT -39.605 -145.685 -39.275 -145.355 ;
        RECT -39.605 -147.045 -39.275 -146.715 ;
        RECT -39.605 -148.405 -39.275 -148.075 ;
        RECT -39.605 -151.125 -39.275 -150.795 ;
        RECT -39.605 -152.485 -39.275 -152.155 ;
        RECT -39.605 -155.205 -39.275 -154.875 ;
        RECT -39.605 -157.925 -39.275 -157.595 ;
        RECT -39.605 -159.285 -39.275 -158.955 ;
        RECT -39.605 -160.645 -39.275 -160.315 ;
        RECT -39.605 -162.005 -39.275 -161.675 ;
        RECT -39.605 -163.365 -39.275 -163.035 ;
        RECT -39.605 -164.725 -39.275 -164.395 ;
        RECT -39.605 -166.085 -39.275 -165.755 ;
        RECT -39.605 -167.445 -39.275 -167.115 ;
        RECT -39.605 -170.165 -39.275 -169.835 ;
        RECT -39.605 -174.245 -39.275 -173.915 ;
        RECT -39.605 -175.725 -39.275 -175.395 ;
        RECT -39.605 -176.965 -39.275 -176.635 ;
        RECT -39.605 -178.325 -39.275 -177.995 ;
        RECT -39.605 -180.57 -39.275 -179.44 ;
        RECT -39.6 -180.685 -39.28 242.565 ;
        RECT -39.605 241.32 -39.275 242.45 ;
        RECT -39.605 239.195 -39.275 239.525 ;
        RECT -39.605 237.835 -39.275 238.165 ;
        RECT -39.605 236.475 -39.275 236.805 ;
        RECT -39.605 235.115 -39.275 235.445 ;
        RECT -39.605 233.755 -39.275 234.085 ;
        RECT -39.605 232.395 -39.275 232.725 ;
        RECT -39.605 231.035 -39.275 231.365 ;
        RECT -39.605 229.675 -39.275 230.005 ;
        RECT -39.605 228.315 -39.275 228.645 ;
        RECT -39.605 226.955 -39.275 227.285 ;
        RECT -39.605 225.595 -39.275 225.925 ;
        RECT -39.605 224.235 -39.275 224.565 ;
        RECT -39.605 222.875 -39.275 223.205 ;
        RECT -39.605 221.515 -39.275 221.845 ;
        RECT -39.605 220.155 -39.275 220.485 ;
        RECT -39.605 218.795 -39.275 219.125 ;
        RECT -39.605 217.435 -39.275 217.765 ;
        RECT -39.605 216.075 -39.275 216.405 ;
        RECT -39.605 214.715 -39.275 215.045 ;
        RECT -39.605 213.355 -39.275 213.685 ;
        RECT -39.605 211.995 -39.275 212.325 ;
        RECT -39.605 210.635 -39.275 210.965 ;
        RECT -39.605 209.275 -39.275 209.605 ;
        RECT -39.605 207.915 -39.275 208.245 ;
        RECT -39.605 206.555 -39.275 206.885 ;
        RECT -39.605 205.195 -39.275 205.525 ;
        RECT -39.605 203.835 -39.275 204.165 ;
        RECT -39.605 202.475 -39.275 202.805 ;
        RECT -39.605 201.115 -39.275 201.445 ;
        RECT -39.605 199.755 -39.275 200.085 ;
        RECT -39.605 198.395 -39.275 198.725 ;
        RECT -39.605 197.035 -39.275 197.365 ;
        RECT -39.605 195.675 -39.275 196.005 ;
        RECT -39.605 194.315 -39.275 194.645 ;
        RECT -39.605 192.955 -39.275 193.285 ;
        RECT -39.605 191.595 -39.275 191.925 ;
        RECT -39.605 190.235 -39.275 190.565 ;
        RECT -39.605 188.875 -39.275 189.205 ;
        RECT -39.605 187.515 -39.275 187.845 ;
        RECT -39.605 186.155 -39.275 186.485 ;
        RECT -39.605 184.795 -39.275 185.125 ;
        RECT -39.605 183.435 -39.275 183.765 ;
        RECT -39.605 182.075 -39.275 182.405 ;
        RECT -39.605 180.715 -39.275 181.045 ;
        RECT -39.605 179.355 -39.275 179.685 ;
        RECT -39.605 177.995 -39.275 178.325 ;
        RECT -39.605 176.635 -39.275 176.965 ;
        RECT -39.605 175.275 -39.275 175.605 ;
        RECT -39.605 173.915 -39.275 174.245 ;
        RECT -39.605 172.555 -39.275 172.885 ;
        RECT -39.605 171.195 -39.275 171.525 ;
        RECT -39.605 169.835 -39.275 170.165 ;
        RECT -39.605 168.475 -39.275 168.805 ;
        RECT -39.605 167.115 -39.275 167.445 ;
        RECT -39.605 165.755 -39.275 166.085 ;
        RECT -39.605 164.395 -39.275 164.725 ;
        RECT -39.605 163.035 -39.275 163.365 ;
        RECT -39.605 161.675 -39.275 162.005 ;
        RECT -39.605 160.315 -39.275 160.645 ;
        RECT -39.605 158.955 -39.275 159.285 ;
        RECT -39.605 157.595 -39.275 157.925 ;
        RECT -39.605 156.235 -39.275 156.565 ;
        RECT -39.605 154.875 -39.275 155.205 ;
        RECT -39.605 153.515 -39.275 153.845 ;
        RECT -39.605 152.155 -39.275 152.485 ;
        RECT -39.605 150.795 -39.275 151.125 ;
        RECT -39.605 149.435 -39.275 149.765 ;
        RECT -39.605 148.075 -39.275 148.405 ;
        RECT -39.605 146.715 -39.275 147.045 ;
        RECT -39.605 145.355 -39.275 145.685 ;
        RECT -39.605 143.995 -39.275 144.325 ;
        RECT -39.605 142.635 -39.275 142.965 ;
        RECT -39.605 141.275 -39.275 141.605 ;
        RECT -39.605 139.915 -39.275 140.245 ;
        RECT -39.605 138.555 -39.275 138.885 ;
        RECT -39.605 137.195 -39.275 137.525 ;
        RECT -39.605 135.835 -39.275 136.165 ;
        RECT -39.605 134.475 -39.275 134.805 ;
        RECT -39.605 133.115 -39.275 133.445 ;
        RECT -39.605 131.755 -39.275 132.085 ;
        RECT -39.605 130.395 -39.275 130.725 ;
        RECT -39.605 129.035 -39.275 129.365 ;
        RECT -39.605 127.675 -39.275 128.005 ;
        RECT -39.605 126.315 -39.275 126.645 ;
        RECT -39.605 124.955 -39.275 125.285 ;
        RECT -39.605 123.595 -39.275 123.925 ;
        RECT -39.605 122.235 -39.275 122.565 ;
        RECT -39.605 120.875 -39.275 121.205 ;
        RECT -39.605 119.515 -39.275 119.845 ;
        RECT -39.605 118.155 -39.275 118.485 ;
        RECT -39.605 116.795 -39.275 117.125 ;
        RECT -39.605 115.435 -39.275 115.765 ;
        RECT -39.605 114.075 -39.275 114.405 ;
        RECT -39.605 112.715 -39.275 113.045 ;
        RECT -39.605 111.355 -39.275 111.685 ;
        RECT -39.605 109.995 -39.275 110.325 ;
        RECT -39.605 108.635 -39.275 108.965 ;
        RECT -39.605 107.275 -39.275 107.605 ;
        RECT -39.605 105.915 -39.275 106.245 ;
        RECT -39.605 104.555 -39.275 104.885 ;
        RECT -39.605 103.195 -39.275 103.525 ;
        RECT -39.605 101.835 -39.275 102.165 ;
        RECT -39.605 100.475 -39.275 100.805 ;
        RECT -39.605 99.115 -39.275 99.445 ;
        RECT -39.605 97.755 -39.275 98.085 ;
        RECT -39.605 96.395 -39.275 96.725 ;
        RECT -39.605 95.035 -39.275 95.365 ;
        RECT -39.605 93.675 -39.275 94.005 ;
        RECT -39.605 92.315 -39.275 92.645 ;
        RECT -39.605 90.955 -39.275 91.285 ;
        RECT -39.605 89.595 -39.275 89.925 ;
        RECT -39.605 88.235 -39.275 88.565 ;
        RECT -39.605 86.875 -39.275 87.205 ;
        RECT -39.605 85.515 -39.275 85.845 ;
        RECT -39.605 84.155 -39.275 84.485 ;
        RECT -39.605 82.795 -39.275 83.125 ;
        RECT -39.605 81.435 -39.275 81.765 ;
        RECT -39.605 80.075 -39.275 80.405 ;
        RECT -39.605 78.715 -39.275 79.045 ;
        RECT -39.605 77.355 -39.275 77.685 ;
        RECT -39.605 75.995 -39.275 76.325 ;
        RECT -39.605 74.635 -39.275 74.965 ;
        RECT -39.605 73.275 -39.275 73.605 ;
        RECT -39.605 71.915 -39.275 72.245 ;
        RECT -39.605 70.555 -39.275 70.885 ;
        RECT -39.605 69.195 -39.275 69.525 ;
        RECT -39.605 67.835 -39.275 68.165 ;
        RECT -39.605 66.475 -39.275 66.805 ;
        RECT -39.605 65.115 -39.275 65.445 ;
        RECT -39.605 63.755 -39.275 64.085 ;
        RECT -39.605 62.395 -39.275 62.725 ;
        RECT -39.605 61.035 -39.275 61.365 ;
        RECT -39.605 59.675 -39.275 60.005 ;
        RECT -39.605 58.315 -39.275 58.645 ;
        RECT -39.605 56.955 -39.275 57.285 ;
        RECT -39.605 55.595 -39.275 55.925 ;
        RECT -39.605 54.235 -39.275 54.565 ;
        RECT -39.605 52.875 -39.275 53.205 ;
        RECT -39.605 51.515 -39.275 51.845 ;
        RECT -39.605 50.155 -39.275 50.485 ;
    END
    PORT
      LAYER met3 ;
        RECT -49.125 241.32 -48.795 242.45 ;
        RECT -49.125 239.195 -48.795 239.525 ;
        RECT -49.125 237.835 -48.795 238.165 ;
        RECT -49.125 236.475 -48.795 236.805 ;
        RECT -49.125 235.115 -48.795 235.445 ;
        RECT -49.125 233.755 -48.795 234.085 ;
        RECT -49.125 232.395 -48.795 232.725 ;
        RECT -49.125 231.035 -48.795 231.365 ;
        RECT -49.125 229.675 -48.795 230.005 ;
        RECT -49.125 228.315 -48.795 228.645 ;
        RECT -49.125 226.955 -48.795 227.285 ;
        RECT -49.125 225.595 -48.795 225.925 ;
        RECT -49.125 224.235 -48.795 224.565 ;
        RECT -49.125 222.875 -48.795 223.205 ;
        RECT -49.125 221.515 -48.795 221.845 ;
        RECT -49.125 220.155 -48.795 220.485 ;
        RECT -49.125 218.795 -48.795 219.125 ;
        RECT -49.125 217.435 -48.795 217.765 ;
        RECT -49.125 216.075 -48.795 216.405 ;
        RECT -49.125 214.715 -48.795 215.045 ;
        RECT -49.125 213.355 -48.795 213.685 ;
        RECT -49.125 211.995 -48.795 212.325 ;
        RECT -49.125 210.635 -48.795 210.965 ;
        RECT -49.125 209.275 -48.795 209.605 ;
        RECT -49.125 207.915 -48.795 208.245 ;
        RECT -49.125 206.555 -48.795 206.885 ;
        RECT -49.125 205.195 -48.795 205.525 ;
        RECT -49.125 203.835 -48.795 204.165 ;
        RECT -49.125 202.475 -48.795 202.805 ;
        RECT -49.125 201.115 -48.795 201.445 ;
        RECT -49.125 199.755 -48.795 200.085 ;
        RECT -49.125 198.395 -48.795 198.725 ;
        RECT -49.125 197.035 -48.795 197.365 ;
        RECT -49.125 195.675 -48.795 196.005 ;
        RECT -49.125 194.315 -48.795 194.645 ;
        RECT -49.125 192.955 -48.795 193.285 ;
        RECT -49.125 191.595 -48.795 191.925 ;
        RECT -49.125 190.235 -48.795 190.565 ;
        RECT -49.125 188.875 -48.795 189.205 ;
        RECT -49.125 187.515 -48.795 187.845 ;
        RECT -49.125 186.155 -48.795 186.485 ;
        RECT -49.125 184.795 -48.795 185.125 ;
        RECT -49.125 183.435 -48.795 183.765 ;
        RECT -49.125 182.075 -48.795 182.405 ;
        RECT -49.125 180.715 -48.795 181.045 ;
        RECT -49.125 179.355 -48.795 179.685 ;
        RECT -49.125 177.995 -48.795 178.325 ;
        RECT -49.125 176.635 -48.795 176.965 ;
        RECT -49.125 175.275 -48.795 175.605 ;
        RECT -49.125 173.915 -48.795 174.245 ;
        RECT -49.125 172.555 -48.795 172.885 ;
        RECT -49.125 171.195 -48.795 171.525 ;
        RECT -49.125 169.835 -48.795 170.165 ;
        RECT -49.125 168.475 -48.795 168.805 ;
        RECT -49.125 167.115 -48.795 167.445 ;
        RECT -49.125 165.755 -48.795 166.085 ;
        RECT -49.125 164.395 -48.795 164.725 ;
        RECT -49.125 163.035 -48.795 163.365 ;
        RECT -49.125 161.675 -48.795 162.005 ;
        RECT -49.125 160.315 -48.795 160.645 ;
        RECT -49.125 158.955 -48.795 159.285 ;
        RECT -49.125 157.595 -48.795 157.925 ;
        RECT -49.125 156.235 -48.795 156.565 ;
        RECT -49.125 154.875 -48.795 155.205 ;
        RECT -49.125 153.515 -48.795 153.845 ;
        RECT -49.125 152.155 -48.795 152.485 ;
        RECT -49.125 150.795 -48.795 151.125 ;
        RECT -49.125 149.435 -48.795 149.765 ;
        RECT -49.125 148.075 -48.795 148.405 ;
        RECT -49.125 146.715 -48.795 147.045 ;
        RECT -49.125 145.355 -48.795 145.685 ;
        RECT -49.125 143.995 -48.795 144.325 ;
        RECT -49.125 142.635 -48.795 142.965 ;
        RECT -49.125 141.275 -48.795 141.605 ;
        RECT -49.125 139.915 -48.795 140.245 ;
        RECT -49.125 138.555 -48.795 138.885 ;
        RECT -49.125 137.225 -48.795 137.555 ;
        RECT -49.125 135.175 -48.795 135.505 ;
        RECT -49.125 132.815 -48.795 133.145 ;
        RECT -49.125 131.665 -48.795 131.995 ;
        RECT -49.125 129.655 -48.795 129.985 ;
        RECT -49.125 128.505 -48.795 128.835 ;
        RECT -49.125 126.495 -48.795 126.825 ;
        RECT -49.125 125.345 -48.795 125.675 ;
        RECT -49.125 123.335 -48.795 123.665 ;
        RECT -49.125 122.185 -48.795 122.515 ;
        RECT -49.125 120.175 -48.795 120.505 ;
        RECT -49.125 119.025 -48.795 119.355 ;
        RECT -49.125 117.185 -48.795 117.515 ;
        RECT -49.125 115.865 -48.795 116.195 ;
        RECT -49.125 113.855 -48.795 114.185 ;
        RECT -49.125 112.705 -48.795 113.035 ;
        RECT -49.125 110.695 -48.795 111.025 ;
        RECT -49.125 109.545 -48.795 109.875 ;
        RECT -49.125 107.535 -48.795 107.865 ;
        RECT -49.125 106.385 -48.795 106.715 ;
        RECT -49.125 104.375 -48.795 104.705 ;
        RECT -49.125 103.225 -48.795 103.555 ;
        RECT -49.125 100.865 -48.795 101.195 ;
        RECT -49.125 98.81 -48.795 99.14 ;
        RECT -49.125 97.755 -48.795 98.085 ;
        RECT -49.125 96.395 -48.795 96.725 ;
        RECT -49.125 95.035 -48.795 95.365 ;
        RECT -49.125 93.675 -48.795 94.005 ;
        RECT -49.125 92.315 -48.795 92.645 ;
        RECT -49.125 90.955 -48.795 91.285 ;
        RECT -49.125 89.595 -48.795 89.925 ;
        RECT -49.125 88.235 -48.795 88.565 ;
        RECT -49.125 86.875 -48.795 87.205 ;
        RECT -49.125 85.515 -48.795 85.845 ;
        RECT -49.125 84.155 -48.795 84.485 ;
        RECT -49.125 82.795 -48.795 83.125 ;
        RECT -49.125 81.435 -48.795 81.765 ;
        RECT -49.125 80.075 -48.795 80.405 ;
        RECT -49.125 78.715 -48.795 79.045 ;
        RECT -49.125 77.355 -48.795 77.685 ;
        RECT -49.125 75.995 -48.795 76.325 ;
        RECT -49.125 74.635 -48.795 74.965 ;
        RECT -49.125 73.275 -48.795 73.605 ;
        RECT -49.125 71.915 -48.795 72.245 ;
        RECT -49.125 70.555 -48.795 70.885 ;
        RECT -49.125 69.195 -48.795 69.525 ;
        RECT -49.125 67.835 -48.795 68.165 ;
        RECT -49.125 66.475 -48.795 66.805 ;
        RECT -49.125 65.115 -48.795 65.445 ;
        RECT -49.125 63.755 -48.795 64.085 ;
        RECT -49.125 62.395 -48.795 62.725 ;
        RECT -49.125 61.035 -48.795 61.365 ;
        RECT -49.125 59.675 -48.795 60.005 ;
        RECT -49.125 58.315 -48.795 58.645 ;
        RECT -49.125 56.955 -48.795 57.285 ;
        RECT -49.125 55.595 -48.795 55.925 ;
        RECT -49.125 54.235 -48.795 54.565 ;
        RECT -49.125 52.875 -48.795 53.205 ;
        RECT -49.125 51.515 -48.795 51.845 ;
        RECT -49.125 50.155 -48.795 50.485 ;
        RECT -49.125 48.795 -48.795 49.125 ;
        RECT -49.125 47.435 -48.795 47.765 ;
        RECT -49.125 46.075 -48.795 46.405 ;
        RECT -49.125 44.715 -48.795 45.045 ;
        RECT -49.125 43.355 -48.795 43.685 ;
        RECT -49.125 41.995 -48.795 42.325 ;
        RECT -49.125 40.635 -48.795 40.965 ;
        RECT -49.125 39.275 -48.795 39.605 ;
        RECT -49.125 37.915 -48.795 38.245 ;
        RECT -49.125 36.555 -48.795 36.885 ;
        RECT -49.125 35.195 -48.795 35.525 ;
        RECT -49.125 33.835 -48.795 34.165 ;
        RECT -49.125 32.475 -48.795 32.805 ;
        RECT -49.125 31.115 -48.795 31.445 ;
        RECT -49.125 29.755 -48.795 30.085 ;
        RECT -49.125 28.395 -48.795 28.725 ;
        RECT -49.125 27.035 -48.795 27.365 ;
        RECT -49.125 25.675 -48.795 26.005 ;
        RECT -49.125 24.315 -48.795 24.645 ;
        RECT -49.125 22.955 -48.795 23.285 ;
        RECT -49.125 21.595 -48.795 21.925 ;
        RECT -49.125 20.235 -48.795 20.565 ;
        RECT -49.125 18.875 -48.795 19.205 ;
        RECT -49.125 17.515 -48.795 17.845 ;
        RECT -49.125 16.155 -48.795 16.485 ;
        RECT -49.125 14.795 -48.795 15.125 ;
        RECT -49.125 13.435 -48.795 13.765 ;
        RECT -49.125 12.075 -48.795 12.405 ;
        RECT -49.125 10.715 -48.795 11.045 ;
        RECT -49.125 9.355 -48.795 9.685 ;
        RECT -49.125 7.995 -48.795 8.325 ;
        RECT -49.125 6.635 -48.795 6.965 ;
        RECT -49.125 5.275 -48.795 5.605 ;
        RECT -49.125 3.915 -48.795 4.245 ;
        RECT -49.125 2.555 -48.795 2.885 ;
        RECT -49.125 1.195 -48.795 1.525 ;
        RECT -49.125 -0.165 -48.795 0.165 ;
        RECT -49.125 -2.885 -48.795 -2.555 ;
        RECT -49.125 -4.245 -48.795 -3.915 ;
        RECT -49.125 -5.605 -48.795 -5.275 ;
        RECT -49.125 -6.965 -48.795 -6.635 ;
        RECT -49.125 -8.325 -48.795 -7.995 ;
        RECT -49.125 -9.685 -48.795 -9.355 ;
        RECT -49.125 -11.045 -48.795 -10.715 ;
        RECT -49.125 -15.125 -48.795 -14.795 ;
        RECT -49.125 -16.485 -48.795 -16.155 ;
        RECT -49.125 -17.845 -48.795 -17.515 ;
        RECT -49.125 -19.205 -48.795 -18.875 ;
        RECT -49.125 -20.565 -48.795 -20.235 ;
        RECT -49.125 -21.925 -48.795 -21.595 ;
        RECT -49.125 -23.285 -48.795 -22.955 ;
        RECT -49.125 -24.645 -48.795 -24.315 ;
        RECT -49.125 -28.725 -48.795 -28.395 ;
        RECT -49.125 -30.085 -48.795 -29.755 ;
        RECT -49.125 -31.445 -48.795 -31.115 ;
        RECT -49.125 -32.805 -48.795 -32.475 ;
        RECT -49.125 -35.525 -48.795 -35.195 ;
        RECT -49.125 -36.885 -48.795 -36.555 ;
        RECT -49.125 -37.93 -48.795 -37.6 ;
        RECT -49.125 -40.965 -48.795 -40.635 ;
        RECT -49.125 -42.77 -48.795 -42.44 ;
        RECT -49.125 -43.685 -48.795 -43.355 ;
        RECT -49.125 -50.485 -48.795 -50.155 ;
        RECT -49.125 -51.845 -48.795 -51.515 ;
        RECT -49.125 -54.565 -48.795 -54.235 ;
        RECT -49.125 -55.925 -48.795 -55.595 ;
        RECT -49.125 -60.005 -48.795 -59.675 ;
        RECT -49.125 -66.805 -48.795 -66.475 ;
        RECT -49.125 -68.165 -48.795 -67.835 ;
        RECT -49.125 -69.525 -48.795 -69.195 ;
        RECT -49.125 -70.885 -48.795 -70.555 ;
        RECT -49.125 -72.245 -48.795 -71.915 ;
        RECT -49.125 -73.605 -48.795 -73.275 ;
        RECT -49.125 -74.965 -48.795 -74.635 ;
        RECT -49.125 -76.325 -48.795 -75.995 ;
        RECT -49.125 -77.685 -48.795 -77.355 ;
        RECT -49.125 -79.045 -48.795 -78.715 ;
        RECT -49.125 -80.405 -48.795 -80.075 ;
        RECT -49.125 -81.765 -48.795 -81.435 ;
        RECT -49.125 -83.125 -48.795 -82.795 ;
        RECT -49.125 -84.485 -48.795 -84.155 ;
        RECT -49.125 -85.845 -48.795 -85.515 ;
        RECT -49.125 -87.205 -48.795 -86.875 ;
        RECT -49.125 -88.565 -48.795 -88.235 ;
        RECT -49.125 -89.925 -48.795 -89.595 ;
        RECT -49.125 -92.645 -48.795 -92.315 ;
        RECT -49.125 -94.005 -48.795 -93.675 ;
        RECT -49.125 -95.365 -48.795 -95.035 ;
        RECT -49.125 -96.725 -48.795 -96.395 ;
        RECT -49.125 -98.73 -48.795 -98.4 ;
        RECT -49.125 -99.445 -48.795 -99.115 ;
        RECT -49.125 -102.165 -48.795 -101.835 ;
        RECT -49.125 -103.525 -48.795 -103.195 ;
        RECT -49.125 -104.885 -48.795 -104.555 ;
        RECT -49.125 -106.87 -48.795 -106.54 ;
        RECT -49.125 -107.605 -48.795 -107.275 ;
        RECT -49.125 -108.965 -48.795 -108.635 ;
        RECT -49.125 -114.405 -48.795 -114.075 ;
        RECT -49.125 -115.765 -48.795 -115.435 ;
        RECT -49.125 -117.125 -48.795 -116.795 ;
        RECT -49.125 -118.485 -48.795 -118.155 ;
        RECT -49.125 -122.565 -48.795 -122.235 ;
        RECT -49.125 -123.925 -48.795 -123.595 ;
        RECT -49.125 -125.285 -48.795 -124.955 ;
        RECT -49.125 -126.645 -48.795 -126.315 ;
        RECT -49.125 -128.005 -48.795 -127.675 ;
        RECT -49.125 -129.365 -48.795 -129.035 ;
        RECT -49.125 -130.725 -48.795 -130.395 ;
        RECT -49.125 -132.085 -48.795 -131.755 ;
        RECT -49.125 -133.445 -48.795 -133.115 ;
        RECT -49.125 -134.805 -48.795 -134.475 ;
        RECT -49.125 -136.165 -48.795 -135.835 ;
        RECT -49.125 -137.525 -48.795 -137.195 ;
        RECT -49.125 -138.885 -48.795 -138.555 ;
        RECT -49.125 -140.245 -48.795 -139.915 ;
        RECT -49.125 -141.605 -48.795 -141.275 ;
        RECT -49.125 -142.965 -48.795 -142.635 ;
        RECT -49.125 -144.325 -48.795 -143.995 ;
        RECT -49.125 -145.685 -48.795 -145.355 ;
        RECT -49.125 -147.045 -48.795 -146.715 ;
        RECT -49.125 -148.405 -48.795 -148.075 ;
        RECT -49.125 -149.765 -48.795 -149.435 ;
        RECT -49.125 -151.125 -48.795 -150.795 ;
        RECT -49.125 -152.485 -48.795 -152.155 ;
        RECT -49.125 -153.845 -48.795 -153.515 ;
        RECT -49.125 -155.205 -48.795 -154.875 ;
        RECT -49.125 -156.565 -48.795 -156.235 ;
        RECT -49.125 -157.925 -48.795 -157.595 ;
        RECT -49.125 -159.285 -48.795 -158.955 ;
        RECT -49.125 -160.645 -48.795 -160.315 ;
        RECT -49.125 -162.005 -48.795 -161.675 ;
        RECT -49.125 -163.365 -48.795 -163.035 ;
        RECT -49.125 -164.725 -48.795 -164.395 ;
        RECT -49.125 -166.085 -48.795 -165.755 ;
        RECT -49.125 -167.445 -48.795 -167.115 ;
        RECT -49.125 -170.165 -48.795 -169.835 ;
        RECT -49.125 -172.885 -48.795 -172.555 ;
        RECT -49.125 -174.245 -48.795 -173.915 ;
        RECT -49.125 -175.725 -48.795 -175.395 ;
        RECT -49.125 -176.965 -48.795 -176.635 ;
        RECT -49.125 -178.325 -48.795 -177.995 ;
        RECT -49.125 -180.57 -48.795 -179.44 ;
        RECT -49.12 -180.685 -48.8 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -47.765 241.32 -47.435 242.45 ;
        RECT -47.765 239.195 -47.435 239.525 ;
        RECT -47.765 237.835 -47.435 238.165 ;
        RECT -47.765 236.475 -47.435 236.805 ;
        RECT -47.765 235.115 -47.435 235.445 ;
        RECT -47.765 233.755 -47.435 234.085 ;
        RECT -47.765 232.395 -47.435 232.725 ;
        RECT -47.765 231.035 -47.435 231.365 ;
        RECT -47.765 229.675 -47.435 230.005 ;
        RECT -47.765 228.315 -47.435 228.645 ;
        RECT -47.765 226.955 -47.435 227.285 ;
        RECT -47.765 225.595 -47.435 225.925 ;
        RECT -47.765 224.235 -47.435 224.565 ;
        RECT -47.765 222.875 -47.435 223.205 ;
        RECT -47.765 221.515 -47.435 221.845 ;
        RECT -47.765 220.155 -47.435 220.485 ;
        RECT -47.765 218.795 -47.435 219.125 ;
        RECT -47.765 217.435 -47.435 217.765 ;
        RECT -47.765 216.075 -47.435 216.405 ;
        RECT -47.765 214.715 -47.435 215.045 ;
        RECT -47.765 213.355 -47.435 213.685 ;
        RECT -47.765 211.995 -47.435 212.325 ;
        RECT -47.765 210.635 -47.435 210.965 ;
        RECT -47.765 209.275 -47.435 209.605 ;
        RECT -47.765 207.915 -47.435 208.245 ;
        RECT -47.765 206.555 -47.435 206.885 ;
        RECT -47.765 205.195 -47.435 205.525 ;
        RECT -47.765 203.835 -47.435 204.165 ;
        RECT -47.765 202.475 -47.435 202.805 ;
        RECT -47.765 201.115 -47.435 201.445 ;
        RECT -47.765 199.755 -47.435 200.085 ;
        RECT -47.765 198.395 -47.435 198.725 ;
        RECT -47.765 197.035 -47.435 197.365 ;
        RECT -47.765 195.675 -47.435 196.005 ;
        RECT -47.765 194.315 -47.435 194.645 ;
        RECT -47.765 192.955 -47.435 193.285 ;
        RECT -47.765 191.595 -47.435 191.925 ;
        RECT -47.765 190.235 -47.435 190.565 ;
        RECT -47.765 188.875 -47.435 189.205 ;
        RECT -47.765 187.515 -47.435 187.845 ;
        RECT -47.765 186.155 -47.435 186.485 ;
        RECT -47.765 184.795 -47.435 185.125 ;
        RECT -47.765 183.435 -47.435 183.765 ;
        RECT -47.765 182.075 -47.435 182.405 ;
        RECT -47.765 180.715 -47.435 181.045 ;
        RECT -47.765 179.355 -47.435 179.685 ;
        RECT -47.765 177.995 -47.435 178.325 ;
        RECT -47.765 176.635 -47.435 176.965 ;
        RECT -47.765 175.275 -47.435 175.605 ;
        RECT -47.765 173.915 -47.435 174.245 ;
        RECT -47.765 172.555 -47.435 172.885 ;
        RECT -47.765 171.195 -47.435 171.525 ;
        RECT -47.765 169.835 -47.435 170.165 ;
        RECT -47.765 168.475 -47.435 168.805 ;
        RECT -47.765 167.115 -47.435 167.445 ;
        RECT -47.765 165.755 -47.435 166.085 ;
        RECT -47.765 164.395 -47.435 164.725 ;
        RECT -47.765 163.035 -47.435 163.365 ;
        RECT -47.765 161.675 -47.435 162.005 ;
        RECT -47.765 160.315 -47.435 160.645 ;
        RECT -47.765 158.955 -47.435 159.285 ;
        RECT -47.765 157.595 -47.435 157.925 ;
        RECT -47.765 156.235 -47.435 156.565 ;
        RECT -47.765 154.875 -47.435 155.205 ;
        RECT -47.765 153.515 -47.435 153.845 ;
        RECT -47.765 152.155 -47.435 152.485 ;
        RECT -47.765 150.795 -47.435 151.125 ;
        RECT -47.765 149.435 -47.435 149.765 ;
        RECT -47.765 148.075 -47.435 148.405 ;
        RECT -47.765 146.715 -47.435 147.045 ;
        RECT -47.765 145.355 -47.435 145.685 ;
        RECT -47.765 143.995 -47.435 144.325 ;
        RECT -47.765 142.635 -47.435 142.965 ;
        RECT -47.765 141.275 -47.435 141.605 ;
        RECT -47.765 139.915 -47.435 140.245 ;
        RECT -47.765 138.555 -47.435 138.885 ;
        RECT -47.765 97.755 -47.435 98.085 ;
        RECT -47.765 96.395 -47.435 96.725 ;
        RECT -47.765 95.035 -47.435 95.365 ;
        RECT -47.765 93.675 -47.435 94.005 ;
        RECT -47.765 92.315 -47.435 92.645 ;
        RECT -47.765 90.955 -47.435 91.285 ;
        RECT -47.765 89.595 -47.435 89.925 ;
        RECT -47.765 88.235 -47.435 88.565 ;
        RECT -47.765 86.875 -47.435 87.205 ;
        RECT -47.765 85.515 -47.435 85.845 ;
        RECT -47.765 84.155 -47.435 84.485 ;
        RECT -47.765 82.795 -47.435 83.125 ;
        RECT -47.765 81.435 -47.435 81.765 ;
        RECT -47.765 80.075 -47.435 80.405 ;
        RECT -47.765 78.715 -47.435 79.045 ;
        RECT -47.765 77.355 -47.435 77.685 ;
        RECT -47.765 75.995 -47.435 76.325 ;
        RECT -47.765 74.635 -47.435 74.965 ;
        RECT -47.765 73.275 -47.435 73.605 ;
        RECT -47.765 71.915 -47.435 72.245 ;
        RECT -47.765 70.555 -47.435 70.885 ;
        RECT -47.765 69.195 -47.435 69.525 ;
        RECT -47.765 67.835 -47.435 68.165 ;
        RECT -47.765 66.475 -47.435 66.805 ;
        RECT -47.765 65.115 -47.435 65.445 ;
        RECT -47.765 63.755 -47.435 64.085 ;
        RECT -47.765 62.395 -47.435 62.725 ;
        RECT -47.765 61.035 -47.435 61.365 ;
        RECT -47.765 59.675 -47.435 60.005 ;
        RECT -47.765 58.315 -47.435 58.645 ;
        RECT -47.765 56.955 -47.435 57.285 ;
        RECT -47.765 55.595 -47.435 55.925 ;
        RECT -47.765 54.235 -47.435 54.565 ;
        RECT -47.765 52.875 -47.435 53.205 ;
        RECT -47.765 51.515 -47.435 51.845 ;
        RECT -47.765 50.155 -47.435 50.485 ;
        RECT -47.765 48.795 -47.435 49.125 ;
        RECT -47.765 47.435 -47.435 47.765 ;
        RECT -47.765 46.075 -47.435 46.405 ;
        RECT -47.765 44.715 -47.435 45.045 ;
        RECT -47.765 43.355 -47.435 43.685 ;
        RECT -47.765 41.995 -47.435 42.325 ;
        RECT -47.765 40.635 -47.435 40.965 ;
        RECT -47.765 39.275 -47.435 39.605 ;
        RECT -47.765 37.915 -47.435 38.245 ;
        RECT -47.765 36.555 -47.435 36.885 ;
        RECT -47.765 35.195 -47.435 35.525 ;
        RECT -47.765 33.835 -47.435 34.165 ;
        RECT -47.765 32.475 -47.435 32.805 ;
        RECT -47.765 31.115 -47.435 31.445 ;
        RECT -47.765 29.755 -47.435 30.085 ;
        RECT -47.765 28.395 -47.435 28.725 ;
        RECT -47.765 27.035 -47.435 27.365 ;
        RECT -47.765 25.675 -47.435 26.005 ;
        RECT -47.765 24.315 -47.435 24.645 ;
        RECT -47.765 22.955 -47.435 23.285 ;
        RECT -47.765 21.595 -47.435 21.925 ;
        RECT -47.765 20.235 -47.435 20.565 ;
        RECT -47.765 18.875 -47.435 19.205 ;
        RECT -47.765 17.515 -47.435 17.845 ;
        RECT -47.765 16.155 -47.435 16.485 ;
        RECT -47.765 14.795 -47.435 15.125 ;
        RECT -47.765 13.435 -47.435 13.765 ;
        RECT -47.765 12.075 -47.435 12.405 ;
        RECT -47.765 10.715 -47.435 11.045 ;
        RECT -47.765 9.355 -47.435 9.685 ;
        RECT -47.765 7.995 -47.435 8.325 ;
        RECT -47.765 6.635 -47.435 6.965 ;
        RECT -47.765 5.275 -47.435 5.605 ;
        RECT -47.765 3.915 -47.435 4.245 ;
        RECT -47.765 2.555 -47.435 2.885 ;
        RECT -47.765 1.195 -47.435 1.525 ;
        RECT -47.765 -0.165 -47.435 0.165 ;
        RECT -47.765 -2.885 -47.435 -2.555 ;
        RECT -47.765 -4.245 -47.435 -3.915 ;
        RECT -47.765 -5.605 -47.435 -5.275 ;
        RECT -47.765 -6.965 -47.435 -6.635 ;
        RECT -47.765 -8.325 -47.435 -7.995 ;
        RECT -47.765 -9.685 -47.435 -9.355 ;
        RECT -47.765 -11.045 -47.435 -10.715 ;
        RECT -47.765 -15.125 -47.435 -14.795 ;
        RECT -47.765 -16.485 -47.435 -16.155 ;
        RECT -47.765 -17.845 -47.435 -17.515 ;
        RECT -47.765 -19.205 -47.435 -18.875 ;
        RECT -47.765 -20.565 -47.435 -20.235 ;
        RECT -47.765 -21.925 -47.435 -21.595 ;
        RECT -47.765 -23.285 -47.435 -22.955 ;
        RECT -47.765 -24.645 -47.435 -24.315 ;
        RECT -47.765 -28.725 -47.435 -28.395 ;
        RECT -47.765 -31.445 -47.435 -31.115 ;
        RECT -47.765 -32.805 -47.435 -32.475 ;
        RECT -47.765 -35.525 -47.435 -35.195 ;
        RECT -47.765 -36.885 -47.435 -36.555 ;
        RECT -47.765 -37.93 -47.435 -37.6 ;
        RECT -47.765 -40.965 -47.435 -40.635 ;
        RECT -47.765 -42.77 -47.435 -42.44 ;
        RECT -47.765 -43.685 -47.435 -43.355 ;
        RECT -47.765 -50.485 -47.435 -50.155 ;
        RECT -47.765 -51.845 -47.435 -51.515 ;
        RECT -47.765 -54.565 -47.435 -54.235 ;
        RECT -47.765 -55.925 -47.435 -55.595 ;
        RECT -47.765 -60.005 -47.435 -59.675 ;
        RECT -47.765 -66.805 -47.435 -66.475 ;
        RECT -47.765 -68.165 -47.435 -67.835 ;
        RECT -47.765 -69.525 -47.435 -69.195 ;
        RECT -47.765 -70.885 -47.435 -70.555 ;
        RECT -47.765 -72.245 -47.435 -71.915 ;
        RECT -47.765 -73.605 -47.435 -73.275 ;
        RECT -47.765 -74.965 -47.435 -74.635 ;
        RECT -47.765 -76.325 -47.435 -75.995 ;
        RECT -47.765 -77.685 -47.435 -77.355 ;
        RECT -47.765 -79.045 -47.435 -78.715 ;
        RECT -47.765 -80.405 -47.435 -80.075 ;
        RECT -47.765 -81.765 -47.435 -81.435 ;
        RECT -47.765 -83.125 -47.435 -82.795 ;
        RECT -47.765 -84.485 -47.435 -84.155 ;
        RECT -47.765 -85.845 -47.435 -85.515 ;
        RECT -47.765 -87.205 -47.435 -86.875 ;
        RECT -47.765 -88.565 -47.435 -88.235 ;
        RECT -47.765 -89.925 -47.435 -89.595 ;
        RECT -47.765 -92.645 -47.435 -92.315 ;
        RECT -47.765 -94.005 -47.435 -93.675 ;
        RECT -47.765 -95.365 -47.435 -95.035 ;
        RECT -47.765 -96.725 -47.435 -96.395 ;
        RECT -47.765 -98.73 -47.435 -98.4 ;
        RECT -47.765 -99.445 -47.435 -99.115 ;
        RECT -47.765 -102.165 -47.435 -101.835 ;
        RECT -47.765 -103.525 -47.435 -103.195 ;
        RECT -47.765 -104.885 -47.435 -104.555 ;
        RECT -47.765 -106.87 -47.435 -106.54 ;
        RECT -47.765 -107.605 -47.435 -107.275 ;
        RECT -47.765 -108.965 -47.435 -108.635 ;
        RECT -47.765 -113.045 -47.435 -112.715 ;
        RECT -47.765 -114.405 -47.435 -114.075 ;
        RECT -47.765 -115.765 -47.435 -115.435 ;
        RECT -47.765 -117.125 -47.435 -116.795 ;
        RECT -47.765 -118.485 -47.435 -118.155 ;
        RECT -47.765 -122.565 -47.435 -122.235 ;
        RECT -47.765 -123.925 -47.435 -123.595 ;
        RECT -47.765 -125.285 -47.435 -124.955 ;
        RECT -47.765 -126.645 -47.435 -126.315 ;
        RECT -47.765 -128.005 -47.435 -127.675 ;
        RECT -47.765 -129.365 -47.435 -129.035 ;
        RECT -47.765 -130.725 -47.435 -130.395 ;
        RECT -47.765 -132.085 -47.435 -131.755 ;
        RECT -47.765 -133.445 -47.435 -133.115 ;
        RECT -47.765 -134.805 -47.435 -134.475 ;
        RECT -47.765 -136.165 -47.435 -135.835 ;
        RECT -47.765 -137.525 -47.435 -137.195 ;
        RECT -47.765 -138.885 -47.435 -138.555 ;
        RECT -47.765 -140.245 -47.435 -139.915 ;
        RECT -47.765 -141.605 -47.435 -141.275 ;
        RECT -47.765 -142.965 -47.435 -142.635 ;
        RECT -47.765 -144.325 -47.435 -143.995 ;
        RECT -47.765 -145.685 -47.435 -145.355 ;
        RECT -47.765 -147.045 -47.435 -146.715 ;
        RECT -47.765 -148.405 -47.435 -148.075 ;
        RECT -47.765 -149.765 -47.435 -149.435 ;
        RECT -47.765 -151.125 -47.435 -150.795 ;
        RECT -47.765 -152.485 -47.435 -152.155 ;
        RECT -47.765 -153.845 -47.435 -153.515 ;
        RECT -47.765 -155.205 -47.435 -154.875 ;
        RECT -47.765 -156.565 -47.435 -156.235 ;
        RECT -47.765 -157.925 -47.435 -157.595 ;
        RECT -47.765 -159.285 -47.435 -158.955 ;
        RECT -47.765 -160.645 -47.435 -160.315 ;
        RECT -47.765 -162.005 -47.435 -161.675 ;
        RECT -47.765 -163.365 -47.435 -163.035 ;
        RECT -47.765 -164.725 -47.435 -164.395 ;
        RECT -47.765 -166.085 -47.435 -165.755 ;
        RECT -47.765 -167.445 -47.435 -167.115 ;
        RECT -47.765 -170.165 -47.435 -169.835 ;
        RECT -47.765 -174.245 -47.435 -173.915 ;
        RECT -47.765 -175.725 -47.435 -175.395 ;
        RECT -47.765 -176.965 -47.435 -176.635 ;
        RECT -47.765 -178.325 -47.435 -177.995 ;
        RECT -47.765 -180.57 -47.435 -179.44 ;
        RECT -47.76 -180.685 -47.44 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -46.405 241.32 -46.075 242.45 ;
        RECT -46.405 239.195 -46.075 239.525 ;
        RECT -46.405 237.835 -46.075 238.165 ;
        RECT -46.405 236.475 -46.075 236.805 ;
        RECT -46.405 235.115 -46.075 235.445 ;
        RECT -46.405 233.755 -46.075 234.085 ;
        RECT -46.405 232.395 -46.075 232.725 ;
        RECT -46.405 231.035 -46.075 231.365 ;
        RECT -46.405 229.675 -46.075 230.005 ;
        RECT -46.405 228.315 -46.075 228.645 ;
        RECT -46.405 226.955 -46.075 227.285 ;
        RECT -46.405 225.595 -46.075 225.925 ;
        RECT -46.405 224.235 -46.075 224.565 ;
        RECT -46.405 222.875 -46.075 223.205 ;
        RECT -46.405 221.515 -46.075 221.845 ;
        RECT -46.405 220.155 -46.075 220.485 ;
        RECT -46.405 218.795 -46.075 219.125 ;
        RECT -46.405 217.435 -46.075 217.765 ;
        RECT -46.405 216.075 -46.075 216.405 ;
        RECT -46.405 214.715 -46.075 215.045 ;
        RECT -46.405 213.355 -46.075 213.685 ;
        RECT -46.405 211.995 -46.075 212.325 ;
        RECT -46.405 210.635 -46.075 210.965 ;
        RECT -46.405 209.275 -46.075 209.605 ;
        RECT -46.405 207.915 -46.075 208.245 ;
        RECT -46.405 206.555 -46.075 206.885 ;
        RECT -46.405 205.195 -46.075 205.525 ;
        RECT -46.405 203.835 -46.075 204.165 ;
        RECT -46.405 202.475 -46.075 202.805 ;
        RECT -46.405 201.115 -46.075 201.445 ;
        RECT -46.405 199.755 -46.075 200.085 ;
        RECT -46.405 198.395 -46.075 198.725 ;
        RECT -46.405 197.035 -46.075 197.365 ;
        RECT -46.405 195.675 -46.075 196.005 ;
        RECT -46.405 194.315 -46.075 194.645 ;
        RECT -46.405 192.955 -46.075 193.285 ;
        RECT -46.405 191.595 -46.075 191.925 ;
        RECT -46.405 190.235 -46.075 190.565 ;
        RECT -46.405 188.875 -46.075 189.205 ;
        RECT -46.405 187.515 -46.075 187.845 ;
        RECT -46.405 186.155 -46.075 186.485 ;
        RECT -46.405 184.795 -46.075 185.125 ;
        RECT -46.405 183.435 -46.075 183.765 ;
        RECT -46.405 182.075 -46.075 182.405 ;
        RECT -46.405 180.715 -46.075 181.045 ;
        RECT -46.405 179.355 -46.075 179.685 ;
        RECT -46.405 177.995 -46.075 178.325 ;
        RECT -46.405 176.635 -46.075 176.965 ;
        RECT -46.405 175.275 -46.075 175.605 ;
        RECT -46.405 173.915 -46.075 174.245 ;
        RECT -46.405 172.555 -46.075 172.885 ;
        RECT -46.405 171.195 -46.075 171.525 ;
        RECT -46.405 169.835 -46.075 170.165 ;
        RECT -46.405 168.475 -46.075 168.805 ;
        RECT -46.405 167.115 -46.075 167.445 ;
        RECT -46.405 165.755 -46.075 166.085 ;
        RECT -46.405 164.395 -46.075 164.725 ;
        RECT -46.405 163.035 -46.075 163.365 ;
        RECT -46.405 161.675 -46.075 162.005 ;
        RECT -46.405 160.315 -46.075 160.645 ;
        RECT -46.405 158.955 -46.075 159.285 ;
        RECT -46.405 157.595 -46.075 157.925 ;
        RECT -46.405 156.235 -46.075 156.565 ;
        RECT -46.405 154.875 -46.075 155.205 ;
        RECT -46.405 153.515 -46.075 153.845 ;
        RECT -46.405 152.155 -46.075 152.485 ;
        RECT -46.405 150.795 -46.075 151.125 ;
        RECT -46.405 149.435 -46.075 149.765 ;
        RECT -46.405 148.075 -46.075 148.405 ;
        RECT -46.405 146.715 -46.075 147.045 ;
        RECT -46.405 145.355 -46.075 145.685 ;
        RECT -46.405 143.995 -46.075 144.325 ;
        RECT -46.405 142.635 -46.075 142.965 ;
        RECT -46.405 141.275 -46.075 141.605 ;
        RECT -46.405 139.915 -46.075 140.245 ;
        RECT -46.405 138.555 -46.075 138.885 ;
        RECT -46.405 137.195 -46.075 137.525 ;
        RECT -46.405 135.835 -46.075 136.165 ;
        RECT -46.405 134.475 -46.075 134.805 ;
        RECT -46.405 133.115 -46.075 133.445 ;
        RECT -46.405 131.755 -46.075 132.085 ;
        RECT -46.405 130.395 -46.075 130.725 ;
        RECT -46.405 129.035 -46.075 129.365 ;
        RECT -46.405 127.675 -46.075 128.005 ;
        RECT -46.405 126.315 -46.075 126.645 ;
        RECT -46.405 124.955 -46.075 125.285 ;
        RECT -46.405 123.595 -46.075 123.925 ;
        RECT -46.405 122.235 -46.075 122.565 ;
        RECT -46.405 120.875 -46.075 121.205 ;
        RECT -46.405 119.515 -46.075 119.845 ;
        RECT -46.405 118.155 -46.075 118.485 ;
        RECT -46.405 116.795 -46.075 117.125 ;
        RECT -46.405 115.435 -46.075 115.765 ;
        RECT -46.405 114.075 -46.075 114.405 ;
        RECT -46.405 112.715 -46.075 113.045 ;
        RECT -46.405 111.355 -46.075 111.685 ;
        RECT -46.405 109.995 -46.075 110.325 ;
        RECT -46.405 108.635 -46.075 108.965 ;
        RECT -46.405 107.275 -46.075 107.605 ;
        RECT -46.405 105.915 -46.075 106.245 ;
        RECT -46.405 104.555 -46.075 104.885 ;
        RECT -46.405 103.195 -46.075 103.525 ;
        RECT -46.405 101.835 -46.075 102.165 ;
        RECT -46.405 100.475 -46.075 100.805 ;
        RECT -46.405 99.115 -46.075 99.445 ;
        RECT -46.405 97.755 -46.075 98.085 ;
        RECT -46.405 96.395 -46.075 96.725 ;
        RECT -46.405 95.035 -46.075 95.365 ;
        RECT -46.405 93.675 -46.075 94.005 ;
        RECT -46.405 92.315 -46.075 92.645 ;
        RECT -46.405 90.955 -46.075 91.285 ;
        RECT -46.405 89.595 -46.075 89.925 ;
        RECT -46.405 88.235 -46.075 88.565 ;
        RECT -46.405 86.875 -46.075 87.205 ;
        RECT -46.405 85.515 -46.075 85.845 ;
        RECT -46.405 84.155 -46.075 84.485 ;
        RECT -46.405 82.795 -46.075 83.125 ;
        RECT -46.405 81.435 -46.075 81.765 ;
        RECT -46.405 80.075 -46.075 80.405 ;
        RECT -46.405 78.715 -46.075 79.045 ;
        RECT -46.405 77.355 -46.075 77.685 ;
        RECT -46.405 75.995 -46.075 76.325 ;
        RECT -46.405 74.635 -46.075 74.965 ;
        RECT -46.405 73.275 -46.075 73.605 ;
        RECT -46.405 71.915 -46.075 72.245 ;
        RECT -46.405 70.555 -46.075 70.885 ;
        RECT -46.405 69.195 -46.075 69.525 ;
        RECT -46.405 67.835 -46.075 68.165 ;
        RECT -46.405 66.475 -46.075 66.805 ;
        RECT -46.405 65.115 -46.075 65.445 ;
        RECT -46.405 63.755 -46.075 64.085 ;
        RECT -46.405 62.395 -46.075 62.725 ;
        RECT -46.405 61.035 -46.075 61.365 ;
        RECT -46.405 59.675 -46.075 60.005 ;
        RECT -46.405 58.315 -46.075 58.645 ;
        RECT -46.405 56.955 -46.075 57.285 ;
        RECT -46.405 55.595 -46.075 55.925 ;
        RECT -46.405 54.235 -46.075 54.565 ;
        RECT -46.405 52.875 -46.075 53.205 ;
        RECT -46.405 51.515 -46.075 51.845 ;
        RECT -46.405 50.155 -46.075 50.485 ;
        RECT -46.405 48.795 -46.075 49.125 ;
        RECT -46.405 47.435 -46.075 47.765 ;
        RECT -46.405 46.075 -46.075 46.405 ;
        RECT -46.405 44.715 -46.075 45.045 ;
        RECT -46.405 43.355 -46.075 43.685 ;
        RECT -46.405 41.995 -46.075 42.325 ;
        RECT -46.405 40.635 -46.075 40.965 ;
        RECT -46.405 39.275 -46.075 39.605 ;
        RECT -46.405 37.915 -46.075 38.245 ;
        RECT -46.405 36.555 -46.075 36.885 ;
        RECT -46.405 35.195 -46.075 35.525 ;
        RECT -46.405 33.835 -46.075 34.165 ;
        RECT -46.405 32.475 -46.075 32.805 ;
        RECT -46.405 31.115 -46.075 31.445 ;
        RECT -46.405 29.755 -46.075 30.085 ;
        RECT -46.405 28.395 -46.075 28.725 ;
        RECT -46.405 27.035 -46.075 27.365 ;
        RECT -46.405 25.675 -46.075 26.005 ;
        RECT -46.405 24.315 -46.075 24.645 ;
        RECT -46.405 22.955 -46.075 23.285 ;
        RECT -46.405 21.595 -46.075 21.925 ;
        RECT -46.405 20.235 -46.075 20.565 ;
        RECT -46.405 18.875 -46.075 19.205 ;
        RECT -46.405 17.515 -46.075 17.845 ;
        RECT -46.405 16.155 -46.075 16.485 ;
        RECT -46.405 14.795 -46.075 15.125 ;
        RECT -46.405 13.435 -46.075 13.765 ;
        RECT -46.405 12.075 -46.075 12.405 ;
        RECT -46.405 10.715 -46.075 11.045 ;
        RECT -46.405 9.355 -46.075 9.685 ;
        RECT -46.405 7.995 -46.075 8.325 ;
        RECT -46.405 6.635 -46.075 6.965 ;
        RECT -46.405 5.275 -46.075 5.605 ;
        RECT -46.405 3.915 -46.075 4.245 ;
        RECT -46.405 2.555 -46.075 2.885 ;
        RECT -46.405 1.195 -46.075 1.525 ;
        RECT -46.405 -0.165 -46.075 0.165 ;
        RECT -46.4 -1.52 -46.08 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -46.405 -31.445 -46.075 -31.115 ;
        RECT -46.405 -32.805 -46.075 -32.475 ;
        RECT -46.405 -35.525 -46.075 -35.195 ;
        RECT -46.405 -36.885 -46.075 -36.555 ;
        RECT -46.405 -37.93 -46.075 -37.6 ;
        RECT -46.405 -40.965 -46.075 -40.635 ;
        RECT -46.405 -42.77 -46.075 -42.44 ;
        RECT -46.405 -43.685 -46.075 -43.355 ;
        RECT -46.405 -50.485 -46.075 -50.155 ;
        RECT -46.405 -51.845 -46.075 -51.515 ;
        RECT -46.405 -54.565 -46.075 -54.235 ;
        RECT -46.405 -55.925 -46.075 -55.595 ;
        RECT -46.405 -60.005 -46.075 -59.675 ;
        RECT -46.405 -66.805 -46.075 -66.475 ;
        RECT -46.405 -68.165 -46.075 -67.835 ;
        RECT -46.405 -69.525 -46.075 -69.195 ;
        RECT -46.405 -70.885 -46.075 -70.555 ;
        RECT -46.405 -72.245 -46.075 -71.915 ;
        RECT -46.405 -73.605 -46.075 -73.275 ;
        RECT -46.405 -74.965 -46.075 -74.635 ;
        RECT -46.405 -76.325 -46.075 -75.995 ;
        RECT -46.405 -77.685 -46.075 -77.355 ;
        RECT -46.405 -79.045 -46.075 -78.715 ;
        RECT -46.405 -80.405 -46.075 -80.075 ;
        RECT -46.405 -81.765 -46.075 -81.435 ;
        RECT -46.405 -83.125 -46.075 -82.795 ;
        RECT -46.405 -84.485 -46.075 -84.155 ;
        RECT -46.405 -85.845 -46.075 -85.515 ;
        RECT -46.405 -87.205 -46.075 -86.875 ;
        RECT -46.405 -88.565 -46.075 -88.235 ;
        RECT -46.405 -89.925 -46.075 -89.595 ;
        RECT -46.405 -92.645 -46.075 -92.315 ;
        RECT -46.405 -94.005 -46.075 -93.675 ;
        RECT -46.405 -95.365 -46.075 -95.035 ;
        RECT -46.405 -96.725 -46.075 -96.395 ;
        RECT -46.405 -98.73 -46.075 -98.4 ;
        RECT -46.405 -99.445 -46.075 -99.115 ;
        RECT -46.405 -102.165 -46.075 -101.835 ;
        RECT -46.405 -103.525 -46.075 -103.195 ;
        RECT -46.405 -104.885 -46.075 -104.555 ;
        RECT -46.405 -106.87 -46.075 -106.54 ;
        RECT -46.405 -107.605 -46.075 -107.275 ;
        RECT -46.405 -108.965 -46.075 -108.635 ;
        RECT -46.4 -111.68 -46.08 -29.08 ;
    END
    PORT
      LAYER met3 ;
        RECT -45.045 237.835 -44.715 238.165 ;
        RECT -45.045 236.475 -44.715 236.805 ;
        RECT -45.045 235.115 -44.715 235.445 ;
        RECT -45.045 233.755 -44.715 234.085 ;
        RECT -45.045 232.395 -44.715 232.725 ;
        RECT -45.045 231.035 -44.715 231.365 ;
        RECT -45.045 229.675 -44.715 230.005 ;
        RECT -45.045 228.315 -44.715 228.645 ;
        RECT -45.045 226.955 -44.715 227.285 ;
        RECT -45.045 225.595 -44.715 225.925 ;
        RECT -45.045 224.235 -44.715 224.565 ;
        RECT -45.045 222.875 -44.715 223.205 ;
        RECT -45.045 221.515 -44.715 221.845 ;
        RECT -45.045 220.155 -44.715 220.485 ;
        RECT -45.045 218.795 -44.715 219.125 ;
        RECT -45.045 217.435 -44.715 217.765 ;
        RECT -45.045 216.075 -44.715 216.405 ;
        RECT -45.045 214.715 -44.715 215.045 ;
        RECT -45.045 213.355 -44.715 213.685 ;
        RECT -45.045 211.995 -44.715 212.325 ;
        RECT -45.045 210.635 -44.715 210.965 ;
        RECT -45.045 209.275 -44.715 209.605 ;
        RECT -45.045 207.915 -44.715 208.245 ;
        RECT -45.045 206.555 -44.715 206.885 ;
        RECT -45.045 205.195 -44.715 205.525 ;
        RECT -45.045 203.835 -44.715 204.165 ;
        RECT -45.045 202.475 -44.715 202.805 ;
        RECT -45.045 201.115 -44.715 201.445 ;
        RECT -45.045 199.755 -44.715 200.085 ;
        RECT -45.045 198.395 -44.715 198.725 ;
        RECT -45.045 197.035 -44.715 197.365 ;
        RECT -45.045 195.675 -44.715 196.005 ;
        RECT -45.045 194.315 -44.715 194.645 ;
        RECT -45.045 192.955 -44.715 193.285 ;
        RECT -45.045 191.595 -44.715 191.925 ;
        RECT -45.045 190.235 -44.715 190.565 ;
        RECT -45.045 188.875 -44.715 189.205 ;
        RECT -45.045 187.515 -44.715 187.845 ;
        RECT -45.045 186.155 -44.715 186.485 ;
        RECT -45.045 184.795 -44.715 185.125 ;
        RECT -45.045 183.435 -44.715 183.765 ;
        RECT -45.045 182.075 -44.715 182.405 ;
        RECT -45.045 180.715 -44.715 181.045 ;
        RECT -45.045 179.355 -44.715 179.685 ;
        RECT -45.045 177.995 -44.715 178.325 ;
        RECT -45.045 176.635 -44.715 176.965 ;
        RECT -45.045 175.275 -44.715 175.605 ;
        RECT -45.045 173.915 -44.715 174.245 ;
        RECT -45.045 172.555 -44.715 172.885 ;
        RECT -45.045 171.195 -44.715 171.525 ;
        RECT -45.045 169.835 -44.715 170.165 ;
        RECT -45.045 168.475 -44.715 168.805 ;
        RECT -45.045 167.115 -44.715 167.445 ;
        RECT -45.045 165.755 -44.715 166.085 ;
        RECT -45.045 164.395 -44.715 164.725 ;
        RECT -45.045 163.035 -44.715 163.365 ;
        RECT -45.045 161.675 -44.715 162.005 ;
        RECT -45.045 160.315 -44.715 160.645 ;
        RECT -45.045 158.955 -44.715 159.285 ;
        RECT -45.045 157.595 -44.715 157.925 ;
        RECT -45.045 156.235 -44.715 156.565 ;
        RECT -45.045 154.875 -44.715 155.205 ;
        RECT -45.045 153.515 -44.715 153.845 ;
        RECT -45.045 152.155 -44.715 152.485 ;
        RECT -45.045 150.795 -44.715 151.125 ;
        RECT -45.045 149.435 -44.715 149.765 ;
        RECT -45.045 148.075 -44.715 148.405 ;
        RECT -45.045 146.715 -44.715 147.045 ;
        RECT -45.045 145.355 -44.715 145.685 ;
        RECT -45.045 143.995 -44.715 144.325 ;
        RECT -45.045 142.635 -44.715 142.965 ;
        RECT -45.045 141.275 -44.715 141.605 ;
        RECT -45.045 139.915 -44.715 140.245 ;
        RECT -45.045 138.555 -44.715 138.885 ;
        RECT -45.045 137.195 -44.715 137.525 ;
        RECT -45.045 135.835 -44.715 136.165 ;
        RECT -45.045 134.475 -44.715 134.805 ;
        RECT -45.045 133.115 -44.715 133.445 ;
        RECT -45.045 131.755 -44.715 132.085 ;
        RECT -45.045 130.395 -44.715 130.725 ;
        RECT -45.045 129.035 -44.715 129.365 ;
        RECT -45.045 127.675 -44.715 128.005 ;
        RECT -45.045 126.315 -44.715 126.645 ;
        RECT -45.045 124.955 -44.715 125.285 ;
        RECT -45.045 123.595 -44.715 123.925 ;
        RECT -45.045 122.235 -44.715 122.565 ;
        RECT -45.045 120.875 -44.715 121.205 ;
        RECT -45.045 119.515 -44.715 119.845 ;
        RECT -45.045 118.155 -44.715 118.485 ;
        RECT -45.045 116.795 -44.715 117.125 ;
        RECT -45.045 115.435 -44.715 115.765 ;
        RECT -45.045 114.075 -44.715 114.405 ;
        RECT -45.045 112.715 -44.715 113.045 ;
        RECT -45.045 111.355 -44.715 111.685 ;
        RECT -45.045 109.995 -44.715 110.325 ;
        RECT -45.045 108.635 -44.715 108.965 ;
        RECT -45.045 107.275 -44.715 107.605 ;
        RECT -45.045 105.915 -44.715 106.245 ;
        RECT -45.045 104.555 -44.715 104.885 ;
        RECT -45.045 103.195 -44.715 103.525 ;
        RECT -45.045 101.835 -44.715 102.165 ;
        RECT -45.045 100.475 -44.715 100.805 ;
        RECT -45.045 99.115 -44.715 99.445 ;
        RECT -45.045 97.755 -44.715 98.085 ;
        RECT -45.045 96.395 -44.715 96.725 ;
        RECT -45.045 95.035 -44.715 95.365 ;
        RECT -45.045 93.675 -44.715 94.005 ;
        RECT -45.045 92.315 -44.715 92.645 ;
        RECT -45.045 90.955 -44.715 91.285 ;
        RECT -45.045 89.595 -44.715 89.925 ;
        RECT -45.045 88.235 -44.715 88.565 ;
        RECT -45.045 86.875 -44.715 87.205 ;
        RECT -45.045 85.515 -44.715 85.845 ;
        RECT -45.045 84.155 -44.715 84.485 ;
        RECT -45.045 82.795 -44.715 83.125 ;
        RECT -45.045 81.435 -44.715 81.765 ;
        RECT -45.045 80.075 -44.715 80.405 ;
        RECT -45.045 78.715 -44.715 79.045 ;
        RECT -45.045 77.355 -44.715 77.685 ;
        RECT -45.045 75.995 -44.715 76.325 ;
        RECT -45.045 74.635 -44.715 74.965 ;
        RECT -45.045 73.275 -44.715 73.605 ;
        RECT -45.045 71.915 -44.715 72.245 ;
        RECT -45.045 70.555 -44.715 70.885 ;
        RECT -45.045 69.195 -44.715 69.525 ;
        RECT -45.045 67.835 -44.715 68.165 ;
        RECT -45.045 66.475 -44.715 66.805 ;
        RECT -45.045 65.115 -44.715 65.445 ;
        RECT -45.045 63.755 -44.715 64.085 ;
        RECT -45.045 62.395 -44.715 62.725 ;
        RECT -45.045 61.035 -44.715 61.365 ;
        RECT -45.045 59.675 -44.715 60.005 ;
        RECT -45.045 58.315 -44.715 58.645 ;
        RECT -45.045 56.955 -44.715 57.285 ;
        RECT -45.045 55.595 -44.715 55.925 ;
        RECT -45.045 54.235 -44.715 54.565 ;
        RECT -45.045 52.875 -44.715 53.205 ;
        RECT -45.045 51.515 -44.715 51.845 ;
        RECT -45.045 50.155 -44.715 50.485 ;
        RECT -45.045 48.795 -44.715 49.125 ;
        RECT -45.045 47.435 -44.715 47.765 ;
        RECT -45.045 46.075 -44.715 46.405 ;
        RECT -45.045 44.715 -44.715 45.045 ;
        RECT -45.045 43.355 -44.715 43.685 ;
        RECT -45.045 41.995 -44.715 42.325 ;
        RECT -45.045 40.635 -44.715 40.965 ;
        RECT -45.045 39.275 -44.715 39.605 ;
        RECT -45.045 37.915 -44.715 38.245 ;
        RECT -45.045 36.555 -44.715 36.885 ;
        RECT -45.045 35.195 -44.715 35.525 ;
        RECT -45.045 33.835 -44.715 34.165 ;
        RECT -45.045 32.475 -44.715 32.805 ;
        RECT -45.045 31.115 -44.715 31.445 ;
        RECT -45.045 29.755 -44.715 30.085 ;
        RECT -45.045 28.395 -44.715 28.725 ;
        RECT -45.045 27.035 -44.715 27.365 ;
        RECT -45.045 25.675 -44.715 26.005 ;
        RECT -45.045 24.315 -44.715 24.645 ;
        RECT -45.045 22.955 -44.715 23.285 ;
        RECT -45.045 21.595 -44.715 21.925 ;
        RECT -45.045 20.235 -44.715 20.565 ;
        RECT -45.045 18.875 -44.715 19.205 ;
        RECT -45.045 17.515 -44.715 17.845 ;
        RECT -45.045 16.155 -44.715 16.485 ;
        RECT -45.045 14.795 -44.715 15.125 ;
        RECT -45.045 13.435 -44.715 13.765 ;
        RECT -45.045 12.075 -44.715 12.405 ;
        RECT -45.045 10.715 -44.715 11.045 ;
        RECT -45.045 9.355 -44.715 9.685 ;
        RECT -45.045 7.995 -44.715 8.325 ;
        RECT -45.045 6.635 -44.715 6.965 ;
        RECT -45.045 5.275 -44.715 5.605 ;
        RECT -45.045 3.915 -44.715 4.245 ;
        RECT -45.045 2.555 -44.715 2.885 ;
        RECT -45.045 1.195 -44.715 1.525 ;
        RECT -45.045 -0.165 -44.715 0.165 ;
        RECT -45.045 -4.245 -44.715 -3.915 ;
        RECT -45.045 -5.605 -44.715 -5.275 ;
        RECT -45.045 -6.965 -44.715 -6.635 ;
        RECT -45.045 -8.325 -44.715 -7.995 ;
        RECT -45.045 -11.045 -44.715 -10.715 ;
        RECT -45.045 -15.125 -44.715 -14.795 ;
        RECT -45.045 -16.485 -44.715 -16.155 ;
        RECT -45.045 -17.845 -44.715 -17.515 ;
        RECT -45.045 -19.205 -44.715 -18.875 ;
        RECT -45.045 -20.565 -44.715 -20.235 ;
        RECT -45.045 -21.925 -44.715 -21.595 ;
        RECT -45.045 -23.285 -44.715 -22.955 ;
        RECT -45.045 -24.645 -44.715 -24.315 ;
        RECT -45.045 -31.445 -44.715 -31.115 ;
        RECT -45.045 -32.805 -44.715 -32.475 ;
        RECT -45.045 -35.525 -44.715 -35.195 ;
        RECT -45.045 -36.885 -44.715 -36.555 ;
        RECT -45.045 -37.93 -44.715 -37.6 ;
        RECT -45.045 -40.965 -44.715 -40.635 ;
        RECT -45.045 -42.77 -44.715 -42.44 ;
        RECT -45.045 -43.685 -44.715 -43.355 ;
        RECT -45.045 -50.485 -44.715 -50.155 ;
        RECT -45.045 -51.845 -44.715 -51.515 ;
        RECT -45.045 -54.565 -44.715 -54.235 ;
        RECT -45.045 -55.925 -44.715 -55.595 ;
        RECT -45.045 -60.005 -44.715 -59.675 ;
        RECT -45.04 -64.76 -44.72 242.565 ;
        RECT -45.045 241.32 -44.715 242.45 ;
        RECT -45.045 239.195 -44.715 239.525 ;
    END
    PORT
      LAYER met3 ;
        RECT -54.565 97.755 -54.235 98.085 ;
        RECT -54.565 96.395 -54.235 96.725 ;
        RECT -54.565 95.035 -54.235 95.365 ;
        RECT -54.565 93.675 -54.235 94.005 ;
        RECT -54.565 92.315 -54.235 92.645 ;
        RECT -54.565 89.595 -54.235 89.925 ;
        RECT -54.565 88.235 -54.235 88.565 ;
        RECT -54.565 84.155 -54.235 84.485 ;
        RECT -54.565 82.795 -54.235 83.125 ;
        RECT -54.565 81.435 -54.235 81.765 ;
        RECT -54.565 80.075 -54.235 80.405 ;
        RECT -54.565 78.715 -54.235 79.045 ;
        RECT -54.565 77.355 -54.235 77.685 ;
        RECT -54.565 75.995 -54.235 76.325 ;
        RECT -54.565 74.635 -54.235 74.965 ;
        RECT -54.565 73.275 -54.235 73.605 ;
        RECT -54.565 71.915 -54.235 72.245 ;
        RECT -54.565 70.555 -54.235 70.885 ;
        RECT -54.565 69.195 -54.235 69.525 ;
        RECT -54.565 67.835 -54.235 68.165 ;
        RECT -54.565 66.475 -54.235 66.805 ;
        RECT -54.565 65.115 -54.235 65.445 ;
        RECT -54.565 63.755 -54.235 64.085 ;
        RECT -54.565 62.395 -54.235 62.725 ;
        RECT -54.565 61.035 -54.235 61.365 ;
        RECT -54.565 59.675 -54.235 60.005 ;
        RECT -54.565 58.315 -54.235 58.645 ;
        RECT -54.565 56.955 -54.235 57.285 ;
        RECT -54.565 55.595 -54.235 55.925 ;
        RECT -54.565 54.235 -54.235 54.565 ;
        RECT -54.565 52.875 -54.235 53.205 ;
        RECT -54.565 51.515 -54.235 51.845 ;
        RECT -54.565 50.155 -54.235 50.485 ;
        RECT -54.565 48.795 -54.235 49.125 ;
        RECT -54.565 47.435 -54.235 47.765 ;
        RECT -54.565 46.075 -54.235 46.405 ;
        RECT -54.565 44.715 -54.235 45.045 ;
        RECT -54.565 43.355 -54.235 43.685 ;
        RECT -54.565 41.995 -54.235 42.325 ;
        RECT -54.565 40.635 -54.235 40.965 ;
        RECT -54.565 39.275 -54.235 39.605 ;
        RECT -54.565 37.915 -54.235 38.245 ;
        RECT -54.565 36.555 -54.235 36.885 ;
        RECT -54.565 35.195 -54.235 35.525 ;
        RECT -54.565 33.835 -54.235 34.165 ;
        RECT -54.565 32.475 -54.235 32.805 ;
        RECT -54.565 31.115 -54.235 31.445 ;
        RECT -54.565 29.755 -54.235 30.085 ;
        RECT -54.565 28.395 -54.235 28.725 ;
        RECT -54.565 27.035 -54.235 27.365 ;
        RECT -54.565 25.675 -54.235 26.005 ;
        RECT -54.565 24.315 -54.235 24.645 ;
        RECT -54.565 22.955 -54.235 23.285 ;
        RECT -54.565 21.595 -54.235 21.925 ;
        RECT -54.565 20.235 -54.235 20.565 ;
        RECT -54.565 18.875 -54.235 19.205 ;
        RECT -54.565 17.515 -54.235 17.845 ;
        RECT -54.565 16.155 -54.235 16.485 ;
        RECT -54.565 14.795 -54.235 15.125 ;
        RECT -54.565 13.435 -54.235 13.765 ;
        RECT -54.565 12.075 -54.235 12.405 ;
        RECT -54.565 10.715 -54.235 11.045 ;
        RECT -54.565 9.355 -54.235 9.685 ;
        RECT -54.565 7.995 -54.235 8.325 ;
        RECT -54.565 6.635 -54.235 6.965 ;
        RECT -54.565 5.275 -54.235 5.605 ;
        RECT -54.565 3.915 -54.235 4.245 ;
        RECT -54.565 2.555 -54.235 2.885 ;
        RECT -54.565 1.195 -54.235 1.525 ;
        RECT -54.565 -0.165 -54.235 0.165 ;
        RECT -54.565 -2.885 -54.235 -2.555 ;
        RECT -54.565 -4.245 -54.235 -3.915 ;
        RECT -54.565 -5.605 -54.235 -5.275 ;
        RECT -54.565 -6.965 -54.235 -6.635 ;
        RECT -54.565 -8.325 -54.235 -7.995 ;
        RECT -54.565 -9.685 -54.235 -9.355 ;
        RECT -54.565 -11.045 -54.235 -10.715 ;
        RECT -54.565 -12.405 -54.235 -12.075 ;
        RECT -54.565 -13.765 -54.235 -13.435 ;
        RECT -54.565 -15.125 -54.235 -14.795 ;
        RECT -54.565 -16.485 -54.235 -16.155 ;
        RECT -54.565 -17.845 -54.235 -17.515 ;
        RECT -54.565 -19.205 -54.235 -18.875 ;
        RECT -54.565 -20.565 -54.235 -20.235 ;
        RECT -54.565 -21.925 -54.235 -21.595 ;
        RECT -54.565 -23.285 -54.235 -22.955 ;
        RECT -54.565 -24.645 -54.235 -24.315 ;
        RECT -54.565 -27.365 -54.235 -27.035 ;
        RECT -54.565 -28.725 -54.235 -28.395 ;
        RECT -54.565 -30.085 -54.235 -29.755 ;
        RECT -54.565 -31.445 -54.235 -31.115 ;
        RECT -54.565 -32.805 -54.235 -32.475 ;
        RECT -54.565 -34.165 -54.235 -33.835 ;
        RECT -54.565 -35.525 -54.235 -35.195 ;
        RECT -54.565 -36.885 -54.235 -36.555 ;
        RECT -54.565 -38.245 -54.235 -37.915 ;
        RECT -54.565 -39.605 -54.235 -39.275 ;
        RECT -54.565 -40.965 -54.235 -40.635 ;
        RECT -54.565 -42.325 -54.235 -41.995 ;
        RECT -54.565 -43.685 -54.235 -43.355 ;
        RECT -54.565 -45.045 -54.235 -44.715 ;
        RECT -54.565 -46.405 -54.235 -46.075 ;
        RECT -54.565 -47.765 -54.235 -47.435 ;
        RECT -54.565 -49.125 -54.235 -48.795 ;
        RECT -54.565 -50.485 -54.235 -50.155 ;
        RECT -54.565 -51.845 -54.235 -51.515 ;
        RECT -54.565 -53.205 -54.235 -52.875 ;
        RECT -54.565 -54.565 -54.235 -54.235 ;
        RECT -54.565 -55.925 -54.235 -55.595 ;
        RECT -54.565 -57.285 -54.235 -56.955 ;
        RECT -54.565 -58.645 -54.235 -58.315 ;
        RECT -54.565 -60.005 -54.235 -59.675 ;
        RECT -54.565 -61.365 -54.235 -61.035 ;
        RECT -54.565 -62.725 -54.235 -62.395 ;
        RECT -54.565 -64.085 -54.235 -63.755 ;
        RECT -54.565 -65.445 -54.235 -65.115 ;
        RECT -54.565 -66.805 -54.235 -66.475 ;
        RECT -54.565 -68.165 -54.235 -67.835 ;
        RECT -54.565 -69.525 -54.235 -69.195 ;
        RECT -54.565 -70.885 -54.235 -70.555 ;
        RECT -54.565 -72.245 -54.235 -71.915 ;
        RECT -54.565 -73.605 -54.235 -73.275 ;
        RECT -54.565 -74.965 -54.235 -74.635 ;
        RECT -54.565 -76.325 -54.235 -75.995 ;
        RECT -54.565 -77.685 -54.235 -77.355 ;
        RECT -54.565 -79.045 -54.235 -78.715 ;
        RECT -54.565 -80.405 -54.235 -80.075 ;
        RECT -54.565 -81.765 -54.235 -81.435 ;
        RECT -54.565 -83.125 -54.235 -82.795 ;
        RECT -54.565 -84.485 -54.235 -84.155 ;
        RECT -54.565 -85.845 -54.235 -85.515 ;
        RECT -54.565 -87.205 -54.235 -86.875 ;
        RECT -54.565 -88.565 -54.235 -88.235 ;
        RECT -54.565 -89.925 -54.235 -89.595 ;
        RECT -54.565 -92.645 -54.235 -92.315 ;
        RECT -54.565 -94.005 -54.235 -93.675 ;
        RECT -54.565 -95.365 -54.235 -95.035 ;
        RECT -54.565 -96.725 -54.235 -96.395 ;
        RECT -54.565 -98.73 -54.235 -98.4 ;
        RECT -54.565 -99.445 -54.235 -99.115 ;
        RECT -54.565 -102.165 -54.235 -101.835 ;
        RECT -54.565 -103.525 -54.235 -103.195 ;
        RECT -54.565 -104.885 -54.235 -104.555 ;
        RECT -54.565 -106.87 -54.235 -106.54 ;
        RECT -54.565 -107.605 -54.235 -107.275 ;
        RECT -54.565 -108.965 -54.235 -108.635 ;
        RECT -54.565 -110.325 -54.235 -109.995 ;
        RECT -54.56 -112.36 -54.24 98.085 ;
    END
    PORT
      LAYER met3 ;
        RECT -54.565 -174.245 -54.235 -173.915 ;
        RECT -54.565 -175.725 -54.235 -175.395 ;
        RECT -54.565 -176.965 -54.235 -176.635 ;
        RECT -54.565 -178.325 -54.235 -177.995 ;
        RECT -54.565 -180.57 -54.235 -179.44 ;
        RECT -54.56 -180.685 -54.24 -173.915 ;
    END
    PORT
      LAYER met3 ;
        RECT -53.205 241.32 -52.875 242.45 ;
        RECT -53.205 239.195 -52.875 239.525 ;
        RECT -53.205 237.835 -52.875 238.165 ;
        RECT -53.205 236.475 -52.875 236.805 ;
        RECT -53.205 235.115 -52.875 235.445 ;
        RECT -53.205 233.755 -52.875 234.085 ;
        RECT -53.205 232.395 -52.875 232.725 ;
        RECT -53.205 231.035 -52.875 231.365 ;
        RECT -53.205 229.675 -52.875 230.005 ;
        RECT -53.205 228.315 -52.875 228.645 ;
        RECT -53.205 226.955 -52.875 227.285 ;
        RECT -53.205 225.595 -52.875 225.925 ;
        RECT -53.205 224.235 -52.875 224.565 ;
        RECT -53.205 222.875 -52.875 223.205 ;
        RECT -53.205 221.515 -52.875 221.845 ;
        RECT -53.205 220.155 -52.875 220.485 ;
        RECT -53.205 218.795 -52.875 219.125 ;
        RECT -53.205 217.435 -52.875 217.765 ;
        RECT -53.205 216.075 -52.875 216.405 ;
        RECT -53.205 214.715 -52.875 215.045 ;
        RECT -53.205 213.355 -52.875 213.685 ;
        RECT -53.205 211.995 -52.875 212.325 ;
        RECT -53.205 210.635 -52.875 210.965 ;
        RECT -53.205 209.275 -52.875 209.605 ;
        RECT -53.205 207.915 -52.875 208.245 ;
        RECT -53.205 206.555 -52.875 206.885 ;
        RECT -53.205 205.195 -52.875 205.525 ;
        RECT -53.205 203.835 -52.875 204.165 ;
        RECT -53.205 202.475 -52.875 202.805 ;
        RECT -53.205 201.115 -52.875 201.445 ;
        RECT -53.205 199.755 -52.875 200.085 ;
        RECT -53.205 198.395 -52.875 198.725 ;
        RECT -53.205 197.035 -52.875 197.365 ;
        RECT -53.205 195.675 -52.875 196.005 ;
        RECT -53.205 194.315 -52.875 194.645 ;
        RECT -53.205 192.955 -52.875 193.285 ;
        RECT -53.205 191.595 -52.875 191.925 ;
        RECT -53.205 190.235 -52.875 190.565 ;
        RECT -53.205 188.875 -52.875 189.205 ;
        RECT -53.205 187.515 -52.875 187.845 ;
        RECT -53.205 186.155 -52.875 186.485 ;
        RECT -53.205 184.795 -52.875 185.125 ;
        RECT -53.205 183.435 -52.875 183.765 ;
        RECT -53.205 182.075 -52.875 182.405 ;
        RECT -53.205 180.715 -52.875 181.045 ;
        RECT -53.205 179.355 -52.875 179.685 ;
        RECT -53.205 177.995 -52.875 178.325 ;
        RECT -53.205 176.635 -52.875 176.965 ;
        RECT -53.205 175.275 -52.875 175.605 ;
        RECT -53.205 173.915 -52.875 174.245 ;
        RECT -53.205 172.555 -52.875 172.885 ;
        RECT -53.205 171.195 -52.875 171.525 ;
        RECT -53.205 169.835 -52.875 170.165 ;
        RECT -53.205 168.475 -52.875 168.805 ;
        RECT -53.205 167.115 -52.875 167.445 ;
        RECT -53.205 165.755 -52.875 166.085 ;
        RECT -53.205 164.395 -52.875 164.725 ;
        RECT -53.205 163.035 -52.875 163.365 ;
        RECT -53.205 161.675 -52.875 162.005 ;
        RECT -53.205 160.315 -52.875 160.645 ;
        RECT -53.205 158.955 -52.875 159.285 ;
        RECT -53.205 157.595 -52.875 157.925 ;
        RECT -53.205 156.235 -52.875 156.565 ;
        RECT -53.205 154.875 -52.875 155.205 ;
        RECT -53.205 153.515 -52.875 153.845 ;
        RECT -53.205 152.155 -52.875 152.485 ;
        RECT -53.205 150.795 -52.875 151.125 ;
        RECT -53.205 149.435 -52.875 149.765 ;
        RECT -53.205 148.075 -52.875 148.405 ;
        RECT -53.205 146.715 -52.875 147.045 ;
        RECT -53.205 145.355 -52.875 145.685 ;
        RECT -53.205 143.995 -52.875 144.325 ;
        RECT -53.205 142.635 -52.875 142.965 ;
        RECT -53.205 141.275 -52.875 141.605 ;
        RECT -53.205 139.915 -52.875 140.245 ;
        RECT -53.205 138.555 -52.875 138.885 ;
        RECT -53.2 138.555 -52.88 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -53.205 97.755 -52.875 98.085 ;
        RECT -53.205 96.395 -52.875 96.725 ;
        RECT -53.205 95.035 -52.875 95.365 ;
        RECT -53.205 93.675 -52.875 94.005 ;
        RECT -53.205 92.315 -52.875 92.645 ;
        RECT -53.205 89.595 -52.875 89.925 ;
        RECT -53.205 88.235 -52.875 88.565 ;
        RECT -53.205 84.155 -52.875 84.485 ;
        RECT -53.205 82.795 -52.875 83.125 ;
        RECT -53.205 81.435 -52.875 81.765 ;
        RECT -53.205 80.075 -52.875 80.405 ;
        RECT -53.205 78.715 -52.875 79.045 ;
        RECT -53.205 77.355 -52.875 77.685 ;
        RECT -53.205 75.995 -52.875 76.325 ;
        RECT -53.205 74.635 -52.875 74.965 ;
        RECT -53.205 73.275 -52.875 73.605 ;
        RECT -53.205 71.915 -52.875 72.245 ;
        RECT -53.205 70.555 -52.875 70.885 ;
        RECT -53.205 69.195 -52.875 69.525 ;
        RECT -53.205 67.835 -52.875 68.165 ;
        RECT -53.205 66.475 -52.875 66.805 ;
        RECT -53.205 65.115 -52.875 65.445 ;
        RECT -53.205 63.755 -52.875 64.085 ;
        RECT -53.205 62.395 -52.875 62.725 ;
        RECT -53.205 61.035 -52.875 61.365 ;
        RECT -53.205 59.675 -52.875 60.005 ;
        RECT -53.205 58.315 -52.875 58.645 ;
        RECT -53.205 56.955 -52.875 57.285 ;
        RECT -53.205 55.595 -52.875 55.925 ;
        RECT -53.205 54.235 -52.875 54.565 ;
        RECT -53.205 52.875 -52.875 53.205 ;
        RECT -53.205 51.515 -52.875 51.845 ;
        RECT -53.205 50.155 -52.875 50.485 ;
        RECT -53.205 48.795 -52.875 49.125 ;
        RECT -53.205 47.435 -52.875 47.765 ;
        RECT -53.205 46.075 -52.875 46.405 ;
        RECT -53.205 44.715 -52.875 45.045 ;
        RECT -53.205 43.355 -52.875 43.685 ;
        RECT -53.205 41.995 -52.875 42.325 ;
        RECT -53.205 40.635 -52.875 40.965 ;
        RECT -53.205 39.275 -52.875 39.605 ;
        RECT -53.205 37.915 -52.875 38.245 ;
        RECT -53.205 36.555 -52.875 36.885 ;
        RECT -53.205 35.195 -52.875 35.525 ;
        RECT -53.205 33.835 -52.875 34.165 ;
        RECT -53.205 32.475 -52.875 32.805 ;
        RECT -53.205 31.115 -52.875 31.445 ;
        RECT -53.205 29.755 -52.875 30.085 ;
        RECT -53.205 28.395 -52.875 28.725 ;
        RECT -53.205 27.035 -52.875 27.365 ;
        RECT -53.205 25.675 -52.875 26.005 ;
        RECT -53.205 24.315 -52.875 24.645 ;
        RECT -53.205 22.955 -52.875 23.285 ;
        RECT -53.205 21.595 -52.875 21.925 ;
        RECT -53.205 20.235 -52.875 20.565 ;
        RECT -53.205 18.875 -52.875 19.205 ;
        RECT -53.205 17.515 -52.875 17.845 ;
        RECT -53.205 16.155 -52.875 16.485 ;
        RECT -53.205 14.795 -52.875 15.125 ;
        RECT -53.205 13.435 -52.875 13.765 ;
        RECT -53.205 12.075 -52.875 12.405 ;
        RECT -53.205 10.715 -52.875 11.045 ;
        RECT -53.205 9.355 -52.875 9.685 ;
        RECT -53.205 7.995 -52.875 8.325 ;
        RECT -53.205 6.635 -52.875 6.965 ;
        RECT -53.205 5.275 -52.875 5.605 ;
        RECT -53.205 3.915 -52.875 4.245 ;
        RECT -53.205 2.555 -52.875 2.885 ;
        RECT -53.205 1.195 -52.875 1.525 ;
        RECT -53.205 -0.165 -52.875 0.165 ;
        RECT -53.205 -2.885 -52.875 -2.555 ;
        RECT -53.205 -4.245 -52.875 -3.915 ;
        RECT -53.205 -5.605 -52.875 -5.275 ;
        RECT -53.205 -6.965 -52.875 -6.635 ;
        RECT -53.205 -8.325 -52.875 -7.995 ;
        RECT -53.205 -9.685 -52.875 -9.355 ;
        RECT -53.205 -11.045 -52.875 -10.715 ;
        RECT -53.205 -12.405 -52.875 -12.075 ;
        RECT -53.205 -13.765 -52.875 -13.435 ;
        RECT -53.205 -15.125 -52.875 -14.795 ;
        RECT -53.205 -16.485 -52.875 -16.155 ;
        RECT -53.205 -17.845 -52.875 -17.515 ;
        RECT -53.205 -19.205 -52.875 -18.875 ;
        RECT -53.205 -20.565 -52.875 -20.235 ;
        RECT -53.205 -21.925 -52.875 -21.595 ;
        RECT -53.205 -23.285 -52.875 -22.955 ;
        RECT -53.205 -24.645 -52.875 -24.315 ;
        RECT -53.205 -28.725 -52.875 -28.395 ;
        RECT -53.205 -30.085 -52.875 -29.755 ;
        RECT -53.205 -31.445 -52.875 -31.115 ;
        RECT -53.205 -32.805 -52.875 -32.475 ;
        RECT -53.205 -34.165 -52.875 -33.835 ;
        RECT -53.205 -35.525 -52.875 -35.195 ;
        RECT -53.205 -36.885 -52.875 -36.555 ;
        RECT -53.205 -38.245 -52.875 -37.915 ;
        RECT -53.205 -39.605 -52.875 -39.275 ;
        RECT -53.205 -40.965 -52.875 -40.635 ;
        RECT -53.205 -42.325 -52.875 -41.995 ;
        RECT -53.205 -43.685 -52.875 -43.355 ;
        RECT -53.205 -45.045 -52.875 -44.715 ;
        RECT -53.205 -46.405 -52.875 -46.075 ;
        RECT -53.205 -47.765 -52.875 -47.435 ;
        RECT -53.205 -49.125 -52.875 -48.795 ;
        RECT -53.205 -50.485 -52.875 -50.155 ;
        RECT -53.205 -51.845 -52.875 -51.515 ;
        RECT -53.205 -53.205 -52.875 -52.875 ;
        RECT -53.205 -54.565 -52.875 -54.235 ;
        RECT -53.205 -55.925 -52.875 -55.595 ;
        RECT -53.205 -57.285 -52.875 -56.955 ;
        RECT -53.205 -58.645 -52.875 -58.315 ;
        RECT -53.205 -60.005 -52.875 -59.675 ;
        RECT -53.205 -61.365 -52.875 -61.035 ;
        RECT -53.205 -62.725 -52.875 -62.395 ;
        RECT -53.205 -64.085 -52.875 -63.755 ;
        RECT -53.205 -65.445 -52.875 -65.115 ;
        RECT -53.205 -66.805 -52.875 -66.475 ;
        RECT -53.205 -68.165 -52.875 -67.835 ;
        RECT -53.205 -69.525 -52.875 -69.195 ;
        RECT -53.205 -70.885 -52.875 -70.555 ;
        RECT -53.205 -72.245 -52.875 -71.915 ;
        RECT -53.205 -73.605 -52.875 -73.275 ;
        RECT -53.205 -74.965 -52.875 -74.635 ;
        RECT -53.205 -76.325 -52.875 -75.995 ;
        RECT -53.205 -77.685 -52.875 -77.355 ;
        RECT -53.205 -79.045 -52.875 -78.715 ;
        RECT -53.205 -80.405 -52.875 -80.075 ;
        RECT -53.205 -81.765 -52.875 -81.435 ;
        RECT -53.205 -83.125 -52.875 -82.795 ;
        RECT -53.205 -84.485 -52.875 -84.155 ;
        RECT -53.205 -85.845 -52.875 -85.515 ;
        RECT -53.205 -87.205 -52.875 -86.875 ;
        RECT -53.205 -88.565 -52.875 -88.235 ;
        RECT -53.205 -89.925 -52.875 -89.595 ;
        RECT -53.205 -92.645 -52.875 -92.315 ;
        RECT -53.205 -94.005 -52.875 -93.675 ;
        RECT -53.205 -95.365 -52.875 -95.035 ;
        RECT -53.205 -96.725 -52.875 -96.395 ;
        RECT -53.205 -98.73 -52.875 -98.4 ;
        RECT -53.205 -99.445 -52.875 -99.115 ;
        RECT -53.205 -102.165 -52.875 -101.835 ;
        RECT -53.205 -103.525 -52.875 -103.195 ;
        RECT -53.205 -104.885 -52.875 -104.555 ;
        RECT -53.205 -106.87 -52.875 -106.54 ;
        RECT -53.205 -107.605 -52.875 -107.275 ;
        RECT -53.205 -108.965 -52.875 -108.635 ;
        RECT -53.205 -110.325 -52.875 -109.995 ;
        RECT -53.205 -115.765 -52.875 -115.435 ;
        RECT -53.205 -117.125 -52.875 -116.795 ;
        RECT -53.205 -118.485 -52.875 -118.155 ;
        RECT -53.205 -122.565 -52.875 -122.235 ;
        RECT -53.205 -123.925 -52.875 -123.595 ;
        RECT -53.205 -125.285 -52.875 -124.955 ;
        RECT -53.205 -126.645 -52.875 -126.315 ;
        RECT -53.205 -128.005 -52.875 -127.675 ;
        RECT -53.205 -129.365 -52.875 -129.035 ;
        RECT -53.205 -130.725 -52.875 -130.395 ;
        RECT -53.205 -132.085 -52.875 -131.755 ;
        RECT -53.205 -133.445 -52.875 -133.115 ;
        RECT -53.205 -134.805 -52.875 -134.475 ;
        RECT -53.205 -136.165 -52.875 -135.835 ;
        RECT -53.205 -137.525 -52.875 -137.195 ;
        RECT -53.205 -138.885 -52.875 -138.555 ;
        RECT -53.205 -140.245 -52.875 -139.915 ;
        RECT -53.205 -141.605 -52.875 -141.275 ;
        RECT -53.205 -142.965 -52.875 -142.635 ;
        RECT -53.205 -144.325 -52.875 -143.995 ;
        RECT -53.205 -145.685 -52.875 -145.355 ;
        RECT -53.205 -147.045 -52.875 -146.715 ;
        RECT -53.205 -148.405 -52.875 -148.075 ;
        RECT -53.205 -149.765 -52.875 -149.435 ;
        RECT -53.205 -151.125 -52.875 -150.795 ;
        RECT -53.205 -152.485 -52.875 -152.155 ;
        RECT -53.205 -153.845 -52.875 -153.515 ;
        RECT -53.205 -155.205 -52.875 -154.875 ;
        RECT -53.205 -156.565 -52.875 -156.235 ;
        RECT -53.205 -157.925 -52.875 -157.595 ;
        RECT -53.205 -159.285 -52.875 -158.955 ;
        RECT -53.205 -160.645 -52.875 -160.315 ;
        RECT -53.205 -162.005 -52.875 -161.675 ;
        RECT -53.205 -163.365 -52.875 -163.035 ;
        RECT -53.205 -164.725 -52.875 -164.395 ;
        RECT -53.205 -166.085 -52.875 -165.755 ;
        RECT -53.205 -167.445 -52.875 -167.115 ;
        RECT -53.205 -170.165 -52.875 -169.835 ;
        RECT -53.205 -174.245 -52.875 -173.915 ;
        RECT -53.205 -175.725 -52.875 -175.395 ;
        RECT -53.205 -176.965 -52.875 -176.635 ;
        RECT -53.205 -178.325 -52.875 -177.995 ;
        RECT -53.205 -180.57 -52.875 -179.44 ;
        RECT -53.2 -180.685 -52.88 98.085 ;
    END
    PORT
      LAYER met3 ;
        RECT -51.845 241.32 -51.515 242.45 ;
        RECT -51.845 239.195 -51.515 239.525 ;
        RECT -51.845 237.835 -51.515 238.165 ;
        RECT -51.845 236.475 -51.515 236.805 ;
        RECT -51.845 235.115 -51.515 235.445 ;
        RECT -51.845 233.755 -51.515 234.085 ;
        RECT -51.845 232.395 -51.515 232.725 ;
        RECT -51.845 231.035 -51.515 231.365 ;
        RECT -51.845 229.675 -51.515 230.005 ;
        RECT -51.845 228.315 -51.515 228.645 ;
        RECT -51.845 226.955 -51.515 227.285 ;
        RECT -51.845 225.595 -51.515 225.925 ;
        RECT -51.845 224.235 -51.515 224.565 ;
        RECT -51.845 222.875 -51.515 223.205 ;
        RECT -51.845 221.515 -51.515 221.845 ;
        RECT -51.845 220.155 -51.515 220.485 ;
        RECT -51.845 218.795 -51.515 219.125 ;
        RECT -51.845 217.435 -51.515 217.765 ;
        RECT -51.845 216.075 -51.515 216.405 ;
        RECT -51.845 214.715 -51.515 215.045 ;
        RECT -51.845 213.355 -51.515 213.685 ;
        RECT -51.845 211.995 -51.515 212.325 ;
        RECT -51.845 210.635 -51.515 210.965 ;
        RECT -51.845 209.275 -51.515 209.605 ;
        RECT -51.845 207.915 -51.515 208.245 ;
        RECT -51.845 206.555 -51.515 206.885 ;
        RECT -51.845 205.195 -51.515 205.525 ;
        RECT -51.845 203.835 -51.515 204.165 ;
        RECT -51.845 202.475 -51.515 202.805 ;
        RECT -51.845 201.115 -51.515 201.445 ;
        RECT -51.845 199.755 -51.515 200.085 ;
        RECT -51.845 198.395 -51.515 198.725 ;
        RECT -51.845 197.035 -51.515 197.365 ;
        RECT -51.845 195.675 -51.515 196.005 ;
        RECT -51.845 194.315 -51.515 194.645 ;
        RECT -51.845 192.955 -51.515 193.285 ;
        RECT -51.845 191.595 -51.515 191.925 ;
        RECT -51.845 190.235 -51.515 190.565 ;
        RECT -51.845 188.875 -51.515 189.205 ;
        RECT -51.845 187.515 -51.515 187.845 ;
        RECT -51.845 186.155 -51.515 186.485 ;
        RECT -51.845 184.795 -51.515 185.125 ;
        RECT -51.845 183.435 -51.515 183.765 ;
        RECT -51.845 182.075 -51.515 182.405 ;
        RECT -51.845 180.715 -51.515 181.045 ;
        RECT -51.845 179.355 -51.515 179.685 ;
        RECT -51.845 177.995 -51.515 178.325 ;
        RECT -51.845 176.635 -51.515 176.965 ;
        RECT -51.845 175.275 -51.515 175.605 ;
        RECT -51.845 173.915 -51.515 174.245 ;
        RECT -51.845 172.555 -51.515 172.885 ;
        RECT -51.845 171.195 -51.515 171.525 ;
        RECT -51.845 169.835 -51.515 170.165 ;
        RECT -51.845 168.475 -51.515 168.805 ;
        RECT -51.845 167.115 -51.515 167.445 ;
        RECT -51.845 165.755 -51.515 166.085 ;
        RECT -51.845 164.395 -51.515 164.725 ;
        RECT -51.845 163.035 -51.515 163.365 ;
        RECT -51.845 161.675 -51.515 162.005 ;
        RECT -51.845 160.315 -51.515 160.645 ;
        RECT -51.845 158.955 -51.515 159.285 ;
        RECT -51.845 157.595 -51.515 157.925 ;
        RECT -51.845 156.235 -51.515 156.565 ;
        RECT -51.845 154.875 -51.515 155.205 ;
        RECT -51.845 153.515 -51.515 153.845 ;
        RECT -51.845 152.155 -51.515 152.485 ;
        RECT -51.845 150.795 -51.515 151.125 ;
        RECT -51.845 149.435 -51.515 149.765 ;
        RECT -51.845 148.075 -51.515 148.405 ;
        RECT -51.845 146.715 -51.515 147.045 ;
        RECT -51.845 145.355 -51.515 145.685 ;
        RECT -51.845 143.995 -51.515 144.325 ;
        RECT -51.845 142.635 -51.515 142.965 ;
        RECT -51.845 141.275 -51.515 141.605 ;
        RECT -51.845 139.915 -51.515 140.245 ;
        RECT -51.845 138.555 -51.515 138.885 ;
        RECT -51.845 137.225 -51.515 137.555 ;
        RECT -51.845 135.175 -51.515 135.505 ;
        RECT -51.845 132.815 -51.515 133.145 ;
        RECT -51.845 131.665 -51.515 131.995 ;
        RECT -51.845 129.655 -51.515 129.985 ;
        RECT -51.845 128.505 -51.515 128.835 ;
        RECT -51.845 126.495 -51.515 126.825 ;
        RECT -51.845 125.345 -51.515 125.675 ;
        RECT -51.845 123.335 -51.515 123.665 ;
        RECT -51.845 122.185 -51.515 122.515 ;
        RECT -51.845 120.175 -51.515 120.505 ;
        RECT -51.845 119.025 -51.515 119.355 ;
        RECT -51.845 117.185 -51.515 117.515 ;
        RECT -51.845 115.865 -51.515 116.195 ;
        RECT -51.845 113.855 -51.515 114.185 ;
        RECT -51.845 112.705 -51.515 113.035 ;
        RECT -51.845 110.695 -51.515 111.025 ;
        RECT -51.845 109.545 -51.515 109.875 ;
        RECT -51.845 107.535 -51.515 107.865 ;
        RECT -51.845 106.385 -51.515 106.715 ;
        RECT -51.845 104.375 -51.515 104.705 ;
        RECT -51.845 103.225 -51.515 103.555 ;
        RECT -51.845 100.865 -51.515 101.195 ;
        RECT -51.845 98.81 -51.515 99.14 ;
        RECT -51.845 97.755 -51.515 98.085 ;
        RECT -51.845 96.395 -51.515 96.725 ;
        RECT -51.845 95.035 -51.515 95.365 ;
        RECT -51.845 93.675 -51.515 94.005 ;
        RECT -51.845 92.315 -51.515 92.645 ;
        RECT -51.845 90.955 -51.515 91.285 ;
        RECT -51.845 89.595 -51.515 89.925 ;
        RECT -51.845 88.235 -51.515 88.565 ;
        RECT -51.845 86.875 -51.515 87.205 ;
        RECT -51.845 85.515 -51.515 85.845 ;
        RECT -51.845 84.155 -51.515 84.485 ;
        RECT -51.845 82.795 -51.515 83.125 ;
        RECT -51.845 81.435 -51.515 81.765 ;
        RECT -51.845 80.075 -51.515 80.405 ;
        RECT -51.845 78.715 -51.515 79.045 ;
        RECT -51.845 77.355 -51.515 77.685 ;
        RECT -51.845 75.995 -51.515 76.325 ;
        RECT -51.845 74.635 -51.515 74.965 ;
        RECT -51.845 73.275 -51.515 73.605 ;
        RECT -51.845 71.915 -51.515 72.245 ;
        RECT -51.845 70.555 -51.515 70.885 ;
        RECT -51.845 69.195 -51.515 69.525 ;
        RECT -51.845 67.835 -51.515 68.165 ;
        RECT -51.845 66.475 -51.515 66.805 ;
        RECT -51.845 65.115 -51.515 65.445 ;
        RECT -51.845 63.755 -51.515 64.085 ;
        RECT -51.845 62.395 -51.515 62.725 ;
        RECT -51.845 61.035 -51.515 61.365 ;
        RECT -51.845 59.675 -51.515 60.005 ;
        RECT -51.845 58.315 -51.515 58.645 ;
        RECT -51.845 56.955 -51.515 57.285 ;
        RECT -51.845 55.595 -51.515 55.925 ;
        RECT -51.845 54.235 -51.515 54.565 ;
        RECT -51.845 52.875 -51.515 53.205 ;
        RECT -51.845 51.515 -51.515 51.845 ;
        RECT -51.845 50.155 -51.515 50.485 ;
        RECT -51.845 48.795 -51.515 49.125 ;
        RECT -51.845 47.435 -51.515 47.765 ;
        RECT -51.845 46.075 -51.515 46.405 ;
        RECT -51.845 44.715 -51.515 45.045 ;
        RECT -51.845 43.355 -51.515 43.685 ;
        RECT -51.845 41.995 -51.515 42.325 ;
        RECT -51.845 40.635 -51.515 40.965 ;
        RECT -51.845 39.275 -51.515 39.605 ;
        RECT -51.845 37.915 -51.515 38.245 ;
        RECT -51.845 36.555 -51.515 36.885 ;
        RECT -51.845 35.195 -51.515 35.525 ;
        RECT -51.845 33.835 -51.515 34.165 ;
        RECT -51.845 32.475 -51.515 32.805 ;
        RECT -51.845 31.115 -51.515 31.445 ;
        RECT -51.845 29.755 -51.515 30.085 ;
        RECT -51.845 28.395 -51.515 28.725 ;
        RECT -51.845 27.035 -51.515 27.365 ;
        RECT -51.845 25.675 -51.515 26.005 ;
        RECT -51.845 24.315 -51.515 24.645 ;
        RECT -51.845 22.955 -51.515 23.285 ;
        RECT -51.845 21.595 -51.515 21.925 ;
        RECT -51.845 20.235 -51.515 20.565 ;
        RECT -51.845 18.875 -51.515 19.205 ;
        RECT -51.845 17.515 -51.515 17.845 ;
        RECT -51.845 16.155 -51.515 16.485 ;
        RECT -51.845 14.795 -51.515 15.125 ;
        RECT -51.845 13.435 -51.515 13.765 ;
        RECT -51.845 12.075 -51.515 12.405 ;
        RECT -51.845 10.715 -51.515 11.045 ;
        RECT -51.845 9.355 -51.515 9.685 ;
        RECT -51.845 7.995 -51.515 8.325 ;
        RECT -51.845 6.635 -51.515 6.965 ;
        RECT -51.845 5.275 -51.515 5.605 ;
        RECT -51.845 3.915 -51.515 4.245 ;
        RECT -51.845 2.555 -51.515 2.885 ;
        RECT -51.845 1.195 -51.515 1.525 ;
        RECT -51.845 -0.165 -51.515 0.165 ;
        RECT -51.845 -2.885 -51.515 -2.555 ;
        RECT -51.845 -4.245 -51.515 -3.915 ;
        RECT -51.845 -5.605 -51.515 -5.275 ;
        RECT -51.845 -6.965 -51.515 -6.635 ;
        RECT -51.845 -8.325 -51.515 -7.995 ;
        RECT -51.845 -9.685 -51.515 -9.355 ;
        RECT -51.845 -11.045 -51.515 -10.715 ;
        RECT -51.845 -12.405 -51.515 -12.075 ;
        RECT -51.845 -13.765 -51.515 -13.435 ;
        RECT -51.845 -15.125 -51.515 -14.795 ;
        RECT -51.845 -16.485 -51.515 -16.155 ;
        RECT -51.845 -17.845 -51.515 -17.515 ;
        RECT -51.845 -19.205 -51.515 -18.875 ;
        RECT -51.845 -20.565 -51.515 -20.235 ;
        RECT -51.845 -21.925 -51.515 -21.595 ;
        RECT -51.845 -23.285 -51.515 -22.955 ;
        RECT -51.845 -24.645 -51.515 -24.315 ;
        RECT -51.845 -28.725 -51.515 -28.395 ;
        RECT -51.845 -30.085 -51.515 -29.755 ;
        RECT -51.845 -31.445 -51.515 -31.115 ;
        RECT -51.845 -32.805 -51.515 -32.475 ;
        RECT -51.845 -34.165 -51.515 -33.835 ;
        RECT -51.845 -35.525 -51.515 -35.195 ;
        RECT -51.845 -36.885 -51.515 -36.555 ;
        RECT -51.845 -38.245 -51.515 -37.915 ;
        RECT -51.845 -39.605 -51.515 -39.275 ;
        RECT -51.845 -40.965 -51.515 -40.635 ;
        RECT -51.845 -42.325 -51.515 -41.995 ;
        RECT -51.845 -43.685 -51.515 -43.355 ;
        RECT -51.845 -45.045 -51.515 -44.715 ;
        RECT -51.845 -46.405 -51.515 -46.075 ;
        RECT -51.845 -47.765 -51.515 -47.435 ;
        RECT -51.845 -49.125 -51.515 -48.795 ;
        RECT -51.845 -50.485 -51.515 -50.155 ;
        RECT -51.845 -51.845 -51.515 -51.515 ;
        RECT -51.845 -53.205 -51.515 -52.875 ;
        RECT -51.845 -54.565 -51.515 -54.235 ;
        RECT -51.845 -55.925 -51.515 -55.595 ;
        RECT -51.845 -57.285 -51.515 -56.955 ;
        RECT -51.845 -58.645 -51.515 -58.315 ;
        RECT -51.845 -60.005 -51.515 -59.675 ;
        RECT -51.845 -61.365 -51.515 -61.035 ;
        RECT -51.845 -62.725 -51.515 -62.395 ;
        RECT -51.845 -64.085 -51.515 -63.755 ;
        RECT -51.845 -65.445 -51.515 -65.115 ;
        RECT -51.845 -66.805 -51.515 -66.475 ;
        RECT -51.845 -68.165 -51.515 -67.835 ;
        RECT -51.845 -69.525 -51.515 -69.195 ;
        RECT -51.845 -70.885 -51.515 -70.555 ;
        RECT -51.845 -72.245 -51.515 -71.915 ;
        RECT -51.845 -73.605 -51.515 -73.275 ;
        RECT -51.845 -74.965 -51.515 -74.635 ;
        RECT -51.845 -76.325 -51.515 -75.995 ;
        RECT -51.845 -77.685 -51.515 -77.355 ;
        RECT -51.845 -79.045 -51.515 -78.715 ;
        RECT -51.845 -80.405 -51.515 -80.075 ;
        RECT -51.845 -81.765 -51.515 -81.435 ;
        RECT -51.845 -83.125 -51.515 -82.795 ;
        RECT -51.845 -84.485 -51.515 -84.155 ;
        RECT -51.845 -85.845 -51.515 -85.515 ;
        RECT -51.845 -87.205 -51.515 -86.875 ;
        RECT -51.845 -88.565 -51.515 -88.235 ;
        RECT -51.845 -89.925 -51.515 -89.595 ;
        RECT -51.845 -92.645 -51.515 -92.315 ;
        RECT -51.845 -94.005 -51.515 -93.675 ;
        RECT -51.845 -95.365 -51.515 -95.035 ;
        RECT -51.845 -96.725 -51.515 -96.395 ;
        RECT -51.845 -98.73 -51.515 -98.4 ;
        RECT -51.845 -99.445 -51.515 -99.115 ;
        RECT -51.845 -102.165 -51.515 -101.835 ;
        RECT -51.845 -103.525 -51.515 -103.195 ;
        RECT -51.845 -104.885 -51.515 -104.555 ;
        RECT -51.845 -106.87 -51.515 -106.54 ;
        RECT -51.845 -107.605 -51.515 -107.275 ;
        RECT -51.845 -108.965 -51.515 -108.635 ;
        RECT -51.845 -114.405 -51.515 -114.075 ;
        RECT -51.845 -115.765 -51.515 -115.435 ;
        RECT -51.845 -117.125 -51.515 -116.795 ;
        RECT -51.845 -118.485 -51.515 -118.155 ;
        RECT -51.845 -122.565 -51.515 -122.235 ;
        RECT -51.845 -123.925 -51.515 -123.595 ;
        RECT -51.845 -125.285 -51.515 -124.955 ;
        RECT -51.845 -126.645 -51.515 -126.315 ;
        RECT -51.845 -128.005 -51.515 -127.675 ;
        RECT -51.845 -129.365 -51.515 -129.035 ;
        RECT -51.845 -130.725 -51.515 -130.395 ;
        RECT -51.845 -132.085 -51.515 -131.755 ;
        RECT -51.845 -133.445 -51.515 -133.115 ;
        RECT -51.845 -134.805 -51.515 -134.475 ;
        RECT -51.845 -136.165 -51.515 -135.835 ;
        RECT -51.845 -137.525 -51.515 -137.195 ;
        RECT -51.845 -138.885 -51.515 -138.555 ;
        RECT -51.845 -140.245 -51.515 -139.915 ;
        RECT -51.845 -141.605 -51.515 -141.275 ;
        RECT -51.845 -142.965 -51.515 -142.635 ;
        RECT -51.845 -144.325 -51.515 -143.995 ;
        RECT -51.845 -145.685 -51.515 -145.355 ;
        RECT -51.845 -147.045 -51.515 -146.715 ;
        RECT -51.845 -148.405 -51.515 -148.075 ;
        RECT -51.845 -149.765 -51.515 -149.435 ;
        RECT -51.845 -151.125 -51.515 -150.795 ;
        RECT -51.845 -152.485 -51.515 -152.155 ;
        RECT -51.845 -153.845 -51.515 -153.515 ;
        RECT -51.845 -155.205 -51.515 -154.875 ;
        RECT -51.845 -156.565 -51.515 -156.235 ;
        RECT -51.845 -157.925 -51.515 -157.595 ;
        RECT -51.845 -159.285 -51.515 -158.955 ;
        RECT -51.845 -160.645 -51.515 -160.315 ;
        RECT -51.845 -162.005 -51.515 -161.675 ;
        RECT -51.845 -163.365 -51.515 -163.035 ;
        RECT -51.845 -164.725 -51.515 -164.395 ;
        RECT -51.845 -166.085 -51.515 -165.755 ;
        RECT -51.845 -167.445 -51.515 -167.115 ;
        RECT -51.845 -170.165 -51.515 -169.835 ;
        RECT -51.845 -172.885 -51.515 -172.555 ;
        RECT -51.845 -174.245 -51.515 -173.915 ;
        RECT -51.845 -175.725 -51.515 -175.395 ;
        RECT -51.845 -176.965 -51.515 -176.635 ;
        RECT -51.845 -178.325 -51.515 -177.995 ;
        RECT -51.845 -180.57 -51.515 -179.44 ;
        RECT -51.84 -180.685 -51.52 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -50.485 184.795 -50.155 185.125 ;
        RECT -50.485 183.435 -50.155 183.765 ;
        RECT -50.485 182.075 -50.155 182.405 ;
        RECT -50.485 180.715 -50.155 181.045 ;
        RECT -50.485 179.355 -50.155 179.685 ;
        RECT -50.485 177.995 -50.155 178.325 ;
        RECT -50.485 176.635 -50.155 176.965 ;
        RECT -50.485 175.275 -50.155 175.605 ;
        RECT -50.485 173.915 -50.155 174.245 ;
        RECT -50.485 172.555 -50.155 172.885 ;
        RECT -50.485 171.195 -50.155 171.525 ;
        RECT -50.485 169.835 -50.155 170.165 ;
        RECT -50.485 168.475 -50.155 168.805 ;
        RECT -50.485 167.115 -50.155 167.445 ;
        RECT -50.485 165.755 -50.155 166.085 ;
        RECT -50.485 164.395 -50.155 164.725 ;
        RECT -50.485 163.035 -50.155 163.365 ;
        RECT -50.485 161.675 -50.155 162.005 ;
        RECT -50.485 160.315 -50.155 160.645 ;
        RECT -50.485 158.955 -50.155 159.285 ;
        RECT -50.485 157.595 -50.155 157.925 ;
        RECT -50.485 156.235 -50.155 156.565 ;
        RECT -50.485 154.875 -50.155 155.205 ;
        RECT -50.485 153.515 -50.155 153.845 ;
        RECT -50.485 152.155 -50.155 152.485 ;
        RECT -50.485 150.795 -50.155 151.125 ;
        RECT -50.485 149.435 -50.155 149.765 ;
        RECT -50.485 148.075 -50.155 148.405 ;
        RECT -50.485 146.715 -50.155 147.045 ;
        RECT -50.485 145.355 -50.155 145.685 ;
        RECT -50.485 143.995 -50.155 144.325 ;
        RECT -50.485 142.635 -50.155 142.965 ;
        RECT -50.485 141.275 -50.155 141.605 ;
        RECT -50.485 139.915 -50.155 140.245 ;
        RECT -50.485 138.555 -50.155 138.885 ;
        RECT -50.485 137.225 -50.155 137.555 ;
        RECT -50.485 135.175 -50.155 135.505 ;
        RECT -50.485 132.815 -50.155 133.145 ;
        RECT -50.485 131.665 -50.155 131.995 ;
        RECT -50.485 129.655 -50.155 129.985 ;
        RECT -50.485 128.505 -50.155 128.835 ;
        RECT -50.485 126.495 -50.155 126.825 ;
        RECT -50.485 125.345 -50.155 125.675 ;
        RECT -50.485 123.335 -50.155 123.665 ;
        RECT -50.485 122.185 -50.155 122.515 ;
        RECT -50.485 120.175 -50.155 120.505 ;
        RECT -50.485 119.025 -50.155 119.355 ;
        RECT -50.485 117.185 -50.155 117.515 ;
        RECT -50.485 115.865 -50.155 116.195 ;
        RECT -50.485 113.855 -50.155 114.185 ;
        RECT -50.485 112.705 -50.155 113.035 ;
        RECT -50.485 110.695 -50.155 111.025 ;
        RECT -50.485 109.545 -50.155 109.875 ;
        RECT -50.485 107.535 -50.155 107.865 ;
        RECT -50.485 106.385 -50.155 106.715 ;
        RECT -50.485 104.375 -50.155 104.705 ;
        RECT -50.485 103.225 -50.155 103.555 ;
        RECT -50.485 100.865 -50.155 101.195 ;
        RECT -50.485 98.81 -50.155 99.14 ;
        RECT -50.485 97.755 -50.155 98.085 ;
        RECT -50.485 96.395 -50.155 96.725 ;
        RECT -50.485 95.035 -50.155 95.365 ;
        RECT -50.485 93.675 -50.155 94.005 ;
        RECT -50.485 92.315 -50.155 92.645 ;
        RECT -50.485 90.955 -50.155 91.285 ;
        RECT -50.485 89.595 -50.155 89.925 ;
        RECT -50.485 88.235 -50.155 88.565 ;
        RECT -50.485 86.875 -50.155 87.205 ;
        RECT -50.485 85.515 -50.155 85.845 ;
        RECT -50.485 84.155 -50.155 84.485 ;
        RECT -50.485 82.795 -50.155 83.125 ;
        RECT -50.485 81.435 -50.155 81.765 ;
        RECT -50.485 80.075 -50.155 80.405 ;
        RECT -50.485 78.715 -50.155 79.045 ;
        RECT -50.485 77.355 -50.155 77.685 ;
        RECT -50.485 75.995 -50.155 76.325 ;
        RECT -50.485 74.635 -50.155 74.965 ;
        RECT -50.485 73.275 -50.155 73.605 ;
        RECT -50.485 71.915 -50.155 72.245 ;
        RECT -50.485 70.555 -50.155 70.885 ;
        RECT -50.485 69.195 -50.155 69.525 ;
        RECT -50.485 67.835 -50.155 68.165 ;
        RECT -50.485 66.475 -50.155 66.805 ;
        RECT -50.485 65.115 -50.155 65.445 ;
        RECT -50.485 63.755 -50.155 64.085 ;
        RECT -50.485 62.395 -50.155 62.725 ;
        RECT -50.485 61.035 -50.155 61.365 ;
        RECT -50.485 59.675 -50.155 60.005 ;
        RECT -50.485 58.315 -50.155 58.645 ;
        RECT -50.485 56.955 -50.155 57.285 ;
        RECT -50.485 55.595 -50.155 55.925 ;
        RECT -50.485 54.235 -50.155 54.565 ;
        RECT -50.485 52.875 -50.155 53.205 ;
        RECT -50.485 51.515 -50.155 51.845 ;
        RECT -50.485 50.155 -50.155 50.485 ;
        RECT -50.485 48.795 -50.155 49.125 ;
        RECT -50.485 47.435 -50.155 47.765 ;
        RECT -50.485 46.075 -50.155 46.405 ;
        RECT -50.485 44.715 -50.155 45.045 ;
        RECT -50.485 43.355 -50.155 43.685 ;
        RECT -50.485 41.995 -50.155 42.325 ;
        RECT -50.485 40.635 -50.155 40.965 ;
        RECT -50.485 39.275 -50.155 39.605 ;
        RECT -50.485 37.915 -50.155 38.245 ;
        RECT -50.485 36.555 -50.155 36.885 ;
        RECT -50.485 35.195 -50.155 35.525 ;
        RECT -50.485 33.835 -50.155 34.165 ;
        RECT -50.485 32.475 -50.155 32.805 ;
        RECT -50.485 31.115 -50.155 31.445 ;
        RECT -50.485 29.755 -50.155 30.085 ;
        RECT -50.485 28.395 -50.155 28.725 ;
        RECT -50.485 27.035 -50.155 27.365 ;
        RECT -50.485 25.675 -50.155 26.005 ;
        RECT -50.485 24.315 -50.155 24.645 ;
        RECT -50.485 22.955 -50.155 23.285 ;
        RECT -50.485 21.595 -50.155 21.925 ;
        RECT -50.485 20.235 -50.155 20.565 ;
        RECT -50.485 18.875 -50.155 19.205 ;
        RECT -50.485 17.515 -50.155 17.845 ;
        RECT -50.485 16.155 -50.155 16.485 ;
        RECT -50.485 14.795 -50.155 15.125 ;
        RECT -50.485 13.435 -50.155 13.765 ;
        RECT -50.485 12.075 -50.155 12.405 ;
        RECT -50.485 10.715 -50.155 11.045 ;
        RECT -50.485 9.355 -50.155 9.685 ;
        RECT -50.485 7.995 -50.155 8.325 ;
        RECT -50.485 6.635 -50.155 6.965 ;
        RECT -50.485 5.275 -50.155 5.605 ;
        RECT -50.485 3.915 -50.155 4.245 ;
        RECT -50.485 2.555 -50.155 2.885 ;
        RECT -50.485 1.195 -50.155 1.525 ;
        RECT -50.485 -0.165 -50.155 0.165 ;
        RECT -50.485 -2.885 -50.155 -2.555 ;
        RECT -50.485 -4.245 -50.155 -3.915 ;
        RECT -50.485 -5.605 -50.155 -5.275 ;
        RECT -50.485 -6.965 -50.155 -6.635 ;
        RECT -50.485 -8.325 -50.155 -7.995 ;
        RECT -50.485 -9.685 -50.155 -9.355 ;
        RECT -50.485 -11.045 -50.155 -10.715 ;
        RECT -50.485 -12.405 -50.155 -12.075 ;
        RECT -50.485 -15.125 -50.155 -14.795 ;
        RECT -50.485 -16.485 -50.155 -16.155 ;
        RECT -50.485 -17.845 -50.155 -17.515 ;
        RECT -50.485 -19.205 -50.155 -18.875 ;
        RECT -50.485 -20.565 -50.155 -20.235 ;
        RECT -50.485 -21.925 -50.155 -21.595 ;
        RECT -50.485 -23.285 -50.155 -22.955 ;
        RECT -50.485 -24.645 -50.155 -24.315 ;
        RECT -50.485 -28.725 -50.155 -28.395 ;
        RECT -50.485 -30.085 -50.155 -29.755 ;
        RECT -50.485 -31.445 -50.155 -31.115 ;
        RECT -50.485 -32.805 -50.155 -32.475 ;
        RECT -50.485 -34.165 -50.155 -33.835 ;
        RECT -50.485 -35.525 -50.155 -35.195 ;
        RECT -50.485 -36.885 -50.155 -36.555 ;
        RECT -50.485 -38.245 -50.155 -37.915 ;
        RECT -50.485 -39.605 -50.155 -39.275 ;
        RECT -50.485 -40.965 -50.155 -40.635 ;
        RECT -50.485 -42.325 -50.155 -41.995 ;
        RECT -50.485 -43.685 -50.155 -43.355 ;
        RECT -50.485 -45.045 -50.155 -44.715 ;
        RECT -50.485 -46.405 -50.155 -46.075 ;
        RECT -50.485 -47.765 -50.155 -47.435 ;
        RECT -50.485 -49.125 -50.155 -48.795 ;
        RECT -50.485 -50.485 -50.155 -50.155 ;
        RECT -50.485 -51.845 -50.155 -51.515 ;
        RECT -50.485 -53.205 -50.155 -52.875 ;
        RECT -50.485 -54.565 -50.155 -54.235 ;
        RECT -50.485 -55.925 -50.155 -55.595 ;
        RECT -50.485 -57.285 -50.155 -56.955 ;
        RECT -50.485 -58.645 -50.155 -58.315 ;
        RECT -50.485 -60.005 -50.155 -59.675 ;
        RECT -50.485 -61.365 -50.155 -61.035 ;
        RECT -50.485 -62.725 -50.155 -62.395 ;
        RECT -50.485 -64.085 -50.155 -63.755 ;
        RECT -50.485 -65.445 -50.155 -65.115 ;
        RECT -50.485 -66.805 -50.155 -66.475 ;
        RECT -50.485 -68.165 -50.155 -67.835 ;
        RECT -50.485 -69.525 -50.155 -69.195 ;
        RECT -50.485 -70.885 -50.155 -70.555 ;
        RECT -50.485 -72.245 -50.155 -71.915 ;
        RECT -50.485 -73.605 -50.155 -73.275 ;
        RECT -50.485 -74.965 -50.155 -74.635 ;
        RECT -50.485 -76.325 -50.155 -75.995 ;
        RECT -50.485 -77.685 -50.155 -77.355 ;
        RECT -50.485 -79.045 -50.155 -78.715 ;
        RECT -50.485 -80.405 -50.155 -80.075 ;
        RECT -50.485 -81.765 -50.155 -81.435 ;
        RECT -50.485 -83.125 -50.155 -82.795 ;
        RECT -50.485 -84.485 -50.155 -84.155 ;
        RECT -50.485 -85.845 -50.155 -85.515 ;
        RECT -50.485 -87.205 -50.155 -86.875 ;
        RECT -50.485 -88.565 -50.155 -88.235 ;
        RECT -50.485 -89.925 -50.155 -89.595 ;
        RECT -50.485 -92.645 -50.155 -92.315 ;
        RECT -50.485 -94.005 -50.155 -93.675 ;
        RECT -50.485 -95.365 -50.155 -95.035 ;
        RECT -50.485 -96.725 -50.155 -96.395 ;
        RECT -50.485 -98.73 -50.155 -98.4 ;
        RECT -50.485 -99.445 -50.155 -99.115 ;
        RECT -50.485 -102.165 -50.155 -101.835 ;
        RECT -50.485 -103.525 -50.155 -103.195 ;
        RECT -50.485 -104.885 -50.155 -104.555 ;
        RECT -50.485 -106.87 -50.155 -106.54 ;
        RECT -50.485 -107.605 -50.155 -107.275 ;
        RECT -50.485 -108.965 -50.155 -108.635 ;
        RECT -50.485 -114.405 -50.155 -114.075 ;
        RECT -50.485 -115.765 -50.155 -115.435 ;
        RECT -50.485 -117.125 -50.155 -116.795 ;
        RECT -50.485 -118.485 -50.155 -118.155 ;
        RECT -50.485 -122.565 -50.155 -122.235 ;
        RECT -50.485 -123.925 -50.155 -123.595 ;
        RECT -50.485 -125.285 -50.155 -124.955 ;
        RECT -50.485 -126.645 -50.155 -126.315 ;
        RECT -50.485 -128.005 -50.155 -127.675 ;
        RECT -50.485 -129.365 -50.155 -129.035 ;
        RECT -50.485 -130.725 -50.155 -130.395 ;
        RECT -50.485 -132.085 -50.155 -131.755 ;
        RECT -50.485 -133.445 -50.155 -133.115 ;
        RECT -50.485 -134.805 -50.155 -134.475 ;
        RECT -50.485 -136.165 -50.155 -135.835 ;
        RECT -50.485 -137.525 -50.155 -137.195 ;
        RECT -50.485 -138.885 -50.155 -138.555 ;
        RECT -50.485 -140.245 -50.155 -139.915 ;
        RECT -50.485 -141.605 -50.155 -141.275 ;
        RECT -50.485 -142.965 -50.155 -142.635 ;
        RECT -50.485 -144.325 -50.155 -143.995 ;
        RECT -50.485 -145.685 -50.155 -145.355 ;
        RECT -50.485 -147.045 -50.155 -146.715 ;
        RECT -50.485 -148.405 -50.155 -148.075 ;
        RECT -50.485 -149.765 -50.155 -149.435 ;
        RECT -50.485 -151.125 -50.155 -150.795 ;
        RECT -50.485 -152.485 -50.155 -152.155 ;
        RECT -50.485 -153.845 -50.155 -153.515 ;
        RECT -50.485 -155.205 -50.155 -154.875 ;
        RECT -50.485 -156.565 -50.155 -156.235 ;
        RECT -50.485 -157.925 -50.155 -157.595 ;
        RECT -50.485 -159.285 -50.155 -158.955 ;
        RECT -50.485 -160.645 -50.155 -160.315 ;
        RECT -50.485 -162.005 -50.155 -161.675 ;
        RECT -50.485 -163.365 -50.155 -163.035 ;
        RECT -50.485 -164.725 -50.155 -164.395 ;
        RECT -50.485 -166.085 -50.155 -165.755 ;
        RECT -50.485 -167.445 -50.155 -167.115 ;
        RECT -50.485 -170.165 -50.155 -169.835 ;
        RECT -50.485 -172.885 -50.155 -172.555 ;
        RECT -50.485 -174.245 -50.155 -173.915 ;
        RECT -50.485 -175.725 -50.155 -175.395 ;
        RECT -50.485 -176.965 -50.155 -176.635 ;
        RECT -50.485 -178.325 -50.155 -177.995 ;
        RECT -50.485 -180.57 -50.155 -179.44 ;
        RECT -50.48 -180.685 -50.16 242.565 ;
        RECT -50.485 241.32 -50.155 242.45 ;
        RECT -50.485 239.195 -50.155 239.525 ;
        RECT -50.485 237.835 -50.155 238.165 ;
        RECT -50.485 236.475 -50.155 236.805 ;
        RECT -50.485 235.115 -50.155 235.445 ;
        RECT -50.485 233.755 -50.155 234.085 ;
        RECT -50.485 232.395 -50.155 232.725 ;
        RECT -50.485 231.035 -50.155 231.365 ;
        RECT -50.485 229.675 -50.155 230.005 ;
        RECT -50.485 228.315 -50.155 228.645 ;
        RECT -50.485 226.955 -50.155 227.285 ;
        RECT -50.485 225.595 -50.155 225.925 ;
        RECT -50.485 224.235 -50.155 224.565 ;
        RECT -50.485 222.875 -50.155 223.205 ;
        RECT -50.485 221.515 -50.155 221.845 ;
        RECT -50.485 220.155 -50.155 220.485 ;
        RECT -50.485 218.795 -50.155 219.125 ;
        RECT -50.485 217.435 -50.155 217.765 ;
        RECT -50.485 216.075 -50.155 216.405 ;
        RECT -50.485 214.715 -50.155 215.045 ;
        RECT -50.485 213.355 -50.155 213.685 ;
        RECT -50.485 211.995 -50.155 212.325 ;
        RECT -50.485 210.635 -50.155 210.965 ;
        RECT -50.485 209.275 -50.155 209.605 ;
        RECT -50.485 207.915 -50.155 208.245 ;
        RECT -50.485 206.555 -50.155 206.885 ;
        RECT -50.485 205.195 -50.155 205.525 ;
        RECT -50.485 203.835 -50.155 204.165 ;
        RECT -50.485 202.475 -50.155 202.805 ;
        RECT -50.485 201.115 -50.155 201.445 ;
        RECT -50.485 199.755 -50.155 200.085 ;
        RECT -50.485 198.395 -50.155 198.725 ;
        RECT -50.485 197.035 -50.155 197.365 ;
        RECT -50.485 195.675 -50.155 196.005 ;
        RECT -50.485 194.315 -50.155 194.645 ;
        RECT -50.485 192.955 -50.155 193.285 ;
        RECT -50.485 191.595 -50.155 191.925 ;
        RECT -50.485 190.235 -50.155 190.565 ;
        RECT -50.485 188.875 -50.155 189.205 ;
        RECT -50.485 187.515 -50.155 187.845 ;
        RECT -50.485 186.155 -50.155 186.485 ;
    END
    PORT
      LAYER met3 ;
        RECT -61.365 -174.245 -61.035 -173.915 ;
        RECT -61.365 -175.725 -61.035 -175.395 ;
        RECT -61.365 -176.965 -61.035 -176.635 ;
        RECT -61.365 -178.325 -61.035 -177.995 ;
        RECT -61.365 -180.57 -61.035 -179.44 ;
        RECT -61.36 -180.685 -61.04 -173.915 ;
    END
    PORT
      LAYER met3 ;
        RECT -60.005 241.32 -59.675 242.45 ;
        RECT -60.005 239.195 -59.675 239.525 ;
        RECT -60.005 237.835 -59.675 238.165 ;
        RECT -60.005 236.475 -59.675 236.805 ;
        RECT -60.005 235.115 -59.675 235.445 ;
        RECT -60.005 233.755 -59.675 234.085 ;
        RECT -60.005 232.395 -59.675 232.725 ;
        RECT -60.005 231.035 -59.675 231.365 ;
        RECT -60.005 229.675 -59.675 230.005 ;
        RECT -60.005 228.315 -59.675 228.645 ;
        RECT -60.005 226.955 -59.675 227.285 ;
        RECT -60.005 225.595 -59.675 225.925 ;
        RECT -60.005 224.235 -59.675 224.565 ;
        RECT -60.005 222.875 -59.675 223.205 ;
        RECT -60.005 221.515 -59.675 221.845 ;
        RECT -60.005 220.155 -59.675 220.485 ;
        RECT -60.005 218.795 -59.675 219.125 ;
        RECT -60.005 217.435 -59.675 217.765 ;
        RECT -60.005 216.075 -59.675 216.405 ;
        RECT -60.005 214.715 -59.675 215.045 ;
        RECT -60.005 213.355 -59.675 213.685 ;
        RECT -60.005 211.995 -59.675 212.325 ;
        RECT -60.005 210.635 -59.675 210.965 ;
        RECT -60.005 209.275 -59.675 209.605 ;
        RECT -60.005 207.915 -59.675 208.245 ;
        RECT -60.005 206.555 -59.675 206.885 ;
        RECT -60.005 205.195 -59.675 205.525 ;
        RECT -60.005 203.835 -59.675 204.165 ;
        RECT -60.005 202.475 -59.675 202.805 ;
        RECT -60.005 201.115 -59.675 201.445 ;
        RECT -60.005 199.755 -59.675 200.085 ;
        RECT -60.005 198.395 -59.675 198.725 ;
        RECT -60.005 197.035 -59.675 197.365 ;
        RECT -60.005 195.675 -59.675 196.005 ;
        RECT -60.005 194.315 -59.675 194.645 ;
        RECT -60.005 192.955 -59.675 193.285 ;
        RECT -60.005 191.595 -59.675 191.925 ;
        RECT -60.005 190.235 -59.675 190.565 ;
        RECT -60.005 188.875 -59.675 189.205 ;
        RECT -60.005 187.515 -59.675 187.845 ;
        RECT -60.005 186.155 -59.675 186.485 ;
        RECT -60.005 184.795 -59.675 185.125 ;
        RECT -60.005 183.435 -59.675 183.765 ;
        RECT -60.005 182.075 -59.675 182.405 ;
        RECT -60.005 180.715 -59.675 181.045 ;
        RECT -60.005 179.355 -59.675 179.685 ;
        RECT -60.005 177.995 -59.675 178.325 ;
        RECT -60.005 176.635 -59.675 176.965 ;
        RECT -60.005 175.275 -59.675 175.605 ;
        RECT -60.005 173.915 -59.675 174.245 ;
        RECT -60.005 172.555 -59.675 172.885 ;
        RECT -60.005 171.195 -59.675 171.525 ;
        RECT -60.005 169.835 -59.675 170.165 ;
        RECT -60.005 168.475 -59.675 168.805 ;
        RECT -60.005 167.115 -59.675 167.445 ;
        RECT -60.005 165.755 -59.675 166.085 ;
        RECT -60.005 164.395 -59.675 164.725 ;
        RECT -60.005 163.035 -59.675 163.365 ;
        RECT -60.005 161.675 -59.675 162.005 ;
        RECT -60.005 160.315 -59.675 160.645 ;
        RECT -60.005 158.955 -59.675 159.285 ;
        RECT -60.005 157.595 -59.675 157.925 ;
        RECT -60.005 156.235 -59.675 156.565 ;
        RECT -60.005 154.875 -59.675 155.205 ;
        RECT -60.005 153.515 -59.675 153.845 ;
        RECT -60.005 152.155 -59.675 152.485 ;
        RECT -60.005 150.795 -59.675 151.125 ;
        RECT -60.005 149.435 -59.675 149.765 ;
        RECT -60.005 148.075 -59.675 148.405 ;
        RECT -60.005 146.715 -59.675 147.045 ;
        RECT -60.005 145.355 -59.675 145.685 ;
        RECT -60.005 143.995 -59.675 144.325 ;
        RECT -60.005 142.635 -59.675 142.965 ;
        RECT -60.005 141.275 -59.675 141.605 ;
        RECT -60.005 139.915 -59.675 140.245 ;
        RECT -60.005 138.555 -59.675 138.885 ;
        RECT -60.005 137.225 -59.675 137.555 ;
        RECT -60.005 135.175 -59.675 135.505 ;
        RECT -60.005 132.815 -59.675 133.145 ;
        RECT -60.005 131.665 -59.675 131.995 ;
        RECT -60.005 129.655 -59.675 129.985 ;
        RECT -60.005 128.505 -59.675 128.835 ;
        RECT -60.005 126.495 -59.675 126.825 ;
        RECT -60.005 125.345 -59.675 125.675 ;
        RECT -60.005 123.335 -59.675 123.665 ;
        RECT -60.005 122.185 -59.675 122.515 ;
        RECT -60.005 120.175 -59.675 120.505 ;
        RECT -60.005 119.025 -59.675 119.355 ;
        RECT -60.005 117.185 -59.675 117.515 ;
        RECT -60.005 115.865 -59.675 116.195 ;
        RECT -60.005 113.855 -59.675 114.185 ;
        RECT -60.005 112.705 -59.675 113.035 ;
        RECT -60.005 110.695 -59.675 111.025 ;
        RECT -60.005 109.545 -59.675 109.875 ;
        RECT -60.005 107.535 -59.675 107.865 ;
        RECT -60.005 106.385 -59.675 106.715 ;
        RECT -60.005 104.375 -59.675 104.705 ;
        RECT -60.005 103.225 -59.675 103.555 ;
        RECT -60.005 100.865 -59.675 101.195 ;
        RECT -60.005 98.81 -59.675 99.14 ;
        RECT -60.005 97.755 -59.675 98.085 ;
        RECT -60.005 96.395 -59.675 96.725 ;
        RECT -60.005 95.035 -59.675 95.365 ;
        RECT -60.005 93.675 -59.675 94.005 ;
        RECT -60.005 92.315 -59.675 92.645 ;
        RECT -60.005 90.955 -59.675 91.285 ;
        RECT -60.005 89.595 -59.675 89.925 ;
        RECT -60.005 88.235 -59.675 88.565 ;
        RECT -60 86.88 -59.68 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -60.005 -122.565 -59.675 -122.235 ;
        RECT -60.005 -123.925 -59.675 -123.595 ;
        RECT -60.005 -125.285 -59.675 -124.955 ;
        RECT -60.005 -126.645 -59.675 -126.315 ;
        RECT -60.005 -128.005 -59.675 -127.675 ;
        RECT -60.005 -129.365 -59.675 -129.035 ;
        RECT -60.005 -130.725 -59.675 -130.395 ;
        RECT -60.005 -132.085 -59.675 -131.755 ;
        RECT -60.005 -133.445 -59.675 -133.115 ;
        RECT -60.005 -134.805 -59.675 -134.475 ;
        RECT -60.005 -136.165 -59.675 -135.835 ;
        RECT -60.005 -137.525 -59.675 -137.195 ;
        RECT -60.005 -138.885 -59.675 -138.555 ;
        RECT -60.005 -140.245 -59.675 -139.915 ;
        RECT -60.005 -141.605 -59.675 -141.275 ;
        RECT -60.005 -142.965 -59.675 -142.635 ;
        RECT -60.005 -144.325 -59.675 -143.995 ;
        RECT -60.005 -145.685 -59.675 -145.355 ;
        RECT -60.005 -147.045 -59.675 -146.715 ;
        RECT -60.005 -148.405 -59.675 -148.075 ;
        RECT -60.005 -149.765 -59.675 -149.435 ;
        RECT -60.005 -151.125 -59.675 -150.795 ;
        RECT -60.005 -152.485 -59.675 -152.155 ;
        RECT -60.005 -153.845 -59.675 -153.515 ;
        RECT -60.005 -155.205 -59.675 -154.875 ;
        RECT -60.005 -156.565 -59.675 -156.235 ;
        RECT -60.005 -157.925 -59.675 -157.595 ;
        RECT -60.005 -159.285 -59.675 -158.955 ;
        RECT -60.005 -160.645 -59.675 -160.315 ;
        RECT -60.005 -162.005 -59.675 -161.675 ;
        RECT -60.005 -163.365 -59.675 -163.035 ;
        RECT -60.005 -164.725 -59.675 -164.395 ;
        RECT -60.005 -166.085 -59.675 -165.755 ;
        RECT -60.005 -167.445 -59.675 -167.115 ;
        RECT -60.005 -170.165 -59.675 -169.835 ;
        RECT -60.005 -174.245 -59.675 -173.915 ;
        RECT -60.005 -176.965 -59.675 -176.635 ;
        RECT -60.005 -178.325 -59.675 -177.995 ;
        RECT -60.005 -180.57 -59.675 -179.44 ;
        RECT -60 -180.685 -59.68 -121.56 ;
    END
    PORT
      LAYER met3 ;
        RECT -58.645 241.32 -58.315 242.45 ;
        RECT -58.645 239.195 -58.315 239.525 ;
        RECT -58.645 237.835 -58.315 238.165 ;
        RECT -58.645 236.475 -58.315 236.805 ;
        RECT -58.645 235.115 -58.315 235.445 ;
        RECT -58.645 233.755 -58.315 234.085 ;
        RECT -58.645 232.395 -58.315 232.725 ;
        RECT -58.645 231.035 -58.315 231.365 ;
        RECT -58.645 229.675 -58.315 230.005 ;
        RECT -58.645 228.315 -58.315 228.645 ;
        RECT -58.645 226.955 -58.315 227.285 ;
        RECT -58.645 225.595 -58.315 225.925 ;
        RECT -58.645 224.235 -58.315 224.565 ;
        RECT -58.645 222.875 -58.315 223.205 ;
        RECT -58.645 221.515 -58.315 221.845 ;
        RECT -58.645 220.155 -58.315 220.485 ;
        RECT -58.645 218.795 -58.315 219.125 ;
        RECT -58.645 217.435 -58.315 217.765 ;
        RECT -58.645 216.075 -58.315 216.405 ;
        RECT -58.645 214.715 -58.315 215.045 ;
        RECT -58.645 213.355 -58.315 213.685 ;
        RECT -58.645 211.995 -58.315 212.325 ;
        RECT -58.645 210.635 -58.315 210.965 ;
        RECT -58.645 209.275 -58.315 209.605 ;
        RECT -58.645 207.915 -58.315 208.245 ;
        RECT -58.645 206.555 -58.315 206.885 ;
        RECT -58.645 205.195 -58.315 205.525 ;
        RECT -58.645 203.835 -58.315 204.165 ;
        RECT -58.645 202.475 -58.315 202.805 ;
        RECT -58.645 201.115 -58.315 201.445 ;
        RECT -58.645 199.755 -58.315 200.085 ;
        RECT -58.645 198.395 -58.315 198.725 ;
        RECT -58.645 197.035 -58.315 197.365 ;
        RECT -58.645 195.675 -58.315 196.005 ;
        RECT -58.645 194.315 -58.315 194.645 ;
        RECT -58.645 192.955 -58.315 193.285 ;
        RECT -58.645 191.595 -58.315 191.925 ;
        RECT -58.645 190.235 -58.315 190.565 ;
        RECT -58.645 188.875 -58.315 189.205 ;
        RECT -58.645 187.515 -58.315 187.845 ;
        RECT -58.645 186.155 -58.315 186.485 ;
        RECT -58.645 184.795 -58.315 185.125 ;
        RECT -58.645 183.435 -58.315 183.765 ;
        RECT -58.645 182.075 -58.315 182.405 ;
        RECT -58.645 180.715 -58.315 181.045 ;
        RECT -58.645 179.355 -58.315 179.685 ;
        RECT -58.645 177.995 -58.315 178.325 ;
        RECT -58.645 176.635 -58.315 176.965 ;
        RECT -58.645 175.275 -58.315 175.605 ;
        RECT -58.645 173.915 -58.315 174.245 ;
        RECT -58.645 172.555 -58.315 172.885 ;
        RECT -58.645 171.195 -58.315 171.525 ;
        RECT -58.645 169.835 -58.315 170.165 ;
        RECT -58.645 168.475 -58.315 168.805 ;
        RECT -58.645 167.115 -58.315 167.445 ;
        RECT -58.645 165.755 -58.315 166.085 ;
        RECT -58.645 164.395 -58.315 164.725 ;
        RECT -58.645 163.035 -58.315 163.365 ;
        RECT -58.645 161.675 -58.315 162.005 ;
        RECT -58.645 160.315 -58.315 160.645 ;
        RECT -58.645 158.955 -58.315 159.285 ;
        RECT -58.645 157.595 -58.315 157.925 ;
        RECT -58.645 156.235 -58.315 156.565 ;
        RECT -58.645 154.875 -58.315 155.205 ;
        RECT -58.645 153.515 -58.315 153.845 ;
        RECT -58.645 152.155 -58.315 152.485 ;
        RECT -58.645 150.795 -58.315 151.125 ;
        RECT -58.645 149.435 -58.315 149.765 ;
        RECT -58.645 148.075 -58.315 148.405 ;
        RECT -58.645 146.715 -58.315 147.045 ;
        RECT -58.645 145.355 -58.315 145.685 ;
        RECT -58.645 143.995 -58.315 144.325 ;
        RECT -58.645 142.635 -58.315 142.965 ;
        RECT -58.645 141.275 -58.315 141.605 ;
        RECT -58.645 139.915 -58.315 140.245 ;
        RECT -58.645 138.555 -58.315 138.885 ;
        RECT -58.64 138.555 -58.32 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -58.645 97.755 -58.315 98.085 ;
        RECT -58.645 96.395 -58.315 96.725 ;
        RECT -58.645 95.035 -58.315 95.365 ;
        RECT -58.645 93.675 -58.315 94.005 ;
        RECT -58.645 92.315 -58.315 92.645 ;
        RECT -58.645 89.595 -58.315 89.925 ;
        RECT -58.645 88.235 -58.315 88.565 ;
        RECT -58.645 84.155 -58.315 84.485 ;
        RECT -58.645 82.795 -58.315 83.125 ;
        RECT -58.645 81.435 -58.315 81.765 ;
        RECT -58.645 80.075 -58.315 80.405 ;
        RECT -58.645 78.715 -58.315 79.045 ;
        RECT -58.645 77.355 -58.315 77.685 ;
        RECT -58.645 75.995 -58.315 76.325 ;
        RECT -58.645 74.635 -58.315 74.965 ;
        RECT -58.645 73.275 -58.315 73.605 ;
        RECT -58.645 71.915 -58.315 72.245 ;
        RECT -58.645 70.555 -58.315 70.885 ;
        RECT -58.645 69.195 -58.315 69.525 ;
        RECT -58.645 67.835 -58.315 68.165 ;
        RECT -58.645 66.475 -58.315 66.805 ;
        RECT -58.645 65.115 -58.315 65.445 ;
        RECT -58.645 63.755 -58.315 64.085 ;
        RECT -58.645 62.395 -58.315 62.725 ;
        RECT -58.645 61.035 -58.315 61.365 ;
        RECT -58.645 59.675 -58.315 60.005 ;
        RECT -58.645 58.315 -58.315 58.645 ;
        RECT -58.645 56.955 -58.315 57.285 ;
        RECT -58.645 55.595 -58.315 55.925 ;
        RECT -58.645 54.235 -58.315 54.565 ;
        RECT -58.645 52.875 -58.315 53.205 ;
        RECT -58.645 51.515 -58.315 51.845 ;
        RECT -58.645 50.155 -58.315 50.485 ;
        RECT -58.645 48.795 -58.315 49.125 ;
        RECT -58.645 47.435 -58.315 47.765 ;
        RECT -58.645 46.075 -58.315 46.405 ;
        RECT -58.645 44.715 -58.315 45.045 ;
        RECT -58.645 43.355 -58.315 43.685 ;
        RECT -58.645 41.995 -58.315 42.325 ;
        RECT -58.645 40.635 -58.315 40.965 ;
        RECT -58.645 39.275 -58.315 39.605 ;
        RECT -58.645 37.915 -58.315 38.245 ;
        RECT -58.645 36.555 -58.315 36.885 ;
        RECT -58.645 35.195 -58.315 35.525 ;
        RECT -58.645 33.835 -58.315 34.165 ;
        RECT -58.645 32.475 -58.315 32.805 ;
        RECT -58.645 31.115 -58.315 31.445 ;
        RECT -58.645 29.755 -58.315 30.085 ;
        RECT -58.645 28.395 -58.315 28.725 ;
        RECT -58.645 27.035 -58.315 27.365 ;
        RECT -58.645 25.675 -58.315 26.005 ;
        RECT -58.645 24.315 -58.315 24.645 ;
        RECT -58.645 22.955 -58.315 23.285 ;
        RECT -58.645 21.595 -58.315 21.925 ;
        RECT -58.645 20.235 -58.315 20.565 ;
        RECT -58.645 18.875 -58.315 19.205 ;
        RECT -58.645 17.515 -58.315 17.845 ;
        RECT -58.645 16.155 -58.315 16.485 ;
        RECT -58.645 14.795 -58.315 15.125 ;
        RECT -58.645 13.435 -58.315 13.765 ;
        RECT -58.645 12.075 -58.315 12.405 ;
        RECT -58.645 10.715 -58.315 11.045 ;
        RECT -58.645 9.355 -58.315 9.685 ;
        RECT -58.645 7.995 -58.315 8.325 ;
        RECT -58.645 6.635 -58.315 6.965 ;
        RECT -58.645 5.275 -58.315 5.605 ;
        RECT -58.645 3.915 -58.315 4.245 ;
        RECT -58.645 2.555 -58.315 2.885 ;
        RECT -58.645 1.195 -58.315 1.525 ;
        RECT -58.645 -0.165 -58.315 0.165 ;
        RECT -58.645 -2.885 -58.315 -2.555 ;
        RECT -58.645 -4.245 -58.315 -3.915 ;
        RECT -58.645 -5.605 -58.315 -5.275 ;
        RECT -58.645 -6.965 -58.315 -6.635 ;
        RECT -58.645 -8.325 -58.315 -7.995 ;
        RECT -58.645 -9.685 -58.315 -9.355 ;
        RECT -58.645 -11.045 -58.315 -10.715 ;
        RECT -58.645 -12.405 -58.315 -12.075 ;
        RECT -58.645 -13.765 -58.315 -13.435 ;
        RECT -58.645 -15.125 -58.315 -14.795 ;
        RECT -58.645 -16.485 -58.315 -16.155 ;
        RECT -58.645 -17.845 -58.315 -17.515 ;
        RECT -58.645 -19.205 -58.315 -18.875 ;
        RECT -58.645 -20.565 -58.315 -20.235 ;
        RECT -58.645 -21.925 -58.315 -21.595 ;
        RECT -58.645 -23.285 -58.315 -22.955 ;
        RECT -58.645 -24.645 -58.315 -24.315 ;
        RECT -58.645 -27.365 -58.315 -27.035 ;
        RECT -58.645 -28.725 -58.315 -28.395 ;
        RECT -58.645 -30.085 -58.315 -29.755 ;
        RECT -58.645 -31.445 -58.315 -31.115 ;
        RECT -58.645 -32.805 -58.315 -32.475 ;
        RECT -58.645 -34.165 -58.315 -33.835 ;
        RECT -58.645 -35.525 -58.315 -35.195 ;
        RECT -58.645 -36.885 -58.315 -36.555 ;
        RECT -58.645 -38.245 -58.315 -37.915 ;
        RECT -58.645 -39.605 -58.315 -39.275 ;
        RECT -58.645 -40.965 -58.315 -40.635 ;
        RECT -58.645 -42.325 -58.315 -41.995 ;
        RECT -58.645 -43.685 -58.315 -43.355 ;
        RECT -58.645 -45.045 -58.315 -44.715 ;
        RECT -58.645 -46.405 -58.315 -46.075 ;
        RECT -58.645 -47.765 -58.315 -47.435 ;
        RECT -58.645 -49.125 -58.315 -48.795 ;
        RECT -58.645 -50.485 -58.315 -50.155 ;
        RECT -58.645 -51.845 -58.315 -51.515 ;
        RECT -58.645 -53.205 -58.315 -52.875 ;
        RECT -58.645 -54.565 -58.315 -54.235 ;
        RECT -58.645 -55.925 -58.315 -55.595 ;
        RECT -58.645 -57.285 -58.315 -56.955 ;
        RECT -58.645 -58.645 -58.315 -58.315 ;
        RECT -58.645 -60.005 -58.315 -59.675 ;
        RECT -58.645 -61.365 -58.315 -61.035 ;
        RECT -58.645 -62.725 -58.315 -62.395 ;
        RECT -58.645 -64.085 -58.315 -63.755 ;
        RECT -58.645 -65.445 -58.315 -65.115 ;
        RECT -58.645 -66.805 -58.315 -66.475 ;
        RECT -58.645 -68.165 -58.315 -67.835 ;
        RECT -58.645 -69.525 -58.315 -69.195 ;
        RECT -58.645 -70.885 -58.315 -70.555 ;
        RECT -58.645 -72.245 -58.315 -71.915 ;
        RECT -58.645 -73.605 -58.315 -73.275 ;
        RECT -58.645 -74.965 -58.315 -74.635 ;
        RECT -58.645 -76.325 -58.315 -75.995 ;
        RECT -58.645 -77.685 -58.315 -77.355 ;
        RECT -58.645 -79.045 -58.315 -78.715 ;
        RECT -58.645 -80.405 -58.315 -80.075 ;
        RECT -58.645 -81.765 -58.315 -81.435 ;
        RECT -58.645 -83.125 -58.315 -82.795 ;
        RECT -58.645 -84.485 -58.315 -84.155 ;
        RECT -58.645 -85.845 -58.315 -85.515 ;
        RECT -58.645 -87.205 -58.315 -86.875 ;
        RECT -58.645 -88.565 -58.315 -88.235 ;
        RECT -58.645 -89.925 -58.315 -89.595 ;
        RECT -58.645 -92.645 -58.315 -92.315 ;
        RECT -58.645 -94.005 -58.315 -93.675 ;
        RECT -58.645 -95.365 -58.315 -95.035 ;
        RECT -58.645 -96.725 -58.315 -96.395 ;
        RECT -58.645 -98.73 -58.315 -98.4 ;
        RECT -58.645 -99.445 -58.315 -99.115 ;
        RECT -58.645 -102.165 -58.315 -101.835 ;
        RECT -58.645 -103.525 -58.315 -103.195 ;
        RECT -58.645 -104.885 -58.315 -104.555 ;
        RECT -58.645 -106.87 -58.315 -106.54 ;
        RECT -58.645 -107.605 -58.315 -107.275 ;
        RECT -58.645 -108.965 -58.315 -108.635 ;
        RECT -58.645 -110.325 -58.315 -109.995 ;
        RECT -58.64 -113.04 -58.32 98.085 ;
    END
    PORT
      LAYER met3 ;
        RECT -57.285 241.32 -56.955 242.45 ;
        RECT -57.285 239.195 -56.955 239.525 ;
        RECT -57.285 237.835 -56.955 238.165 ;
        RECT -57.285 236.475 -56.955 236.805 ;
        RECT -57.285 235.115 -56.955 235.445 ;
        RECT -57.285 233.755 -56.955 234.085 ;
        RECT -57.285 232.395 -56.955 232.725 ;
        RECT -57.285 231.035 -56.955 231.365 ;
        RECT -57.285 229.675 -56.955 230.005 ;
        RECT -57.285 228.315 -56.955 228.645 ;
        RECT -57.285 226.955 -56.955 227.285 ;
        RECT -57.285 225.595 -56.955 225.925 ;
        RECT -57.285 224.235 -56.955 224.565 ;
        RECT -57.285 222.875 -56.955 223.205 ;
        RECT -57.285 221.515 -56.955 221.845 ;
        RECT -57.285 220.155 -56.955 220.485 ;
        RECT -57.285 218.795 -56.955 219.125 ;
        RECT -57.285 217.435 -56.955 217.765 ;
        RECT -57.285 216.075 -56.955 216.405 ;
        RECT -57.285 214.715 -56.955 215.045 ;
        RECT -57.285 213.355 -56.955 213.685 ;
        RECT -57.285 211.995 -56.955 212.325 ;
        RECT -57.285 210.635 -56.955 210.965 ;
        RECT -57.285 209.275 -56.955 209.605 ;
        RECT -57.285 207.915 -56.955 208.245 ;
        RECT -57.285 206.555 -56.955 206.885 ;
        RECT -57.285 205.195 -56.955 205.525 ;
        RECT -57.285 203.835 -56.955 204.165 ;
        RECT -57.285 202.475 -56.955 202.805 ;
        RECT -57.285 201.115 -56.955 201.445 ;
        RECT -57.285 199.755 -56.955 200.085 ;
        RECT -57.285 198.395 -56.955 198.725 ;
        RECT -57.285 197.035 -56.955 197.365 ;
        RECT -57.285 195.675 -56.955 196.005 ;
        RECT -57.285 194.315 -56.955 194.645 ;
        RECT -57.285 192.955 -56.955 193.285 ;
        RECT -57.285 191.595 -56.955 191.925 ;
        RECT -57.285 190.235 -56.955 190.565 ;
        RECT -57.285 188.875 -56.955 189.205 ;
        RECT -57.285 187.515 -56.955 187.845 ;
        RECT -57.285 186.155 -56.955 186.485 ;
        RECT -57.285 184.795 -56.955 185.125 ;
        RECT -57.285 183.435 -56.955 183.765 ;
        RECT -57.285 182.075 -56.955 182.405 ;
        RECT -57.285 180.715 -56.955 181.045 ;
        RECT -57.285 179.355 -56.955 179.685 ;
        RECT -57.285 177.995 -56.955 178.325 ;
        RECT -57.285 176.635 -56.955 176.965 ;
        RECT -57.285 175.275 -56.955 175.605 ;
        RECT -57.285 173.915 -56.955 174.245 ;
        RECT -57.285 172.555 -56.955 172.885 ;
        RECT -57.285 171.195 -56.955 171.525 ;
        RECT -57.285 169.835 -56.955 170.165 ;
        RECT -57.285 168.475 -56.955 168.805 ;
        RECT -57.285 167.115 -56.955 167.445 ;
        RECT -57.285 165.755 -56.955 166.085 ;
        RECT -57.285 164.395 -56.955 164.725 ;
        RECT -57.285 163.035 -56.955 163.365 ;
        RECT -57.285 161.675 -56.955 162.005 ;
        RECT -57.285 160.315 -56.955 160.645 ;
        RECT -57.285 158.955 -56.955 159.285 ;
        RECT -57.285 157.595 -56.955 157.925 ;
        RECT -57.285 156.235 -56.955 156.565 ;
        RECT -57.285 154.875 -56.955 155.205 ;
        RECT -57.285 153.515 -56.955 153.845 ;
        RECT -57.285 152.155 -56.955 152.485 ;
        RECT -57.285 150.795 -56.955 151.125 ;
        RECT -57.285 149.435 -56.955 149.765 ;
        RECT -57.285 148.075 -56.955 148.405 ;
        RECT -57.285 146.715 -56.955 147.045 ;
        RECT -57.285 145.355 -56.955 145.685 ;
        RECT -57.285 143.995 -56.955 144.325 ;
        RECT -57.285 142.635 -56.955 142.965 ;
        RECT -57.285 141.275 -56.955 141.605 ;
        RECT -57.285 139.915 -56.955 140.245 ;
        RECT -57.285 138.555 -56.955 138.885 ;
        RECT -57.28 138.555 -56.96 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -57.285 97.755 -56.955 98.085 ;
        RECT -57.285 96.395 -56.955 96.725 ;
        RECT -57.285 95.035 -56.955 95.365 ;
        RECT -57.285 93.675 -56.955 94.005 ;
        RECT -57.285 92.315 -56.955 92.645 ;
        RECT -57.285 89.595 -56.955 89.925 ;
        RECT -57.285 88.235 -56.955 88.565 ;
        RECT -57.285 84.155 -56.955 84.485 ;
        RECT -57.285 82.795 -56.955 83.125 ;
        RECT -57.285 81.435 -56.955 81.765 ;
        RECT -57.285 80.075 -56.955 80.405 ;
        RECT -57.285 78.715 -56.955 79.045 ;
        RECT -57.285 77.355 -56.955 77.685 ;
        RECT -57.285 75.995 -56.955 76.325 ;
        RECT -57.285 74.635 -56.955 74.965 ;
        RECT -57.285 73.275 -56.955 73.605 ;
        RECT -57.285 71.915 -56.955 72.245 ;
        RECT -57.285 70.555 -56.955 70.885 ;
        RECT -57.285 69.195 -56.955 69.525 ;
        RECT -57.285 67.835 -56.955 68.165 ;
        RECT -57.285 66.475 -56.955 66.805 ;
        RECT -57.285 65.115 -56.955 65.445 ;
        RECT -57.285 63.755 -56.955 64.085 ;
        RECT -57.285 62.395 -56.955 62.725 ;
        RECT -57.285 61.035 -56.955 61.365 ;
        RECT -57.285 59.675 -56.955 60.005 ;
        RECT -57.285 58.315 -56.955 58.645 ;
        RECT -57.285 56.955 -56.955 57.285 ;
        RECT -57.285 55.595 -56.955 55.925 ;
        RECT -57.285 54.235 -56.955 54.565 ;
        RECT -57.285 52.875 -56.955 53.205 ;
        RECT -57.285 51.515 -56.955 51.845 ;
        RECT -57.285 50.155 -56.955 50.485 ;
        RECT -57.285 48.795 -56.955 49.125 ;
        RECT -57.285 47.435 -56.955 47.765 ;
        RECT -57.285 46.075 -56.955 46.405 ;
        RECT -57.285 44.715 -56.955 45.045 ;
        RECT -57.285 43.355 -56.955 43.685 ;
        RECT -57.285 41.995 -56.955 42.325 ;
        RECT -57.285 40.635 -56.955 40.965 ;
        RECT -57.285 39.275 -56.955 39.605 ;
        RECT -57.285 37.915 -56.955 38.245 ;
        RECT -57.285 36.555 -56.955 36.885 ;
        RECT -57.285 35.195 -56.955 35.525 ;
        RECT -57.285 33.835 -56.955 34.165 ;
        RECT -57.285 32.475 -56.955 32.805 ;
        RECT -57.285 31.115 -56.955 31.445 ;
        RECT -57.285 29.755 -56.955 30.085 ;
        RECT -57.285 28.395 -56.955 28.725 ;
        RECT -57.285 27.035 -56.955 27.365 ;
        RECT -57.285 25.675 -56.955 26.005 ;
        RECT -57.285 24.315 -56.955 24.645 ;
        RECT -57.285 22.955 -56.955 23.285 ;
        RECT -57.285 21.595 -56.955 21.925 ;
        RECT -57.285 20.235 -56.955 20.565 ;
        RECT -57.285 18.875 -56.955 19.205 ;
        RECT -57.285 17.515 -56.955 17.845 ;
        RECT -57.285 16.155 -56.955 16.485 ;
        RECT -57.285 14.795 -56.955 15.125 ;
        RECT -57.285 13.435 -56.955 13.765 ;
        RECT -57.285 12.075 -56.955 12.405 ;
        RECT -57.285 10.715 -56.955 11.045 ;
        RECT -57.285 9.355 -56.955 9.685 ;
        RECT -57.285 7.995 -56.955 8.325 ;
        RECT -57.285 6.635 -56.955 6.965 ;
        RECT -57.285 5.275 -56.955 5.605 ;
        RECT -57.285 3.915 -56.955 4.245 ;
        RECT -57.285 2.555 -56.955 2.885 ;
        RECT -57.285 1.195 -56.955 1.525 ;
        RECT -57.285 -0.165 -56.955 0.165 ;
        RECT -57.285 -2.885 -56.955 -2.555 ;
        RECT -57.285 -4.245 -56.955 -3.915 ;
        RECT -57.285 -5.605 -56.955 -5.275 ;
        RECT -57.285 -6.965 -56.955 -6.635 ;
        RECT -57.285 -8.325 -56.955 -7.995 ;
        RECT -57.285 -9.685 -56.955 -9.355 ;
        RECT -57.285 -11.045 -56.955 -10.715 ;
        RECT -57.285 -12.405 -56.955 -12.075 ;
        RECT -57.285 -13.765 -56.955 -13.435 ;
        RECT -57.285 -15.125 -56.955 -14.795 ;
        RECT -57.285 -16.485 -56.955 -16.155 ;
        RECT -57.285 -17.845 -56.955 -17.515 ;
        RECT -57.285 -19.205 -56.955 -18.875 ;
        RECT -57.285 -20.565 -56.955 -20.235 ;
        RECT -57.285 -21.925 -56.955 -21.595 ;
        RECT -57.285 -23.285 -56.955 -22.955 ;
        RECT -57.285 -24.645 -56.955 -24.315 ;
        RECT -57.285 -27.365 -56.955 -27.035 ;
        RECT -57.285 -28.725 -56.955 -28.395 ;
        RECT -57.285 -30.085 -56.955 -29.755 ;
        RECT -57.285 -31.445 -56.955 -31.115 ;
        RECT -57.285 -32.805 -56.955 -32.475 ;
        RECT -57.285 -34.165 -56.955 -33.835 ;
        RECT -57.285 -35.525 -56.955 -35.195 ;
        RECT -57.285 -36.885 -56.955 -36.555 ;
        RECT -57.285 -38.245 -56.955 -37.915 ;
        RECT -57.285 -39.605 -56.955 -39.275 ;
        RECT -57.285 -40.965 -56.955 -40.635 ;
        RECT -57.285 -42.325 -56.955 -41.995 ;
        RECT -57.285 -43.685 -56.955 -43.355 ;
        RECT -57.285 -45.045 -56.955 -44.715 ;
        RECT -57.285 -46.405 -56.955 -46.075 ;
        RECT -57.285 -47.765 -56.955 -47.435 ;
        RECT -57.285 -49.125 -56.955 -48.795 ;
        RECT -57.285 -50.485 -56.955 -50.155 ;
        RECT -57.285 -51.845 -56.955 -51.515 ;
        RECT -57.285 -53.205 -56.955 -52.875 ;
        RECT -57.285 -54.565 -56.955 -54.235 ;
        RECT -57.285 -55.925 -56.955 -55.595 ;
        RECT -57.285 -57.285 -56.955 -56.955 ;
        RECT -57.285 -58.645 -56.955 -58.315 ;
        RECT -57.285 -60.005 -56.955 -59.675 ;
        RECT -57.285 -61.365 -56.955 -61.035 ;
        RECT -57.285 -62.725 -56.955 -62.395 ;
        RECT -57.285 -64.085 -56.955 -63.755 ;
        RECT -57.285 -65.445 -56.955 -65.115 ;
        RECT -57.285 -66.805 -56.955 -66.475 ;
        RECT -57.285 -68.165 -56.955 -67.835 ;
        RECT -57.285 -69.525 -56.955 -69.195 ;
        RECT -57.285 -70.885 -56.955 -70.555 ;
        RECT -57.285 -72.245 -56.955 -71.915 ;
        RECT -57.285 -73.605 -56.955 -73.275 ;
        RECT -57.285 -74.965 -56.955 -74.635 ;
        RECT -57.285 -76.325 -56.955 -75.995 ;
        RECT -57.285 -77.685 -56.955 -77.355 ;
        RECT -57.285 -79.045 -56.955 -78.715 ;
        RECT -57.285 -80.405 -56.955 -80.075 ;
        RECT -57.285 -81.765 -56.955 -81.435 ;
        RECT -57.285 -83.125 -56.955 -82.795 ;
        RECT -57.285 -84.485 -56.955 -84.155 ;
        RECT -57.285 -85.845 -56.955 -85.515 ;
        RECT -57.285 -87.205 -56.955 -86.875 ;
        RECT -57.285 -88.565 -56.955 -88.235 ;
        RECT -57.285 -89.925 -56.955 -89.595 ;
        RECT -57.285 -92.645 -56.955 -92.315 ;
        RECT -57.285 -94.005 -56.955 -93.675 ;
        RECT -57.285 -95.365 -56.955 -95.035 ;
        RECT -57.285 -96.725 -56.955 -96.395 ;
        RECT -57.285 -98.73 -56.955 -98.4 ;
        RECT -57.285 -99.445 -56.955 -99.115 ;
        RECT -57.285 -102.165 -56.955 -101.835 ;
        RECT -57.285 -103.525 -56.955 -103.195 ;
        RECT -57.285 -104.885 -56.955 -104.555 ;
        RECT -57.285 -106.87 -56.955 -106.54 ;
        RECT -57.285 -107.605 -56.955 -107.275 ;
        RECT -57.285 -108.965 -56.955 -108.635 ;
        RECT -57.285 -110.325 -56.955 -109.995 ;
        RECT -57.285 -113.045 -56.955 -112.715 ;
        RECT -57.285 -115.765 -56.955 -115.435 ;
        RECT -57.285 -117.125 -56.955 -116.795 ;
        RECT -57.285 -118.485 -56.955 -118.155 ;
        RECT -57.285 -122.565 -56.955 -122.235 ;
        RECT -57.285 -123.925 -56.955 -123.595 ;
        RECT -57.285 -125.285 -56.955 -124.955 ;
        RECT -57.285 -126.645 -56.955 -126.315 ;
        RECT -57.285 -128.005 -56.955 -127.675 ;
        RECT -57.285 -129.365 -56.955 -129.035 ;
        RECT -57.285 -130.725 -56.955 -130.395 ;
        RECT -57.285 -132.085 -56.955 -131.755 ;
        RECT -57.285 -133.445 -56.955 -133.115 ;
        RECT -57.285 -134.805 -56.955 -134.475 ;
        RECT -57.285 -136.165 -56.955 -135.835 ;
        RECT -57.285 -137.525 -56.955 -137.195 ;
        RECT -57.285 -138.885 -56.955 -138.555 ;
        RECT -57.285 -140.245 -56.955 -139.915 ;
        RECT -57.285 -141.605 -56.955 -141.275 ;
        RECT -57.285 -142.965 -56.955 -142.635 ;
        RECT -57.285 -144.325 -56.955 -143.995 ;
        RECT -57.285 -145.685 -56.955 -145.355 ;
        RECT -57.285 -147.045 -56.955 -146.715 ;
        RECT -57.285 -148.405 -56.955 -148.075 ;
        RECT -57.285 -149.765 -56.955 -149.435 ;
        RECT -57.285 -151.125 -56.955 -150.795 ;
        RECT -57.285 -152.485 -56.955 -152.155 ;
        RECT -57.285 -153.845 -56.955 -153.515 ;
        RECT -57.285 -155.205 -56.955 -154.875 ;
        RECT -57.285 -156.565 -56.955 -156.235 ;
        RECT -57.285 -157.925 -56.955 -157.595 ;
        RECT -57.285 -159.285 -56.955 -158.955 ;
        RECT -57.285 -160.645 -56.955 -160.315 ;
        RECT -57.285 -162.005 -56.955 -161.675 ;
        RECT -57.285 -163.365 -56.955 -163.035 ;
        RECT -57.285 -164.725 -56.955 -164.395 ;
        RECT -57.285 -166.085 -56.955 -165.755 ;
        RECT -57.285 -167.445 -56.955 -167.115 ;
        RECT -57.285 -170.165 -56.955 -169.835 ;
        RECT -57.285 -172.885 -56.955 -172.555 ;
        RECT -57.285 -174.245 -56.955 -173.915 ;
        RECT -57.285 -175.725 -56.955 -175.395 ;
        RECT -57.285 -176.965 -56.955 -176.635 ;
        RECT -57.285 -178.325 -56.955 -177.995 ;
        RECT -57.285 -180.57 -56.955 -179.44 ;
        RECT -57.28 -180.685 -56.96 98.085 ;
    END
    PORT
      LAYER met3 ;
        RECT -55.925 241.32 -55.595 242.45 ;
        RECT -55.925 239.195 -55.595 239.525 ;
        RECT -55.925 237.835 -55.595 238.165 ;
        RECT -55.925 236.475 -55.595 236.805 ;
        RECT -55.925 235.115 -55.595 235.445 ;
        RECT -55.925 233.755 -55.595 234.085 ;
        RECT -55.925 232.395 -55.595 232.725 ;
        RECT -55.925 231.035 -55.595 231.365 ;
        RECT -55.925 229.675 -55.595 230.005 ;
        RECT -55.925 228.315 -55.595 228.645 ;
        RECT -55.925 226.955 -55.595 227.285 ;
        RECT -55.925 225.595 -55.595 225.925 ;
        RECT -55.925 224.235 -55.595 224.565 ;
        RECT -55.925 222.875 -55.595 223.205 ;
        RECT -55.925 221.515 -55.595 221.845 ;
        RECT -55.925 220.155 -55.595 220.485 ;
        RECT -55.925 218.795 -55.595 219.125 ;
        RECT -55.925 217.435 -55.595 217.765 ;
        RECT -55.925 216.075 -55.595 216.405 ;
        RECT -55.925 214.715 -55.595 215.045 ;
        RECT -55.925 213.355 -55.595 213.685 ;
        RECT -55.925 211.995 -55.595 212.325 ;
        RECT -55.925 210.635 -55.595 210.965 ;
        RECT -55.925 209.275 -55.595 209.605 ;
        RECT -55.925 207.915 -55.595 208.245 ;
        RECT -55.925 206.555 -55.595 206.885 ;
        RECT -55.925 205.195 -55.595 205.525 ;
        RECT -55.925 203.835 -55.595 204.165 ;
        RECT -55.925 202.475 -55.595 202.805 ;
        RECT -55.925 201.115 -55.595 201.445 ;
        RECT -55.925 199.755 -55.595 200.085 ;
        RECT -55.925 198.395 -55.595 198.725 ;
        RECT -55.925 197.035 -55.595 197.365 ;
        RECT -55.925 195.675 -55.595 196.005 ;
        RECT -55.925 194.315 -55.595 194.645 ;
        RECT -55.925 192.955 -55.595 193.285 ;
        RECT -55.925 191.595 -55.595 191.925 ;
        RECT -55.925 190.235 -55.595 190.565 ;
        RECT -55.925 188.875 -55.595 189.205 ;
        RECT -55.925 187.515 -55.595 187.845 ;
        RECT -55.925 186.155 -55.595 186.485 ;
        RECT -55.925 184.795 -55.595 185.125 ;
        RECT -55.925 183.435 -55.595 183.765 ;
        RECT -55.925 182.075 -55.595 182.405 ;
        RECT -55.925 180.715 -55.595 181.045 ;
        RECT -55.925 179.355 -55.595 179.685 ;
        RECT -55.925 177.995 -55.595 178.325 ;
        RECT -55.925 176.635 -55.595 176.965 ;
        RECT -55.925 175.275 -55.595 175.605 ;
        RECT -55.925 173.915 -55.595 174.245 ;
        RECT -55.925 172.555 -55.595 172.885 ;
        RECT -55.925 171.195 -55.595 171.525 ;
        RECT -55.925 169.835 -55.595 170.165 ;
        RECT -55.925 168.475 -55.595 168.805 ;
        RECT -55.925 167.115 -55.595 167.445 ;
        RECT -55.925 165.755 -55.595 166.085 ;
        RECT -55.925 164.395 -55.595 164.725 ;
        RECT -55.925 163.035 -55.595 163.365 ;
        RECT -55.925 161.675 -55.595 162.005 ;
        RECT -55.925 160.315 -55.595 160.645 ;
        RECT -55.925 158.955 -55.595 159.285 ;
        RECT -55.925 157.595 -55.595 157.925 ;
        RECT -55.925 156.235 -55.595 156.565 ;
        RECT -55.925 154.875 -55.595 155.205 ;
        RECT -55.925 153.515 -55.595 153.845 ;
        RECT -55.925 152.155 -55.595 152.485 ;
        RECT -55.925 150.795 -55.595 151.125 ;
        RECT -55.925 149.435 -55.595 149.765 ;
        RECT -55.925 148.075 -55.595 148.405 ;
        RECT -55.925 146.715 -55.595 147.045 ;
        RECT -55.925 145.355 -55.595 145.685 ;
        RECT -55.925 143.995 -55.595 144.325 ;
        RECT -55.925 142.635 -55.595 142.965 ;
        RECT -55.925 141.275 -55.595 141.605 ;
        RECT -55.925 139.915 -55.595 140.245 ;
        RECT -55.925 138.555 -55.595 138.885 ;
        RECT -55.92 138.555 -55.6 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -55.925 97.755 -55.595 98.085 ;
        RECT -55.925 96.395 -55.595 96.725 ;
        RECT -55.925 95.035 -55.595 95.365 ;
        RECT -55.925 93.675 -55.595 94.005 ;
        RECT -55.925 92.315 -55.595 92.645 ;
        RECT -55.925 89.595 -55.595 89.925 ;
        RECT -55.925 88.235 -55.595 88.565 ;
        RECT -55.925 84.155 -55.595 84.485 ;
        RECT -55.925 82.795 -55.595 83.125 ;
        RECT -55.925 81.435 -55.595 81.765 ;
        RECT -55.925 80.075 -55.595 80.405 ;
        RECT -55.925 78.715 -55.595 79.045 ;
        RECT -55.925 77.355 -55.595 77.685 ;
        RECT -55.925 75.995 -55.595 76.325 ;
        RECT -55.925 74.635 -55.595 74.965 ;
        RECT -55.925 73.275 -55.595 73.605 ;
        RECT -55.925 71.915 -55.595 72.245 ;
        RECT -55.925 70.555 -55.595 70.885 ;
        RECT -55.925 69.195 -55.595 69.525 ;
        RECT -55.925 67.835 -55.595 68.165 ;
        RECT -55.925 66.475 -55.595 66.805 ;
        RECT -55.925 65.115 -55.595 65.445 ;
        RECT -55.925 63.755 -55.595 64.085 ;
        RECT -55.925 62.395 -55.595 62.725 ;
        RECT -55.925 61.035 -55.595 61.365 ;
        RECT -55.925 59.675 -55.595 60.005 ;
        RECT -55.925 58.315 -55.595 58.645 ;
        RECT -55.925 56.955 -55.595 57.285 ;
        RECT -55.925 55.595 -55.595 55.925 ;
        RECT -55.925 54.235 -55.595 54.565 ;
        RECT -55.925 52.875 -55.595 53.205 ;
        RECT -55.925 51.515 -55.595 51.845 ;
        RECT -55.925 50.155 -55.595 50.485 ;
        RECT -55.925 48.795 -55.595 49.125 ;
        RECT -55.925 47.435 -55.595 47.765 ;
        RECT -55.925 46.075 -55.595 46.405 ;
        RECT -55.925 44.715 -55.595 45.045 ;
        RECT -55.925 43.355 -55.595 43.685 ;
        RECT -55.925 41.995 -55.595 42.325 ;
        RECT -55.925 40.635 -55.595 40.965 ;
        RECT -55.925 39.275 -55.595 39.605 ;
        RECT -55.925 37.915 -55.595 38.245 ;
        RECT -55.925 36.555 -55.595 36.885 ;
        RECT -55.925 35.195 -55.595 35.525 ;
        RECT -55.925 33.835 -55.595 34.165 ;
        RECT -55.925 32.475 -55.595 32.805 ;
        RECT -55.925 31.115 -55.595 31.445 ;
        RECT -55.925 29.755 -55.595 30.085 ;
        RECT -55.925 28.395 -55.595 28.725 ;
        RECT -55.925 27.035 -55.595 27.365 ;
        RECT -55.925 25.675 -55.595 26.005 ;
        RECT -55.925 24.315 -55.595 24.645 ;
        RECT -55.925 22.955 -55.595 23.285 ;
        RECT -55.925 21.595 -55.595 21.925 ;
        RECT -55.925 20.235 -55.595 20.565 ;
        RECT -55.925 18.875 -55.595 19.205 ;
        RECT -55.925 17.515 -55.595 17.845 ;
        RECT -55.925 16.155 -55.595 16.485 ;
        RECT -55.925 14.795 -55.595 15.125 ;
        RECT -55.925 13.435 -55.595 13.765 ;
        RECT -55.925 12.075 -55.595 12.405 ;
        RECT -55.925 10.715 -55.595 11.045 ;
        RECT -55.925 9.355 -55.595 9.685 ;
        RECT -55.925 7.995 -55.595 8.325 ;
        RECT -55.925 6.635 -55.595 6.965 ;
        RECT -55.925 5.275 -55.595 5.605 ;
        RECT -55.925 3.915 -55.595 4.245 ;
        RECT -55.925 2.555 -55.595 2.885 ;
        RECT -55.925 1.195 -55.595 1.525 ;
        RECT -55.925 -0.165 -55.595 0.165 ;
        RECT -55.925 -2.885 -55.595 -2.555 ;
        RECT -55.925 -4.245 -55.595 -3.915 ;
        RECT -55.925 -5.605 -55.595 -5.275 ;
        RECT -55.925 -6.965 -55.595 -6.635 ;
        RECT -55.925 -8.325 -55.595 -7.995 ;
        RECT -55.925 -9.685 -55.595 -9.355 ;
        RECT -55.925 -11.045 -55.595 -10.715 ;
        RECT -55.925 -12.405 -55.595 -12.075 ;
        RECT -55.925 -13.765 -55.595 -13.435 ;
        RECT -55.925 -15.125 -55.595 -14.795 ;
        RECT -55.925 -16.485 -55.595 -16.155 ;
        RECT -55.925 -17.845 -55.595 -17.515 ;
        RECT -55.925 -19.205 -55.595 -18.875 ;
        RECT -55.925 -20.565 -55.595 -20.235 ;
        RECT -55.925 -21.925 -55.595 -21.595 ;
        RECT -55.925 -23.285 -55.595 -22.955 ;
        RECT -55.925 -24.645 -55.595 -24.315 ;
        RECT -55.925 -27.365 -55.595 -27.035 ;
        RECT -55.925 -28.725 -55.595 -28.395 ;
        RECT -55.925 -30.085 -55.595 -29.755 ;
        RECT -55.925 -31.445 -55.595 -31.115 ;
        RECT -55.925 -32.805 -55.595 -32.475 ;
        RECT -55.925 -34.165 -55.595 -33.835 ;
        RECT -55.925 -35.525 -55.595 -35.195 ;
        RECT -55.925 -36.885 -55.595 -36.555 ;
        RECT -55.925 -38.245 -55.595 -37.915 ;
        RECT -55.925 -39.605 -55.595 -39.275 ;
        RECT -55.925 -40.965 -55.595 -40.635 ;
        RECT -55.925 -42.325 -55.595 -41.995 ;
        RECT -55.925 -43.685 -55.595 -43.355 ;
        RECT -55.925 -45.045 -55.595 -44.715 ;
        RECT -55.925 -46.405 -55.595 -46.075 ;
        RECT -55.925 -47.765 -55.595 -47.435 ;
        RECT -55.925 -49.125 -55.595 -48.795 ;
        RECT -55.925 -50.485 -55.595 -50.155 ;
        RECT -55.925 -51.845 -55.595 -51.515 ;
        RECT -55.925 -53.205 -55.595 -52.875 ;
        RECT -55.925 -54.565 -55.595 -54.235 ;
        RECT -55.925 -55.925 -55.595 -55.595 ;
        RECT -55.925 -57.285 -55.595 -56.955 ;
        RECT -55.925 -58.645 -55.595 -58.315 ;
        RECT -55.925 -60.005 -55.595 -59.675 ;
        RECT -55.925 -61.365 -55.595 -61.035 ;
        RECT -55.925 -62.725 -55.595 -62.395 ;
        RECT -55.925 -64.085 -55.595 -63.755 ;
        RECT -55.925 -65.445 -55.595 -65.115 ;
        RECT -55.925 -66.805 -55.595 -66.475 ;
        RECT -55.925 -68.165 -55.595 -67.835 ;
        RECT -55.925 -69.525 -55.595 -69.195 ;
        RECT -55.925 -70.885 -55.595 -70.555 ;
        RECT -55.925 -72.245 -55.595 -71.915 ;
        RECT -55.925 -73.605 -55.595 -73.275 ;
        RECT -55.925 -74.965 -55.595 -74.635 ;
        RECT -55.925 -76.325 -55.595 -75.995 ;
        RECT -55.925 -77.685 -55.595 -77.355 ;
        RECT -55.925 -79.045 -55.595 -78.715 ;
        RECT -55.925 -80.405 -55.595 -80.075 ;
        RECT -55.925 -81.765 -55.595 -81.435 ;
        RECT -55.925 -83.125 -55.595 -82.795 ;
        RECT -55.925 -84.485 -55.595 -84.155 ;
        RECT -55.925 -85.845 -55.595 -85.515 ;
        RECT -55.925 -87.205 -55.595 -86.875 ;
        RECT -55.925 -88.565 -55.595 -88.235 ;
        RECT -55.925 -89.925 -55.595 -89.595 ;
        RECT -55.925 -92.645 -55.595 -92.315 ;
        RECT -55.925 -94.005 -55.595 -93.675 ;
        RECT -55.925 -95.365 -55.595 -95.035 ;
        RECT -55.925 -96.725 -55.595 -96.395 ;
        RECT -55.925 -98.73 -55.595 -98.4 ;
        RECT -55.925 -99.445 -55.595 -99.115 ;
        RECT -55.925 -102.165 -55.595 -101.835 ;
        RECT -55.925 -103.525 -55.595 -103.195 ;
        RECT -55.925 -104.885 -55.595 -104.555 ;
        RECT -55.925 -106.87 -55.595 -106.54 ;
        RECT -55.925 -107.605 -55.595 -107.275 ;
        RECT -55.925 -108.965 -55.595 -108.635 ;
        RECT -55.925 -110.325 -55.595 -109.995 ;
        RECT -55.925 -113.045 -55.595 -112.715 ;
        RECT -55.925 -115.765 -55.595 -115.435 ;
        RECT -55.925 -117.125 -55.595 -116.795 ;
        RECT -55.925 -118.485 -55.595 -118.155 ;
        RECT -55.925 -122.565 -55.595 -122.235 ;
        RECT -55.925 -123.925 -55.595 -123.595 ;
        RECT -55.925 -125.285 -55.595 -124.955 ;
        RECT -55.925 -126.645 -55.595 -126.315 ;
        RECT -55.925 -128.005 -55.595 -127.675 ;
        RECT -55.925 -129.365 -55.595 -129.035 ;
        RECT -55.925 -130.725 -55.595 -130.395 ;
        RECT -55.925 -132.085 -55.595 -131.755 ;
        RECT -55.925 -133.445 -55.595 -133.115 ;
        RECT -55.925 -134.805 -55.595 -134.475 ;
        RECT -55.925 -136.165 -55.595 -135.835 ;
        RECT -55.925 -137.525 -55.595 -137.195 ;
        RECT -55.925 -138.885 -55.595 -138.555 ;
        RECT -55.925 -140.245 -55.595 -139.915 ;
        RECT -55.925 -141.605 -55.595 -141.275 ;
        RECT -55.925 -142.965 -55.595 -142.635 ;
        RECT -55.925 -144.325 -55.595 -143.995 ;
        RECT -55.925 -145.685 -55.595 -145.355 ;
        RECT -55.925 -147.045 -55.595 -146.715 ;
        RECT -55.925 -148.405 -55.595 -148.075 ;
        RECT -55.925 -149.765 -55.595 -149.435 ;
        RECT -55.925 -151.125 -55.595 -150.795 ;
        RECT -55.925 -152.485 -55.595 -152.155 ;
        RECT -55.925 -153.845 -55.595 -153.515 ;
        RECT -55.925 -155.205 -55.595 -154.875 ;
        RECT -55.925 -156.565 -55.595 -156.235 ;
        RECT -55.925 -157.925 -55.595 -157.595 ;
        RECT -55.925 -159.285 -55.595 -158.955 ;
        RECT -55.925 -160.645 -55.595 -160.315 ;
        RECT -55.925 -162.005 -55.595 -161.675 ;
        RECT -55.925 -163.365 -55.595 -163.035 ;
        RECT -55.925 -164.725 -55.595 -164.395 ;
        RECT -55.925 -166.085 -55.595 -165.755 ;
        RECT -55.925 -167.445 -55.595 -167.115 ;
        RECT -55.925 -170.165 -55.595 -169.835 ;
        RECT -55.925 -172.885 -55.595 -172.555 ;
        RECT -55.925 -174.245 -55.595 -173.915 ;
        RECT -55.925 -175.725 -55.595 -175.395 ;
        RECT -55.925 -176.965 -55.595 -176.635 ;
        RECT -55.925 -178.325 -55.595 -177.995 ;
        RECT -55.925 -180.57 -55.595 -179.44 ;
        RECT -55.92 -180.685 -55.6 98.085 ;
    END
    PORT
      LAYER met3 ;
        RECT -54.565 195.675 -54.235 196.005 ;
        RECT -54.565 194.315 -54.235 194.645 ;
        RECT -54.565 192.955 -54.235 193.285 ;
        RECT -54.565 191.595 -54.235 191.925 ;
        RECT -54.565 190.235 -54.235 190.565 ;
        RECT -54.565 188.875 -54.235 189.205 ;
        RECT -54.565 187.515 -54.235 187.845 ;
        RECT -54.565 186.155 -54.235 186.485 ;
        RECT -54.565 184.795 -54.235 185.125 ;
        RECT -54.565 183.435 -54.235 183.765 ;
        RECT -54.565 182.075 -54.235 182.405 ;
        RECT -54.565 180.715 -54.235 181.045 ;
        RECT -54.565 179.355 -54.235 179.685 ;
        RECT -54.565 177.995 -54.235 178.325 ;
        RECT -54.565 176.635 -54.235 176.965 ;
        RECT -54.565 175.275 -54.235 175.605 ;
        RECT -54.565 173.915 -54.235 174.245 ;
        RECT -54.565 172.555 -54.235 172.885 ;
        RECT -54.565 171.195 -54.235 171.525 ;
        RECT -54.565 169.835 -54.235 170.165 ;
        RECT -54.565 168.475 -54.235 168.805 ;
        RECT -54.565 167.115 -54.235 167.445 ;
        RECT -54.565 165.755 -54.235 166.085 ;
        RECT -54.565 164.395 -54.235 164.725 ;
        RECT -54.565 163.035 -54.235 163.365 ;
        RECT -54.565 161.675 -54.235 162.005 ;
        RECT -54.565 160.315 -54.235 160.645 ;
        RECT -54.565 158.955 -54.235 159.285 ;
        RECT -54.565 157.595 -54.235 157.925 ;
        RECT -54.565 156.235 -54.235 156.565 ;
        RECT -54.565 154.875 -54.235 155.205 ;
        RECT -54.565 153.515 -54.235 153.845 ;
        RECT -54.565 152.155 -54.235 152.485 ;
        RECT -54.565 150.795 -54.235 151.125 ;
        RECT -54.565 149.435 -54.235 149.765 ;
        RECT -54.565 148.075 -54.235 148.405 ;
        RECT -54.565 146.715 -54.235 147.045 ;
        RECT -54.565 145.355 -54.235 145.685 ;
        RECT -54.565 143.995 -54.235 144.325 ;
        RECT -54.565 142.635 -54.235 142.965 ;
        RECT -54.565 141.275 -54.235 141.605 ;
        RECT -54.565 139.915 -54.235 140.245 ;
        RECT -54.565 138.555 -54.235 138.885 ;
        RECT -54.56 138.555 -54.24 242.565 ;
        RECT -54.565 241.32 -54.235 242.45 ;
        RECT -54.565 239.195 -54.235 239.525 ;
        RECT -54.565 237.835 -54.235 238.165 ;
        RECT -54.565 236.475 -54.235 236.805 ;
        RECT -54.565 235.115 -54.235 235.445 ;
        RECT -54.565 233.755 -54.235 234.085 ;
        RECT -54.565 232.395 -54.235 232.725 ;
        RECT -54.565 231.035 -54.235 231.365 ;
        RECT -54.565 229.675 -54.235 230.005 ;
        RECT -54.565 228.315 -54.235 228.645 ;
        RECT -54.565 226.955 -54.235 227.285 ;
        RECT -54.565 225.595 -54.235 225.925 ;
        RECT -54.565 224.235 -54.235 224.565 ;
        RECT -54.565 222.875 -54.235 223.205 ;
        RECT -54.565 221.515 -54.235 221.845 ;
        RECT -54.565 220.155 -54.235 220.485 ;
        RECT -54.565 218.795 -54.235 219.125 ;
        RECT -54.565 217.435 -54.235 217.765 ;
        RECT -54.565 216.075 -54.235 216.405 ;
        RECT -54.565 214.715 -54.235 215.045 ;
        RECT -54.565 213.355 -54.235 213.685 ;
        RECT -54.565 211.995 -54.235 212.325 ;
        RECT -54.565 210.635 -54.235 210.965 ;
        RECT -54.565 209.275 -54.235 209.605 ;
        RECT -54.565 207.915 -54.235 208.245 ;
        RECT -54.565 206.555 -54.235 206.885 ;
        RECT -54.565 205.195 -54.235 205.525 ;
        RECT -54.565 203.835 -54.235 204.165 ;
        RECT -54.565 202.475 -54.235 202.805 ;
        RECT -54.565 201.115 -54.235 201.445 ;
        RECT -54.565 199.755 -54.235 200.085 ;
        RECT -54.565 198.395 -54.235 198.725 ;
        RECT -54.565 197.035 -54.235 197.365 ;
    END
    PORT
      LAYER met3 ;
        RECT -64.085 241.32 -63.755 242.45 ;
        RECT -64.085 239.195 -63.755 239.525 ;
        RECT -64.085 237.835 -63.755 238.165 ;
        RECT -64.085 236.475 -63.755 236.805 ;
        RECT -64.085 235.115 -63.755 235.445 ;
        RECT -64.085 233.755 -63.755 234.085 ;
        RECT -64.085 232.395 -63.755 232.725 ;
        RECT -64.085 231.035 -63.755 231.365 ;
        RECT -64.085 229.675 -63.755 230.005 ;
        RECT -64.085 228.315 -63.755 228.645 ;
        RECT -64.085 226.955 -63.755 227.285 ;
        RECT -64.085 225.595 -63.755 225.925 ;
        RECT -64.085 224.235 -63.755 224.565 ;
        RECT -64.085 222.875 -63.755 223.205 ;
        RECT -64.085 221.515 -63.755 221.845 ;
        RECT -64.085 220.155 -63.755 220.485 ;
        RECT -64.085 218.795 -63.755 219.125 ;
        RECT -64.085 217.435 -63.755 217.765 ;
        RECT -64.085 216.075 -63.755 216.405 ;
        RECT -64.085 214.715 -63.755 215.045 ;
        RECT -64.085 213.355 -63.755 213.685 ;
        RECT -64.085 211.995 -63.755 212.325 ;
        RECT -64.085 210.635 -63.755 210.965 ;
        RECT -64.085 209.275 -63.755 209.605 ;
        RECT -64.085 207.915 -63.755 208.245 ;
        RECT -64.085 206.555 -63.755 206.885 ;
        RECT -64.085 205.195 -63.755 205.525 ;
        RECT -64.085 203.835 -63.755 204.165 ;
        RECT -64.085 202.475 -63.755 202.805 ;
        RECT -64.085 201.115 -63.755 201.445 ;
        RECT -64.085 199.755 -63.755 200.085 ;
        RECT -64.085 198.395 -63.755 198.725 ;
        RECT -64.085 197.035 -63.755 197.365 ;
        RECT -64.085 195.675 -63.755 196.005 ;
        RECT -64.085 194.315 -63.755 194.645 ;
        RECT -64.085 192.955 -63.755 193.285 ;
        RECT -64.085 191.595 -63.755 191.925 ;
        RECT -64.085 190.235 -63.755 190.565 ;
        RECT -64.085 188.875 -63.755 189.205 ;
        RECT -64.085 187.515 -63.755 187.845 ;
        RECT -64.085 186.155 -63.755 186.485 ;
        RECT -64.085 184.795 -63.755 185.125 ;
        RECT -64.085 183.435 -63.755 183.765 ;
        RECT -64.085 182.075 -63.755 182.405 ;
        RECT -64.085 180.715 -63.755 181.045 ;
        RECT -64.085 179.355 -63.755 179.685 ;
        RECT -64.085 177.995 -63.755 178.325 ;
        RECT -64.085 176.635 -63.755 176.965 ;
        RECT -64.085 175.275 -63.755 175.605 ;
        RECT -64.085 173.915 -63.755 174.245 ;
        RECT -64.085 172.555 -63.755 172.885 ;
        RECT -64.085 171.195 -63.755 171.525 ;
        RECT -64.085 169.835 -63.755 170.165 ;
        RECT -64.085 168.475 -63.755 168.805 ;
        RECT -64.085 167.115 -63.755 167.445 ;
        RECT -64.085 165.755 -63.755 166.085 ;
        RECT -64.085 164.395 -63.755 164.725 ;
        RECT -64.085 163.035 -63.755 163.365 ;
        RECT -64.085 161.675 -63.755 162.005 ;
        RECT -64.085 160.315 -63.755 160.645 ;
        RECT -64.085 158.955 -63.755 159.285 ;
        RECT -64.085 157.595 -63.755 157.925 ;
        RECT -64.085 156.235 -63.755 156.565 ;
        RECT -64.085 154.875 -63.755 155.205 ;
        RECT -64.085 153.515 -63.755 153.845 ;
        RECT -64.085 152.155 -63.755 152.485 ;
        RECT -64.085 150.795 -63.755 151.125 ;
        RECT -64.085 149.435 -63.755 149.765 ;
        RECT -64.085 148.075 -63.755 148.405 ;
        RECT -64.085 146.715 -63.755 147.045 ;
        RECT -64.085 145.355 -63.755 145.685 ;
        RECT -64.085 143.995 -63.755 144.325 ;
        RECT -64.085 142.635 -63.755 142.965 ;
        RECT -64.085 141.275 -63.755 141.605 ;
        RECT -64.085 139.915 -63.755 140.245 ;
        RECT -64.085 138.555 -63.755 138.885 ;
        RECT -64.085 137.225 -63.755 137.555 ;
        RECT -64.085 135.175 -63.755 135.505 ;
        RECT -64.085 132.815 -63.755 133.145 ;
        RECT -64.085 131.665 -63.755 131.995 ;
        RECT -64.085 129.655 -63.755 129.985 ;
        RECT -64.085 128.505 -63.755 128.835 ;
        RECT -64.085 126.495 -63.755 126.825 ;
        RECT -64.085 125.345 -63.755 125.675 ;
        RECT -64.085 123.335 -63.755 123.665 ;
        RECT -64.085 122.185 -63.755 122.515 ;
        RECT -64.085 120.175 -63.755 120.505 ;
        RECT -64.085 119.025 -63.755 119.355 ;
        RECT -64.085 117.185 -63.755 117.515 ;
        RECT -64.085 115.865 -63.755 116.195 ;
        RECT -64.085 113.855 -63.755 114.185 ;
        RECT -64.085 112.705 -63.755 113.035 ;
        RECT -64.085 110.695 -63.755 111.025 ;
        RECT -64.085 109.545 -63.755 109.875 ;
        RECT -64.085 107.535 -63.755 107.865 ;
        RECT -64.085 106.385 -63.755 106.715 ;
        RECT -64.085 104.375 -63.755 104.705 ;
        RECT -64.085 103.225 -63.755 103.555 ;
        RECT -64.085 100.865 -63.755 101.195 ;
        RECT -64.085 98.81 -63.755 99.14 ;
        RECT -64.085 97.755 -63.755 98.085 ;
        RECT -64.085 96.395 -63.755 96.725 ;
        RECT -64.085 95.035 -63.755 95.365 ;
        RECT -64.085 93.675 -63.755 94.005 ;
        RECT -64.085 92.315 -63.755 92.645 ;
        RECT -64.085 90.955 -63.755 91.285 ;
        RECT -64.085 89.595 -63.755 89.925 ;
        RECT -64.085 88.235 -63.755 88.565 ;
        RECT -64.085 86.875 -63.755 87.205 ;
        RECT -64.085 85.515 -63.755 85.845 ;
        RECT -64.085 84.155 -63.755 84.485 ;
        RECT -64.085 82.795 -63.755 83.125 ;
        RECT -64.085 81.435 -63.755 81.765 ;
        RECT -64.085 80.075 -63.755 80.405 ;
        RECT -64.085 78.715 -63.755 79.045 ;
        RECT -64.085 77.355 -63.755 77.685 ;
        RECT -64.085 75.995 -63.755 76.325 ;
        RECT -64.085 74.635 -63.755 74.965 ;
        RECT -64.085 73.275 -63.755 73.605 ;
        RECT -64.085 71.915 -63.755 72.245 ;
        RECT -64.085 70.555 -63.755 70.885 ;
        RECT -64.085 69.195 -63.755 69.525 ;
        RECT -64.085 67.835 -63.755 68.165 ;
        RECT -64.085 66.475 -63.755 66.805 ;
        RECT -64.085 65.115 -63.755 65.445 ;
        RECT -64.085 63.755 -63.755 64.085 ;
        RECT -64.085 62.395 -63.755 62.725 ;
        RECT -64.085 61.035 -63.755 61.365 ;
        RECT -64.085 59.675 -63.755 60.005 ;
        RECT -64.085 58.315 -63.755 58.645 ;
        RECT -64.085 56.955 -63.755 57.285 ;
        RECT -64.085 55.595 -63.755 55.925 ;
        RECT -64.085 54.235 -63.755 54.565 ;
        RECT -64.085 52.875 -63.755 53.205 ;
        RECT -64.085 51.515 -63.755 51.845 ;
        RECT -64.085 50.155 -63.755 50.485 ;
        RECT -64.085 48.795 -63.755 49.125 ;
        RECT -64.085 47.435 -63.755 47.765 ;
        RECT -64.085 46.075 -63.755 46.405 ;
        RECT -64.085 44.715 -63.755 45.045 ;
        RECT -64.085 43.355 -63.755 43.685 ;
        RECT -64.085 41.995 -63.755 42.325 ;
        RECT -64.085 40.635 -63.755 40.965 ;
        RECT -64.085 39.275 -63.755 39.605 ;
        RECT -64.085 37.915 -63.755 38.245 ;
        RECT -64.085 36.555 -63.755 36.885 ;
        RECT -64.085 35.195 -63.755 35.525 ;
        RECT -64.085 33.835 -63.755 34.165 ;
        RECT -64.085 32.475 -63.755 32.805 ;
        RECT -64.085 31.115 -63.755 31.445 ;
        RECT -64.085 29.755 -63.755 30.085 ;
        RECT -64.085 28.395 -63.755 28.725 ;
        RECT -64.085 27.035 -63.755 27.365 ;
        RECT -64.085 25.675 -63.755 26.005 ;
        RECT -64.085 24.315 -63.755 24.645 ;
        RECT -64.085 22.955 -63.755 23.285 ;
        RECT -64.085 21.595 -63.755 21.925 ;
        RECT -64.085 20.235 -63.755 20.565 ;
        RECT -64.085 18.875 -63.755 19.205 ;
        RECT -64.085 17.515 -63.755 17.845 ;
        RECT -64.085 16.155 -63.755 16.485 ;
        RECT -64.085 14.795 -63.755 15.125 ;
        RECT -64.085 13.435 -63.755 13.765 ;
        RECT -64.085 12.075 -63.755 12.405 ;
        RECT -64.085 10.715 -63.755 11.045 ;
        RECT -64.085 9.355 -63.755 9.685 ;
        RECT -64.085 7.995 -63.755 8.325 ;
        RECT -64.085 6.635 -63.755 6.965 ;
        RECT -64.085 5.275 -63.755 5.605 ;
        RECT -64.085 3.915 -63.755 4.245 ;
        RECT -64.085 2.555 -63.755 2.885 ;
        RECT -64.085 1.195 -63.755 1.525 ;
        RECT -64.085 -0.165 -63.755 0.165 ;
        RECT -64.085 -1.525 -63.755 -1.195 ;
        RECT -64.085 -2.885 -63.755 -2.555 ;
        RECT -64.085 -4.245 -63.755 -3.915 ;
        RECT -64.085 -5.605 -63.755 -5.275 ;
        RECT -64.085 -6.965 -63.755 -6.635 ;
        RECT -64.085 -8.325 -63.755 -7.995 ;
        RECT -64.085 -9.685 -63.755 -9.355 ;
        RECT -64.085 -11.045 -63.755 -10.715 ;
        RECT -64.085 -12.405 -63.755 -12.075 ;
        RECT -64.085 -13.765 -63.755 -13.435 ;
        RECT -64.085 -15.125 -63.755 -14.795 ;
        RECT -64.085 -16.485 -63.755 -16.155 ;
        RECT -64.085 -17.845 -63.755 -17.515 ;
        RECT -64.085 -19.205 -63.755 -18.875 ;
        RECT -64.085 -20.565 -63.755 -20.235 ;
        RECT -64.085 -21.925 -63.755 -21.595 ;
        RECT -64.085 -23.285 -63.755 -22.955 ;
        RECT -64.085 -24.645 -63.755 -24.315 ;
        RECT -64.085 -26.005 -63.755 -25.675 ;
        RECT -64.085 -27.365 -63.755 -27.035 ;
        RECT -64.085 -28.725 -63.755 -28.395 ;
        RECT -64.085 -30.085 -63.755 -29.755 ;
        RECT -64.085 -31.445 -63.755 -31.115 ;
        RECT -64.085 -32.805 -63.755 -32.475 ;
        RECT -64.085 -34.165 -63.755 -33.835 ;
        RECT -64.085 -35.525 -63.755 -35.195 ;
        RECT -64.085 -36.885 -63.755 -36.555 ;
        RECT -64.085 -38.245 -63.755 -37.915 ;
        RECT -64.085 -39.605 -63.755 -39.275 ;
        RECT -64.085 -40.965 -63.755 -40.635 ;
        RECT -64.085 -42.325 -63.755 -41.995 ;
        RECT -64.085 -43.685 -63.755 -43.355 ;
        RECT -64.085 -45.045 -63.755 -44.715 ;
        RECT -64.085 -46.405 -63.755 -46.075 ;
        RECT -64.085 -47.765 -63.755 -47.435 ;
        RECT -64.085 -49.125 -63.755 -48.795 ;
        RECT -64.085 -50.485 -63.755 -50.155 ;
        RECT -64.085 -51.845 -63.755 -51.515 ;
        RECT -64.085 -53.205 -63.755 -52.875 ;
        RECT -64.085 -54.565 -63.755 -54.235 ;
        RECT -64.085 -55.925 -63.755 -55.595 ;
        RECT -64.085 -57.285 -63.755 -56.955 ;
        RECT -64.085 -58.645 -63.755 -58.315 ;
        RECT -64.085 -60.005 -63.755 -59.675 ;
        RECT -64.085 -61.365 -63.755 -61.035 ;
        RECT -64.085 -62.725 -63.755 -62.395 ;
        RECT -64.085 -64.085 -63.755 -63.755 ;
        RECT -64.085 -65.445 -63.755 -65.115 ;
        RECT -64.085 -66.805 -63.755 -66.475 ;
        RECT -64.085 -68.165 -63.755 -67.835 ;
        RECT -64.085 -69.525 -63.755 -69.195 ;
        RECT -64.085 -70.885 -63.755 -70.555 ;
        RECT -64.085 -72.245 -63.755 -71.915 ;
        RECT -64.085 -73.605 -63.755 -73.275 ;
        RECT -64.085 -74.965 -63.755 -74.635 ;
        RECT -64.085 -76.325 -63.755 -75.995 ;
        RECT -64.085 -77.685 -63.755 -77.355 ;
        RECT -64.085 -79.045 -63.755 -78.715 ;
        RECT -64.085 -80.405 -63.755 -80.075 ;
        RECT -64.085 -81.765 -63.755 -81.435 ;
        RECT -64.085 -83.125 -63.755 -82.795 ;
        RECT -64.085 -84.485 -63.755 -84.155 ;
        RECT -64.085 -85.845 -63.755 -85.515 ;
        RECT -64.085 -87.205 -63.755 -86.875 ;
        RECT -64.085 -88.565 -63.755 -88.235 ;
        RECT -64.085 -89.925 -63.755 -89.595 ;
        RECT -64.085 -91.285 -63.755 -90.955 ;
        RECT -64.085 -92.645 -63.755 -92.315 ;
        RECT -64.085 -94.005 -63.755 -93.675 ;
        RECT -64.085 -95.365 -63.755 -95.035 ;
        RECT -64.085 -96.725 -63.755 -96.395 ;
        RECT -64.085 -98.085 -63.755 -97.755 ;
        RECT -64.085 -99.445 -63.755 -99.115 ;
        RECT -64.085 -100.805 -63.755 -100.475 ;
        RECT -64.085 -102.165 -63.755 -101.835 ;
        RECT -64.085 -103.525 -63.755 -103.195 ;
        RECT -64.085 -104.885 -63.755 -104.555 ;
        RECT -64.085 -106.245 -63.755 -105.915 ;
        RECT -64.085 -107.605 -63.755 -107.275 ;
        RECT -64.085 -108.965 -63.755 -108.635 ;
        RECT -64.085 -110.325 -63.755 -109.995 ;
        RECT -64.085 -111.685 -63.755 -111.355 ;
        RECT -64.085 -113.045 -63.755 -112.715 ;
        RECT -64.085 -114.405 -63.755 -114.075 ;
        RECT -64.085 -115.765 -63.755 -115.435 ;
        RECT -64.085 -117.125 -63.755 -116.795 ;
        RECT -64.085 -118.485 -63.755 -118.155 ;
        RECT -64.085 -119.845 -63.755 -119.515 ;
        RECT -64.085 -121.205 -63.755 -120.875 ;
        RECT -64.085 -122.565 -63.755 -122.235 ;
        RECT -64.085 -123.925 -63.755 -123.595 ;
        RECT -64.085 -125.285 -63.755 -124.955 ;
        RECT -64.085 -126.645 -63.755 -126.315 ;
        RECT -64.085 -128.005 -63.755 -127.675 ;
        RECT -64.085 -129.365 -63.755 -129.035 ;
        RECT -64.085 -130.725 -63.755 -130.395 ;
        RECT -64.085 -132.085 -63.755 -131.755 ;
        RECT -64.085 -133.445 -63.755 -133.115 ;
        RECT -64.085 -134.805 -63.755 -134.475 ;
        RECT -64.085 -136.165 -63.755 -135.835 ;
        RECT -64.085 -137.525 -63.755 -137.195 ;
        RECT -64.085 -138.885 -63.755 -138.555 ;
        RECT -64.085 -140.245 -63.755 -139.915 ;
        RECT -64.085 -141.605 -63.755 -141.275 ;
        RECT -64.085 -142.965 -63.755 -142.635 ;
        RECT -64.085 -144.325 -63.755 -143.995 ;
        RECT -64.085 -145.685 -63.755 -145.355 ;
        RECT -64.085 -147.045 -63.755 -146.715 ;
        RECT -64.085 -148.405 -63.755 -148.075 ;
        RECT -64.085 -149.765 -63.755 -149.435 ;
        RECT -64.085 -151.125 -63.755 -150.795 ;
        RECT -64.085 -152.485 -63.755 -152.155 ;
        RECT -64.085 -153.845 -63.755 -153.515 ;
        RECT -64.085 -155.205 -63.755 -154.875 ;
        RECT -64.085 -156.565 -63.755 -156.235 ;
        RECT -64.085 -157.925 -63.755 -157.595 ;
        RECT -64.085 -159.285 -63.755 -158.955 ;
        RECT -64.085 -160.645 -63.755 -160.315 ;
        RECT -64.085 -162.005 -63.755 -161.675 ;
        RECT -64.085 -163.365 -63.755 -163.035 ;
        RECT -64.085 -164.725 -63.755 -164.395 ;
        RECT -64.085 -166.085 -63.755 -165.755 ;
        RECT -64.085 -167.445 -63.755 -167.115 ;
        RECT -64.085 -170.165 -63.755 -169.835 ;
        RECT -64.085 -172.885 -63.755 -172.555 ;
        RECT -64.085 -174.245 -63.755 -173.915 ;
        RECT -64.085 -175.725 -63.755 -175.395 ;
        RECT -64.085 -176.965 -63.755 -176.635 ;
        RECT -64.085 -178.325 -63.755 -177.995 ;
        RECT -64.085 -180.57 -63.755 -179.44 ;
        RECT -64.08 -180.685 -63.76 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -62.725 241.32 -62.395 242.45 ;
        RECT -62.725 239.195 -62.395 239.525 ;
        RECT -62.725 237.835 -62.395 238.165 ;
        RECT -62.725 236.475 -62.395 236.805 ;
        RECT -62.725 235.115 -62.395 235.445 ;
        RECT -62.725 233.755 -62.395 234.085 ;
        RECT -62.725 232.395 -62.395 232.725 ;
        RECT -62.725 231.035 -62.395 231.365 ;
        RECT -62.725 229.675 -62.395 230.005 ;
        RECT -62.725 228.315 -62.395 228.645 ;
        RECT -62.725 226.955 -62.395 227.285 ;
        RECT -62.725 225.595 -62.395 225.925 ;
        RECT -62.725 224.235 -62.395 224.565 ;
        RECT -62.725 222.875 -62.395 223.205 ;
        RECT -62.725 221.515 -62.395 221.845 ;
        RECT -62.725 220.155 -62.395 220.485 ;
        RECT -62.725 218.795 -62.395 219.125 ;
        RECT -62.725 217.435 -62.395 217.765 ;
        RECT -62.725 216.075 -62.395 216.405 ;
        RECT -62.725 214.715 -62.395 215.045 ;
        RECT -62.725 213.355 -62.395 213.685 ;
        RECT -62.725 211.995 -62.395 212.325 ;
        RECT -62.725 210.635 -62.395 210.965 ;
        RECT -62.725 209.275 -62.395 209.605 ;
        RECT -62.725 207.915 -62.395 208.245 ;
        RECT -62.725 206.555 -62.395 206.885 ;
        RECT -62.725 205.195 -62.395 205.525 ;
        RECT -62.725 203.835 -62.395 204.165 ;
        RECT -62.725 202.475 -62.395 202.805 ;
        RECT -62.725 201.115 -62.395 201.445 ;
        RECT -62.725 199.755 -62.395 200.085 ;
        RECT -62.725 198.395 -62.395 198.725 ;
        RECT -62.725 197.035 -62.395 197.365 ;
        RECT -62.725 195.675 -62.395 196.005 ;
        RECT -62.725 194.315 -62.395 194.645 ;
        RECT -62.725 192.955 -62.395 193.285 ;
        RECT -62.725 191.595 -62.395 191.925 ;
        RECT -62.725 190.235 -62.395 190.565 ;
        RECT -62.725 188.875 -62.395 189.205 ;
        RECT -62.725 187.515 -62.395 187.845 ;
        RECT -62.725 186.155 -62.395 186.485 ;
        RECT -62.725 184.795 -62.395 185.125 ;
        RECT -62.725 183.435 -62.395 183.765 ;
        RECT -62.725 182.075 -62.395 182.405 ;
        RECT -62.725 180.715 -62.395 181.045 ;
        RECT -62.725 179.355 -62.395 179.685 ;
        RECT -62.725 177.995 -62.395 178.325 ;
        RECT -62.725 176.635 -62.395 176.965 ;
        RECT -62.725 175.275 -62.395 175.605 ;
        RECT -62.725 173.915 -62.395 174.245 ;
        RECT -62.725 172.555 -62.395 172.885 ;
        RECT -62.725 171.195 -62.395 171.525 ;
        RECT -62.725 169.835 -62.395 170.165 ;
        RECT -62.725 168.475 -62.395 168.805 ;
        RECT -62.725 167.115 -62.395 167.445 ;
        RECT -62.725 165.755 -62.395 166.085 ;
        RECT -62.725 164.395 -62.395 164.725 ;
        RECT -62.725 163.035 -62.395 163.365 ;
        RECT -62.725 161.675 -62.395 162.005 ;
        RECT -62.725 160.315 -62.395 160.645 ;
        RECT -62.725 158.955 -62.395 159.285 ;
        RECT -62.725 157.595 -62.395 157.925 ;
        RECT -62.725 156.235 -62.395 156.565 ;
        RECT -62.725 154.875 -62.395 155.205 ;
        RECT -62.725 153.515 -62.395 153.845 ;
        RECT -62.725 152.155 -62.395 152.485 ;
        RECT -62.725 150.795 -62.395 151.125 ;
        RECT -62.725 149.435 -62.395 149.765 ;
        RECT -62.725 148.075 -62.395 148.405 ;
        RECT -62.725 146.715 -62.395 147.045 ;
        RECT -62.725 145.355 -62.395 145.685 ;
        RECT -62.725 143.995 -62.395 144.325 ;
        RECT -62.725 142.635 -62.395 142.965 ;
        RECT -62.725 141.275 -62.395 141.605 ;
        RECT -62.725 139.915 -62.395 140.245 ;
        RECT -62.725 138.555 -62.395 138.885 ;
        RECT -62.725 137.225 -62.395 137.555 ;
        RECT -62.725 135.175 -62.395 135.505 ;
        RECT -62.725 132.815 -62.395 133.145 ;
        RECT -62.725 131.665 -62.395 131.995 ;
        RECT -62.725 129.655 -62.395 129.985 ;
        RECT -62.725 128.505 -62.395 128.835 ;
        RECT -62.725 126.495 -62.395 126.825 ;
        RECT -62.725 125.345 -62.395 125.675 ;
        RECT -62.725 123.335 -62.395 123.665 ;
        RECT -62.725 122.185 -62.395 122.515 ;
        RECT -62.725 120.175 -62.395 120.505 ;
        RECT -62.725 119.025 -62.395 119.355 ;
        RECT -62.725 117.185 -62.395 117.515 ;
        RECT -62.725 115.865 -62.395 116.195 ;
        RECT -62.725 113.855 -62.395 114.185 ;
        RECT -62.725 112.705 -62.395 113.035 ;
        RECT -62.725 110.695 -62.395 111.025 ;
        RECT -62.725 109.545 -62.395 109.875 ;
        RECT -62.725 107.535 -62.395 107.865 ;
        RECT -62.725 106.385 -62.395 106.715 ;
        RECT -62.725 104.375 -62.395 104.705 ;
        RECT -62.725 103.225 -62.395 103.555 ;
        RECT -62.725 100.865 -62.395 101.195 ;
        RECT -62.725 98.81 -62.395 99.14 ;
        RECT -62.725 97.755 -62.395 98.085 ;
        RECT -62.725 96.395 -62.395 96.725 ;
        RECT -62.725 95.035 -62.395 95.365 ;
        RECT -62.725 93.675 -62.395 94.005 ;
        RECT -62.725 92.315 -62.395 92.645 ;
        RECT -62.725 90.955 -62.395 91.285 ;
        RECT -62.725 89.595 -62.395 89.925 ;
        RECT -62.725 88.235 -62.395 88.565 ;
        RECT -62.725 86.875 -62.395 87.205 ;
        RECT -62.725 85.515 -62.395 85.845 ;
        RECT -62.725 84.155 -62.395 84.485 ;
        RECT -62.725 82.795 -62.395 83.125 ;
        RECT -62.725 81.435 -62.395 81.765 ;
        RECT -62.725 80.075 -62.395 80.405 ;
        RECT -62.725 78.715 -62.395 79.045 ;
        RECT -62.725 77.355 -62.395 77.685 ;
        RECT -62.725 75.995 -62.395 76.325 ;
        RECT -62.725 74.635 -62.395 74.965 ;
        RECT -62.725 73.275 -62.395 73.605 ;
        RECT -62.725 71.915 -62.395 72.245 ;
        RECT -62.725 70.555 -62.395 70.885 ;
        RECT -62.725 69.195 -62.395 69.525 ;
        RECT -62.725 67.835 -62.395 68.165 ;
        RECT -62.725 66.475 -62.395 66.805 ;
        RECT -62.725 65.115 -62.395 65.445 ;
        RECT -62.725 63.755 -62.395 64.085 ;
        RECT -62.725 62.395 -62.395 62.725 ;
        RECT -62.725 61.035 -62.395 61.365 ;
        RECT -62.725 59.675 -62.395 60.005 ;
        RECT -62.725 58.315 -62.395 58.645 ;
        RECT -62.725 56.955 -62.395 57.285 ;
        RECT -62.725 55.595 -62.395 55.925 ;
        RECT -62.725 54.235 -62.395 54.565 ;
        RECT -62.725 52.875 -62.395 53.205 ;
        RECT -62.725 51.515 -62.395 51.845 ;
        RECT -62.725 50.155 -62.395 50.485 ;
        RECT -62.725 48.795 -62.395 49.125 ;
        RECT -62.725 47.435 -62.395 47.765 ;
        RECT -62.725 46.075 -62.395 46.405 ;
        RECT -62.725 44.715 -62.395 45.045 ;
        RECT -62.725 43.355 -62.395 43.685 ;
        RECT -62.725 41.995 -62.395 42.325 ;
        RECT -62.725 40.635 -62.395 40.965 ;
        RECT -62.725 39.275 -62.395 39.605 ;
        RECT -62.725 37.915 -62.395 38.245 ;
        RECT -62.725 36.555 -62.395 36.885 ;
        RECT -62.725 35.195 -62.395 35.525 ;
        RECT -62.725 33.835 -62.395 34.165 ;
        RECT -62.725 32.475 -62.395 32.805 ;
        RECT -62.725 31.115 -62.395 31.445 ;
        RECT -62.725 29.755 -62.395 30.085 ;
        RECT -62.725 28.395 -62.395 28.725 ;
        RECT -62.725 27.035 -62.395 27.365 ;
        RECT -62.725 25.675 -62.395 26.005 ;
        RECT -62.725 24.315 -62.395 24.645 ;
        RECT -62.725 22.955 -62.395 23.285 ;
        RECT -62.725 21.595 -62.395 21.925 ;
        RECT -62.725 20.235 -62.395 20.565 ;
        RECT -62.725 18.875 -62.395 19.205 ;
        RECT -62.725 17.515 -62.395 17.845 ;
        RECT -62.725 16.155 -62.395 16.485 ;
        RECT -62.725 14.795 -62.395 15.125 ;
        RECT -62.725 13.435 -62.395 13.765 ;
        RECT -62.725 12.075 -62.395 12.405 ;
        RECT -62.725 10.715 -62.395 11.045 ;
        RECT -62.725 9.355 -62.395 9.685 ;
        RECT -62.725 7.995 -62.395 8.325 ;
        RECT -62.725 6.635 -62.395 6.965 ;
        RECT -62.725 5.275 -62.395 5.605 ;
        RECT -62.725 3.915 -62.395 4.245 ;
        RECT -62.725 2.555 -62.395 2.885 ;
        RECT -62.725 1.195 -62.395 1.525 ;
        RECT -62.725 -0.165 -62.395 0.165 ;
        RECT -62.725 -1.525 -62.395 -1.195 ;
        RECT -62.725 -2.885 -62.395 -2.555 ;
        RECT -62.725 -4.245 -62.395 -3.915 ;
        RECT -62.725 -5.605 -62.395 -5.275 ;
        RECT -62.725 -6.965 -62.395 -6.635 ;
        RECT -62.725 -8.325 -62.395 -7.995 ;
        RECT -62.725 -9.685 -62.395 -9.355 ;
        RECT -62.725 -11.045 -62.395 -10.715 ;
        RECT -62.725 -12.405 -62.395 -12.075 ;
        RECT -62.725 -13.765 -62.395 -13.435 ;
        RECT -62.725 -15.125 -62.395 -14.795 ;
        RECT -62.725 -16.485 -62.395 -16.155 ;
        RECT -62.725 -17.845 -62.395 -17.515 ;
        RECT -62.725 -19.205 -62.395 -18.875 ;
        RECT -62.725 -20.565 -62.395 -20.235 ;
        RECT -62.725 -21.925 -62.395 -21.595 ;
        RECT -62.725 -23.285 -62.395 -22.955 ;
        RECT -62.725 -24.645 -62.395 -24.315 ;
        RECT -62.725 -26.005 -62.395 -25.675 ;
        RECT -62.725 -27.365 -62.395 -27.035 ;
        RECT -62.725 -28.725 -62.395 -28.395 ;
        RECT -62.725 -30.085 -62.395 -29.755 ;
        RECT -62.725 -31.445 -62.395 -31.115 ;
        RECT -62.725 -32.805 -62.395 -32.475 ;
        RECT -62.725 -34.165 -62.395 -33.835 ;
        RECT -62.725 -35.525 -62.395 -35.195 ;
        RECT -62.725 -36.885 -62.395 -36.555 ;
        RECT -62.725 -38.245 -62.395 -37.915 ;
        RECT -62.725 -39.605 -62.395 -39.275 ;
        RECT -62.725 -40.965 -62.395 -40.635 ;
        RECT -62.725 -42.325 -62.395 -41.995 ;
        RECT -62.725 -43.685 -62.395 -43.355 ;
        RECT -62.725 -45.045 -62.395 -44.715 ;
        RECT -62.725 -46.405 -62.395 -46.075 ;
        RECT -62.725 -47.765 -62.395 -47.435 ;
        RECT -62.725 -49.125 -62.395 -48.795 ;
        RECT -62.725 -50.485 -62.395 -50.155 ;
        RECT -62.725 -51.845 -62.395 -51.515 ;
        RECT -62.725 -53.205 -62.395 -52.875 ;
        RECT -62.725 -54.565 -62.395 -54.235 ;
        RECT -62.725 -55.925 -62.395 -55.595 ;
        RECT -62.725 -57.285 -62.395 -56.955 ;
        RECT -62.725 -58.645 -62.395 -58.315 ;
        RECT -62.725 -60.005 -62.395 -59.675 ;
        RECT -62.725 -61.365 -62.395 -61.035 ;
        RECT -62.725 -62.725 -62.395 -62.395 ;
        RECT -62.725 -64.085 -62.395 -63.755 ;
        RECT -62.725 -65.445 -62.395 -65.115 ;
        RECT -62.725 -66.805 -62.395 -66.475 ;
        RECT -62.725 -68.165 -62.395 -67.835 ;
        RECT -62.725 -69.525 -62.395 -69.195 ;
        RECT -62.725 -70.885 -62.395 -70.555 ;
        RECT -62.725 -72.245 -62.395 -71.915 ;
        RECT -62.725 -73.605 -62.395 -73.275 ;
        RECT -62.725 -74.965 -62.395 -74.635 ;
        RECT -62.725 -76.325 -62.395 -75.995 ;
        RECT -62.725 -77.685 -62.395 -77.355 ;
        RECT -62.725 -79.045 -62.395 -78.715 ;
        RECT -62.725 -80.405 -62.395 -80.075 ;
        RECT -62.725 -81.765 -62.395 -81.435 ;
        RECT -62.725 -83.125 -62.395 -82.795 ;
        RECT -62.725 -84.485 -62.395 -84.155 ;
        RECT -62.725 -85.845 -62.395 -85.515 ;
        RECT -62.725 -87.205 -62.395 -86.875 ;
        RECT -62.725 -88.565 -62.395 -88.235 ;
        RECT -62.725 -89.925 -62.395 -89.595 ;
        RECT -62.725 -91.285 -62.395 -90.955 ;
        RECT -62.725 -92.645 -62.395 -92.315 ;
        RECT -62.725 -94.005 -62.395 -93.675 ;
        RECT -62.725 -95.365 -62.395 -95.035 ;
        RECT -62.725 -96.725 -62.395 -96.395 ;
        RECT -62.725 -98.085 -62.395 -97.755 ;
        RECT -62.725 -99.445 -62.395 -99.115 ;
        RECT -62.725 -100.805 -62.395 -100.475 ;
        RECT -62.725 -102.165 -62.395 -101.835 ;
        RECT -62.725 -103.525 -62.395 -103.195 ;
        RECT -62.725 -104.885 -62.395 -104.555 ;
        RECT -62.725 -106.245 -62.395 -105.915 ;
        RECT -62.725 -107.605 -62.395 -107.275 ;
        RECT -62.725 -108.965 -62.395 -108.635 ;
        RECT -62.725 -110.325 -62.395 -109.995 ;
        RECT -62.725 -111.685 -62.395 -111.355 ;
        RECT -62.725 -113.045 -62.395 -112.715 ;
        RECT -62.725 -114.405 -62.395 -114.075 ;
        RECT -62.725 -115.765 -62.395 -115.435 ;
        RECT -62.725 -117.125 -62.395 -116.795 ;
        RECT -62.725 -118.485 -62.395 -118.155 ;
        RECT -62.725 -119.845 -62.395 -119.515 ;
        RECT -62.725 -121.205 -62.395 -120.875 ;
        RECT -62.725 -122.565 -62.395 -122.235 ;
        RECT -62.725 -123.925 -62.395 -123.595 ;
        RECT -62.725 -125.285 -62.395 -124.955 ;
        RECT -62.725 -126.645 -62.395 -126.315 ;
        RECT -62.725 -128.005 -62.395 -127.675 ;
        RECT -62.725 -129.365 -62.395 -129.035 ;
        RECT -62.725 -130.725 -62.395 -130.395 ;
        RECT -62.725 -132.085 -62.395 -131.755 ;
        RECT -62.725 -133.445 -62.395 -133.115 ;
        RECT -62.725 -134.805 -62.395 -134.475 ;
        RECT -62.725 -136.165 -62.395 -135.835 ;
        RECT -62.725 -137.525 -62.395 -137.195 ;
        RECT -62.725 -138.885 -62.395 -138.555 ;
        RECT -62.725 -140.245 -62.395 -139.915 ;
        RECT -62.725 -141.605 -62.395 -141.275 ;
        RECT -62.725 -142.965 -62.395 -142.635 ;
        RECT -62.725 -144.325 -62.395 -143.995 ;
        RECT -62.725 -145.685 -62.395 -145.355 ;
        RECT -62.725 -147.045 -62.395 -146.715 ;
        RECT -62.725 -148.405 -62.395 -148.075 ;
        RECT -62.725 -149.765 -62.395 -149.435 ;
        RECT -62.725 -151.125 -62.395 -150.795 ;
        RECT -62.725 -152.485 -62.395 -152.155 ;
        RECT -62.725 -153.845 -62.395 -153.515 ;
        RECT -62.725 -155.205 -62.395 -154.875 ;
        RECT -62.725 -156.565 -62.395 -156.235 ;
        RECT -62.725 -157.925 -62.395 -157.595 ;
        RECT -62.725 -159.285 -62.395 -158.955 ;
        RECT -62.725 -160.645 -62.395 -160.315 ;
        RECT -62.725 -162.005 -62.395 -161.675 ;
        RECT -62.725 -163.365 -62.395 -163.035 ;
        RECT -62.725 -164.725 -62.395 -164.395 ;
        RECT -62.725 -166.085 -62.395 -165.755 ;
        RECT -62.725 -167.445 -62.395 -167.115 ;
        RECT -62.725 -170.165 -62.395 -169.835 ;
        RECT -62.725 -172.885 -62.395 -172.555 ;
        RECT -62.725 -174.245 -62.395 -173.915 ;
        RECT -62.725 -175.725 -62.395 -175.395 ;
        RECT -62.725 -176.965 -62.395 -176.635 ;
        RECT -62.725 -178.325 -62.395 -177.995 ;
        RECT -62.725 -180.57 -62.395 -179.44 ;
        RECT -62.72 -180.685 -62.4 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -61.365 191.595 -61.035 191.925 ;
        RECT -61.365 190.235 -61.035 190.565 ;
        RECT -61.365 188.875 -61.035 189.205 ;
        RECT -61.365 187.515 -61.035 187.845 ;
        RECT -61.365 186.155 -61.035 186.485 ;
        RECT -61.365 184.795 -61.035 185.125 ;
        RECT -61.365 183.435 -61.035 183.765 ;
        RECT -61.365 182.075 -61.035 182.405 ;
        RECT -61.365 180.715 -61.035 181.045 ;
        RECT -61.365 179.355 -61.035 179.685 ;
        RECT -61.365 177.995 -61.035 178.325 ;
        RECT -61.365 176.635 -61.035 176.965 ;
        RECT -61.365 175.275 -61.035 175.605 ;
        RECT -61.365 173.915 -61.035 174.245 ;
        RECT -61.365 172.555 -61.035 172.885 ;
        RECT -61.365 171.195 -61.035 171.525 ;
        RECT -61.365 169.835 -61.035 170.165 ;
        RECT -61.365 168.475 -61.035 168.805 ;
        RECT -61.365 167.115 -61.035 167.445 ;
        RECT -61.365 165.755 -61.035 166.085 ;
        RECT -61.365 164.395 -61.035 164.725 ;
        RECT -61.365 163.035 -61.035 163.365 ;
        RECT -61.365 161.675 -61.035 162.005 ;
        RECT -61.365 160.315 -61.035 160.645 ;
        RECT -61.365 158.955 -61.035 159.285 ;
        RECT -61.365 157.595 -61.035 157.925 ;
        RECT -61.365 156.235 -61.035 156.565 ;
        RECT -61.365 154.875 -61.035 155.205 ;
        RECT -61.365 153.515 -61.035 153.845 ;
        RECT -61.365 152.155 -61.035 152.485 ;
        RECT -61.365 150.795 -61.035 151.125 ;
        RECT -61.365 149.435 -61.035 149.765 ;
        RECT -61.365 148.075 -61.035 148.405 ;
        RECT -61.365 146.715 -61.035 147.045 ;
        RECT -61.365 145.355 -61.035 145.685 ;
        RECT -61.365 143.995 -61.035 144.325 ;
        RECT -61.365 142.635 -61.035 142.965 ;
        RECT -61.365 141.275 -61.035 141.605 ;
        RECT -61.365 139.915 -61.035 140.245 ;
        RECT -61.365 138.555 -61.035 138.885 ;
        RECT -61.365 137.225 -61.035 137.555 ;
        RECT -61.365 135.175 -61.035 135.505 ;
        RECT -61.365 132.815 -61.035 133.145 ;
        RECT -61.365 131.665 -61.035 131.995 ;
        RECT -61.365 129.655 -61.035 129.985 ;
        RECT -61.365 128.505 -61.035 128.835 ;
        RECT -61.365 126.495 -61.035 126.825 ;
        RECT -61.365 125.345 -61.035 125.675 ;
        RECT -61.365 123.335 -61.035 123.665 ;
        RECT -61.365 122.185 -61.035 122.515 ;
        RECT -61.365 120.175 -61.035 120.505 ;
        RECT -61.365 119.025 -61.035 119.355 ;
        RECT -61.365 117.185 -61.035 117.515 ;
        RECT -61.365 115.865 -61.035 116.195 ;
        RECT -61.365 113.855 -61.035 114.185 ;
        RECT -61.365 112.705 -61.035 113.035 ;
        RECT -61.365 110.695 -61.035 111.025 ;
        RECT -61.365 109.545 -61.035 109.875 ;
        RECT -61.365 107.535 -61.035 107.865 ;
        RECT -61.365 106.385 -61.035 106.715 ;
        RECT -61.365 104.375 -61.035 104.705 ;
        RECT -61.365 103.225 -61.035 103.555 ;
        RECT -61.365 100.865 -61.035 101.195 ;
        RECT -61.365 98.81 -61.035 99.14 ;
        RECT -61.365 97.755 -61.035 98.085 ;
        RECT -61.365 96.395 -61.035 96.725 ;
        RECT -61.365 95.035 -61.035 95.365 ;
        RECT -61.365 93.675 -61.035 94.005 ;
        RECT -61.365 92.315 -61.035 92.645 ;
        RECT -61.365 90.955 -61.035 91.285 ;
        RECT -61.365 89.595 -61.035 89.925 ;
        RECT -61.365 88.235 -61.035 88.565 ;
        RECT -61.365 86.875 -61.035 87.205 ;
        RECT -61.365 85.515 -61.035 85.845 ;
        RECT -61.365 84.155 -61.035 84.485 ;
        RECT -61.365 82.795 -61.035 83.125 ;
        RECT -61.365 81.435 -61.035 81.765 ;
        RECT -61.365 80.075 -61.035 80.405 ;
        RECT -61.365 78.715 -61.035 79.045 ;
        RECT -61.365 77.355 -61.035 77.685 ;
        RECT -61.365 75.995 -61.035 76.325 ;
        RECT -61.365 74.635 -61.035 74.965 ;
        RECT -61.365 73.275 -61.035 73.605 ;
        RECT -61.365 71.915 -61.035 72.245 ;
        RECT -61.365 70.555 -61.035 70.885 ;
        RECT -61.365 69.195 -61.035 69.525 ;
        RECT -61.365 67.835 -61.035 68.165 ;
        RECT -61.365 66.475 -61.035 66.805 ;
        RECT -61.365 65.115 -61.035 65.445 ;
        RECT -61.365 63.755 -61.035 64.085 ;
        RECT -61.365 62.395 -61.035 62.725 ;
        RECT -61.365 61.035 -61.035 61.365 ;
        RECT -61.365 59.675 -61.035 60.005 ;
        RECT -61.365 58.315 -61.035 58.645 ;
        RECT -61.365 56.955 -61.035 57.285 ;
        RECT -61.365 55.595 -61.035 55.925 ;
        RECT -61.365 54.235 -61.035 54.565 ;
        RECT -61.365 52.875 -61.035 53.205 ;
        RECT -61.365 51.515 -61.035 51.845 ;
        RECT -61.365 50.155 -61.035 50.485 ;
        RECT -61.365 48.795 -61.035 49.125 ;
        RECT -61.365 47.435 -61.035 47.765 ;
        RECT -61.365 46.075 -61.035 46.405 ;
        RECT -61.365 44.715 -61.035 45.045 ;
        RECT -61.365 43.355 -61.035 43.685 ;
        RECT -61.365 41.995 -61.035 42.325 ;
        RECT -61.365 40.635 -61.035 40.965 ;
        RECT -61.365 39.275 -61.035 39.605 ;
        RECT -61.365 37.915 -61.035 38.245 ;
        RECT -61.365 36.555 -61.035 36.885 ;
        RECT -61.365 35.195 -61.035 35.525 ;
        RECT -61.365 33.835 -61.035 34.165 ;
        RECT -61.365 32.475 -61.035 32.805 ;
        RECT -61.365 31.115 -61.035 31.445 ;
        RECT -61.365 29.755 -61.035 30.085 ;
        RECT -61.365 28.395 -61.035 28.725 ;
        RECT -61.365 27.035 -61.035 27.365 ;
        RECT -61.365 25.675 -61.035 26.005 ;
        RECT -61.365 24.315 -61.035 24.645 ;
        RECT -61.365 22.955 -61.035 23.285 ;
        RECT -61.365 21.595 -61.035 21.925 ;
        RECT -61.365 20.235 -61.035 20.565 ;
        RECT -61.365 18.875 -61.035 19.205 ;
        RECT -61.365 17.515 -61.035 17.845 ;
        RECT -61.365 16.155 -61.035 16.485 ;
        RECT -61.365 14.795 -61.035 15.125 ;
        RECT -61.365 13.435 -61.035 13.765 ;
        RECT -61.365 12.075 -61.035 12.405 ;
        RECT -61.365 10.715 -61.035 11.045 ;
        RECT -61.365 9.355 -61.035 9.685 ;
        RECT -61.365 7.995 -61.035 8.325 ;
        RECT -61.365 6.635 -61.035 6.965 ;
        RECT -61.365 5.275 -61.035 5.605 ;
        RECT -61.365 3.915 -61.035 4.245 ;
        RECT -61.365 2.555 -61.035 2.885 ;
        RECT -61.365 1.195 -61.035 1.525 ;
        RECT -61.365 -0.165 -61.035 0.165 ;
        RECT -61.365 -1.525 -61.035 -1.195 ;
        RECT -61.365 -2.885 -61.035 -2.555 ;
        RECT -61.365 -4.245 -61.035 -3.915 ;
        RECT -61.365 -5.605 -61.035 -5.275 ;
        RECT -61.365 -6.965 -61.035 -6.635 ;
        RECT -61.365 -8.325 -61.035 -7.995 ;
        RECT -61.365 -9.685 -61.035 -9.355 ;
        RECT -61.365 -11.045 -61.035 -10.715 ;
        RECT -61.365 -12.405 -61.035 -12.075 ;
        RECT -61.365 -13.765 -61.035 -13.435 ;
        RECT -61.365 -15.125 -61.035 -14.795 ;
        RECT -61.365 -16.485 -61.035 -16.155 ;
        RECT -61.365 -17.845 -61.035 -17.515 ;
        RECT -61.365 -19.205 -61.035 -18.875 ;
        RECT -61.365 -20.565 -61.035 -20.235 ;
        RECT -61.365 -21.925 -61.035 -21.595 ;
        RECT -61.365 -23.285 -61.035 -22.955 ;
        RECT -61.365 -24.645 -61.035 -24.315 ;
        RECT -61.365 -26.005 -61.035 -25.675 ;
        RECT -61.365 -27.365 -61.035 -27.035 ;
        RECT -61.365 -28.725 -61.035 -28.395 ;
        RECT -61.365 -30.085 -61.035 -29.755 ;
        RECT -61.365 -31.445 -61.035 -31.115 ;
        RECT -61.365 -32.805 -61.035 -32.475 ;
        RECT -61.365 -34.165 -61.035 -33.835 ;
        RECT -61.365 -35.525 -61.035 -35.195 ;
        RECT -61.365 -36.885 -61.035 -36.555 ;
        RECT -61.365 -38.245 -61.035 -37.915 ;
        RECT -61.365 -39.605 -61.035 -39.275 ;
        RECT -61.365 -40.965 -61.035 -40.635 ;
        RECT -61.365 -42.325 -61.035 -41.995 ;
        RECT -61.365 -43.685 -61.035 -43.355 ;
        RECT -61.365 -45.045 -61.035 -44.715 ;
        RECT -61.365 -46.405 -61.035 -46.075 ;
        RECT -61.365 -47.765 -61.035 -47.435 ;
        RECT -61.365 -49.125 -61.035 -48.795 ;
        RECT -61.365 -50.485 -61.035 -50.155 ;
        RECT -61.365 -51.845 -61.035 -51.515 ;
        RECT -61.365 -53.205 -61.035 -52.875 ;
        RECT -61.365 -54.565 -61.035 -54.235 ;
        RECT -61.365 -55.925 -61.035 -55.595 ;
        RECT -61.365 -57.285 -61.035 -56.955 ;
        RECT -61.365 -58.645 -61.035 -58.315 ;
        RECT -61.365 -60.005 -61.035 -59.675 ;
        RECT -61.365 -61.365 -61.035 -61.035 ;
        RECT -61.365 -62.725 -61.035 -62.395 ;
        RECT -61.365 -64.085 -61.035 -63.755 ;
        RECT -61.365 -65.445 -61.035 -65.115 ;
        RECT -61.365 -66.805 -61.035 -66.475 ;
        RECT -61.365 -68.165 -61.035 -67.835 ;
        RECT -61.365 -69.525 -61.035 -69.195 ;
        RECT -61.365 -70.885 -61.035 -70.555 ;
        RECT -61.365 -72.245 -61.035 -71.915 ;
        RECT -61.365 -73.605 -61.035 -73.275 ;
        RECT -61.365 -74.965 -61.035 -74.635 ;
        RECT -61.365 -76.325 -61.035 -75.995 ;
        RECT -61.365 -77.685 -61.035 -77.355 ;
        RECT -61.365 -79.045 -61.035 -78.715 ;
        RECT -61.365 -80.405 -61.035 -80.075 ;
        RECT -61.365 -81.765 -61.035 -81.435 ;
        RECT -61.365 -83.125 -61.035 -82.795 ;
        RECT -61.365 -84.485 -61.035 -84.155 ;
        RECT -61.365 -85.845 -61.035 -85.515 ;
        RECT -61.365 -87.205 -61.035 -86.875 ;
        RECT -61.365 -88.565 -61.035 -88.235 ;
        RECT -61.365 -89.925 -61.035 -89.595 ;
        RECT -61.365 -92.645 -61.035 -92.315 ;
        RECT -61.365 -94.005 -61.035 -93.675 ;
        RECT -61.365 -95.365 -61.035 -95.035 ;
        RECT -61.365 -96.725 -61.035 -96.395 ;
        RECT -61.365 -99.445 -61.035 -99.115 ;
        RECT -61.365 -102.165 -61.035 -101.835 ;
        RECT -61.365 -103.525 -61.035 -103.195 ;
        RECT -61.365 -104.885 -61.035 -104.555 ;
        RECT -61.365 -107.605 -61.035 -107.275 ;
        RECT -61.365 -108.965 -61.035 -108.635 ;
        RECT -61.365 -110.325 -61.035 -109.995 ;
        RECT -61.36 -112.36 -61.04 242.565 ;
        RECT -61.365 241.32 -61.035 242.45 ;
        RECT -61.365 239.195 -61.035 239.525 ;
        RECT -61.365 237.835 -61.035 238.165 ;
        RECT -61.365 236.475 -61.035 236.805 ;
        RECT -61.365 235.115 -61.035 235.445 ;
        RECT -61.365 233.755 -61.035 234.085 ;
        RECT -61.365 232.395 -61.035 232.725 ;
        RECT -61.365 231.035 -61.035 231.365 ;
        RECT -61.365 229.675 -61.035 230.005 ;
        RECT -61.365 228.315 -61.035 228.645 ;
        RECT -61.365 226.955 -61.035 227.285 ;
        RECT -61.365 225.595 -61.035 225.925 ;
        RECT -61.365 224.235 -61.035 224.565 ;
        RECT -61.365 222.875 -61.035 223.205 ;
        RECT -61.365 221.515 -61.035 221.845 ;
        RECT -61.365 220.155 -61.035 220.485 ;
        RECT -61.365 218.795 -61.035 219.125 ;
        RECT -61.365 217.435 -61.035 217.765 ;
        RECT -61.365 216.075 -61.035 216.405 ;
        RECT -61.365 214.715 -61.035 215.045 ;
        RECT -61.365 213.355 -61.035 213.685 ;
        RECT -61.365 211.995 -61.035 212.325 ;
        RECT -61.365 210.635 -61.035 210.965 ;
        RECT -61.365 209.275 -61.035 209.605 ;
        RECT -61.365 207.915 -61.035 208.245 ;
        RECT -61.365 206.555 -61.035 206.885 ;
        RECT -61.365 205.195 -61.035 205.525 ;
        RECT -61.365 203.835 -61.035 204.165 ;
        RECT -61.365 202.475 -61.035 202.805 ;
        RECT -61.365 201.115 -61.035 201.445 ;
        RECT -61.365 199.755 -61.035 200.085 ;
        RECT -61.365 198.395 -61.035 198.725 ;
        RECT -61.365 197.035 -61.035 197.365 ;
        RECT -61.365 195.675 -61.035 196.005 ;
        RECT -61.365 194.315 -61.035 194.645 ;
        RECT -61.365 192.955 -61.035 193.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -68.165 241.32 -67.835 242.45 ;
        RECT -68.165 239.195 -67.835 239.525 ;
        RECT -68.165 237.835 -67.835 238.165 ;
        RECT -68.165 236.475 -67.835 236.805 ;
        RECT -68.165 235.115 -67.835 235.445 ;
        RECT -68.165 233.755 -67.835 234.085 ;
        RECT -68.165 232.395 -67.835 232.725 ;
        RECT -68.165 231.035 -67.835 231.365 ;
        RECT -68.165 229.675 -67.835 230.005 ;
        RECT -68.165 228.315 -67.835 228.645 ;
        RECT -68.165 226.955 -67.835 227.285 ;
        RECT -68.165 225.595 -67.835 225.925 ;
        RECT -68.165 224.235 -67.835 224.565 ;
        RECT -68.165 222.875 -67.835 223.205 ;
        RECT -68.165 221.515 -67.835 221.845 ;
        RECT -68.165 220.155 -67.835 220.485 ;
        RECT -68.165 218.795 -67.835 219.125 ;
        RECT -68.165 217.435 -67.835 217.765 ;
        RECT -68.165 216.075 -67.835 216.405 ;
        RECT -68.165 214.715 -67.835 215.045 ;
        RECT -68.165 213.355 -67.835 213.685 ;
        RECT -68.165 211.995 -67.835 212.325 ;
        RECT -68.165 210.635 -67.835 210.965 ;
        RECT -68.165 209.275 -67.835 209.605 ;
        RECT -68.165 207.915 -67.835 208.245 ;
        RECT -68.165 206.555 -67.835 206.885 ;
        RECT -68.165 205.195 -67.835 205.525 ;
        RECT -68.165 203.835 -67.835 204.165 ;
        RECT -68.165 202.475 -67.835 202.805 ;
        RECT -68.165 201.115 -67.835 201.445 ;
        RECT -68.165 199.755 -67.835 200.085 ;
        RECT -68.165 198.395 -67.835 198.725 ;
        RECT -68.165 197.035 -67.835 197.365 ;
        RECT -68.165 195.675 -67.835 196.005 ;
        RECT -68.165 194.315 -67.835 194.645 ;
        RECT -68.165 192.955 -67.835 193.285 ;
        RECT -68.165 191.595 -67.835 191.925 ;
        RECT -68.165 190.235 -67.835 190.565 ;
        RECT -68.165 188.875 -67.835 189.205 ;
        RECT -68.165 187.515 -67.835 187.845 ;
        RECT -68.165 186.155 -67.835 186.485 ;
        RECT -68.165 184.795 -67.835 185.125 ;
        RECT -68.165 183.435 -67.835 183.765 ;
        RECT -68.165 182.075 -67.835 182.405 ;
        RECT -68.165 180.715 -67.835 181.045 ;
        RECT -68.165 179.355 -67.835 179.685 ;
        RECT -68.165 177.995 -67.835 178.325 ;
        RECT -68.165 176.635 -67.835 176.965 ;
        RECT -68.165 175.275 -67.835 175.605 ;
        RECT -68.165 173.915 -67.835 174.245 ;
        RECT -68.165 172.555 -67.835 172.885 ;
        RECT -68.165 171.195 -67.835 171.525 ;
        RECT -68.165 169.835 -67.835 170.165 ;
        RECT -68.165 168.475 -67.835 168.805 ;
        RECT -68.165 167.115 -67.835 167.445 ;
        RECT -68.165 165.755 -67.835 166.085 ;
        RECT -68.165 164.395 -67.835 164.725 ;
        RECT -68.165 163.035 -67.835 163.365 ;
        RECT -68.165 161.675 -67.835 162.005 ;
        RECT -68.165 160.315 -67.835 160.645 ;
        RECT -68.165 158.955 -67.835 159.285 ;
        RECT -68.165 157.595 -67.835 157.925 ;
        RECT -68.165 156.235 -67.835 156.565 ;
        RECT -68.165 154.875 -67.835 155.205 ;
        RECT -68.165 153.515 -67.835 153.845 ;
        RECT -68.165 152.155 -67.835 152.485 ;
        RECT -68.165 150.795 -67.835 151.125 ;
        RECT -68.165 149.435 -67.835 149.765 ;
        RECT -68.165 148.075 -67.835 148.405 ;
        RECT -68.165 146.715 -67.835 147.045 ;
        RECT -68.165 145.355 -67.835 145.685 ;
        RECT -68.165 143.995 -67.835 144.325 ;
        RECT -68.165 142.635 -67.835 142.965 ;
        RECT -68.165 141.275 -67.835 141.605 ;
        RECT -68.165 139.915 -67.835 140.245 ;
        RECT -68.165 138.555 -67.835 138.885 ;
        RECT -68.165 137.195 -67.835 137.525 ;
        RECT -68.165 135.835 -67.835 136.165 ;
        RECT -68.165 134.475 -67.835 134.805 ;
        RECT -68.165 133.115 -67.835 133.445 ;
        RECT -68.165 131.755 -67.835 132.085 ;
        RECT -68.165 130.395 -67.835 130.725 ;
        RECT -68.165 129.035 -67.835 129.365 ;
        RECT -68.165 127.675 -67.835 128.005 ;
        RECT -68.165 126.315 -67.835 126.645 ;
        RECT -68.165 124.955 -67.835 125.285 ;
        RECT -68.165 123.595 -67.835 123.925 ;
        RECT -68.165 122.235 -67.835 122.565 ;
        RECT -68.165 120.875 -67.835 121.205 ;
        RECT -68.165 119.515 -67.835 119.845 ;
        RECT -68.165 118.155 -67.835 118.485 ;
        RECT -68.165 116.795 -67.835 117.125 ;
        RECT -68.165 115.435 -67.835 115.765 ;
        RECT -68.165 114.075 -67.835 114.405 ;
        RECT -68.165 112.715 -67.835 113.045 ;
        RECT -68.165 111.355 -67.835 111.685 ;
        RECT -68.165 109.995 -67.835 110.325 ;
        RECT -68.165 108.635 -67.835 108.965 ;
        RECT -68.165 107.275 -67.835 107.605 ;
        RECT -68.165 105.915 -67.835 106.245 ;
        RECT -68.165 104.555 -67.835 104.885 ;
        RECT -68.165 103.195 -67.835 103.525 ;
        RECT -68.165 101.835 -67.835 102.165 ;
        RECT -68.165 100.475 -67.835 100.805 ;
        RECT -68.165 99.115 -67.835 99.445 ;
        RECT -68.165 97.755 -67.835 98.085 ;
        RECT -68.165 96.395 -67.835 96.725 ;
        RECT -68.165 95.035 -67.835 95.365 ;
        RECT -68.165 93.675 -67.835 94.005 ;
        RECT -68.165 92.315 -67.835 92.645 ;
        RECT -68.165 90.955 -67.835 91.285 ;
        RECT -68.165 89.595 -67.835 89.925 ;
        RECT -68.165 88.235 -67.835 88.565 ;
        RECT -68.165 86.875 -67.835 87.205 ;
        RECT -68.165 85.515 -67.835 85.845 ;
        RECT -68.165 84.155 -67.835 84.485 ;
        RECT -68.165 82.795 -67.835 83.125 ;
        RECT -68.165 81.435 -67.835 81.765 ;
        RECT -68.165 80.075 -67.835 80.405 ;
        RECT -68.165 78.715 -67.835 79.045 ;
        RECT -68.165 77.355 -67.835 77.685 ;
        RECT -68.165 75.995 -67.835 76.325 ;
        RECT -68.165 74.635 -67.835 74.965 ;
        RECT -68.165 73.275 -67.835 73.605 ;
        RECT -68.165 71.915 -67.835 72.245 ;
        RECT -68.165 70.555 -67.835 70.885 ;
        RECT -68.165 69.195 -67.835 69.525 ;
        RECT -68.165 67.835 -67.835 68.165 ;
        RECT -68.165 66.475 -67.835 66.805 ;
        RECT -68.165 65.115 -67.835 65.445 ;
        RECT -68.165 63.755 -67.835 64.085 ;
        RECT -68.165 62.395 -67.835 62.725 ;
        RECT -68.165 61.035 -67.835 61.365 ;
        RECT -68.165 59.675 -67.835 60.005 ;
        RECT -68.165 58.315 -67.835 58.645 ;
        RECT -68.165 56.955 -67.835 57.285 ;
        RECT -68.165 55.595 -67.835 55.925 ;
        RECT -68.165 54.235 -67.835 54.565 ;
        RECT -68.165 52.875 -67.835 53.205 ;
        RECT -68.165 51.515 -67.835 51.845 ;
        RECT -68.165 50.155 -67.835 50.485 ;
        RECT -68.165 48.795 -67.835 49.125 ;
        RECT -68.165 47.435 -67.835 47.765 ;
        RECT -68.165 46.075 -67.835 46.405 ;
        RECT -68.165 44.715 -67.835 45.045 ;
        RECT -68.165 43.355 -67.835 43.685 ;
        RECT -68.165 41.995 -67.835 42.325 ;
        RECT -68.165 40.635 -67.835 40.965 ;
        RECT -68.165 39.275 -67.835 39.605 ;
        RECT -68.165 37.915 -67.835 38.245 ;
        RECT -68.165 36.555 -67.835 36.885 ;
        RECT -68.165 35.195 -67.835 35.525 ;
        RECT -68.165 33.835 -67.835 34.165 ;
        RECT -68.165 32.475 -67.835 32.805 ;
        RECT -68.165 31.115 -67.835 31.445 ;
        RECT -68.165 29.755 -67.835 30.085 ;
        RECT -68.165 28.395 -67.835 28.725 ;
        RECT -68.165 27.035 -67.835 27.365 ;
        RECT -68.165 25.675 -67.835 26.005 ;
        RECT -68.165 24.315 -67.835 24.645 ;
        RECT -68.165 22.955 -67.835 23.285 ;
        RECT -68.165 21.595 -67.835 21.925 ;
        RECT -68.165 20.235 -67.835 20.565 ;
        RECT -68.165 18.875 -67.835 19.205 ;
        RECT -68.165 17.515 -67.835 17.845 ;
        RECT -68.165 16.155 -67.835 16.485 ;
        RECT -68.165 14.795 -67.835 15.125 ;
        RECT -68.165 13.435 -67.835 13.765 ;
        RECT -68.165 12.075 -67.835 12.405 ;
        RECT -68.165 10.715 -67.835 11.045 ;
        RECT -68.165 9.355 -67.835 9.685 ;
        RECT -68.165 7.995 -67.835 8.325 ;
        RECT -68.165 6.635 -67.835 6.965 ;
        RECT -68.165 5.275 -67.835 5.605 ;
        RECT -68.165 3.915 -67.835 4.245 ;
        RECT -68.165 2.555 -67.835 2.885 ;
        RECT -68.165 1.195 -67.835 1.525 ;
        RECT -68.165 -0.165 -67.835 0.165 ;
        RECT -68.165 -1.525 -67.835 -1.195 ;
        RECT -68.165 -2.885 -67.835 -2.555 ;
        RECT -68.165 -4.245 -67.835 -3.915 ;
        RECT -68.165 -5.605 -67.835 -5.275 ;
        RECT -68.165 -6.965 -67.835 -6.635 ;
        RECT -68.165 -8.325 -67.835 -7.995 ;
        RECT -68.165 -9.685 -67.835 -9.355 ;
        RECT -68.165 -11.045 -67.835 -10.715 ;
        RECT -68.165 -12.405 -67.835 -12.075 ;
        RECT -68.165 -13.765 -67.835 -13.435 ;
        RECT -68.165 -15.125 -67.835 -14.795 ;
        RECT -68.165 -16.485 -67.835 -16.155 ;
        RECT -68.165 -17.845 -67.835 -17.515 ;
        RECT -68.165 -19.205 -67.835 -18.875 ;
        RECT -68.165 -20.565 -67.835 -20.235 ;
        RECT -68.165 -21.925 -67.835 -21.595 ;
        RECT -68.165 -23.285 -67.835 -22.955 ;
        RECT -68.165 -24.645 -67.835 -24.315 ;
        RECT -68.165 -26.005 -67.835 -25.675 ;
        RECT -68.165 -27.365 -67.835 -27.035 ;
        RECT -68.165 -28.725 -67.835 -28.395 ;
        RECT -68.165 -30.085 -67.835 -29.755 ;
        RECT -68.165 -31.445 -67.835 -31.115 ;
        RECT -68.165 -32.805 -67.835 -32.475 ;
        RECT -68.165 -34.165 -67.835 -33.835 ;
        RECT -68.165 -35.525 -67.835 -35.195 ;
        RECT -68.165 -36.885 -67.835 -36.555 ;
        RECT -68.165 -38.245 -67.835 -37.915 ;
        RECT -68.165 -39.605 -67.835 -39.275 ;
        RECT -68.165 -40.965 -67.835 -40.635 ;
        RECT -68.165 -42.325 -67.835 -41.995 ;
        RECT -68.165 -43.685 -67.835 -43.355 ;
        RECT -68.165 -45.045 -67.835 -44.715 ;
        RECT -68.165 -46.405 -67.835 -46.075 ;
        RECT -68.165 -47.765 -67.835 -47.435 ;
        RECT -68.165 -49.125 -67.835 -48.795 ;
        RECT -68.165 -50.485 -67.835 -50.155 ;
        RECT -68.165 -51.845 -67.835 -51.515 ;
        RECT -68.165 -53.205 -67.835 -52.875 ;
        RECT -68.165 -54.565 -67.835 -54.235 ;
        RECT -68.165 -55.925 -67.835 -55.595 ;
        RECT -68.165 -57.285 -67.835 -56.955 ;
        RECT -68.165 -58.645 -67.835 -58.315 ;
        RECT -68.165 -60.005 -67.835 -59.675 ;
        RECT -68.165 -61.365 -67.835 -61.035 ;
        RECT -68.165 -62.725 -67.835 -62.395 ;
        RECT -68.165 -64.085 -67.835 -63.755 ;
        RECT -68.165 -65.445 -67.835 -65.115 ;
        RECT -68.165 -66.805 -67.835 -66.475 ;
        RECT -68.165 -68.165 -67.835 -67.835 ;
        RECT -68.165 -69.525 -67.835 -69.195 ;
        RECT -68.165 -70.885 -67.835 -70.555 ;
        RECT -68.165 -72.245 -67.835 -71.915 ;
        RECT -68.165 -73.605 -67.835 -73.275 ;
        RECT -68.165 -74.965 -67.835 -74.635 ;
        RECT -68.165 -76.325 -67.835 -75.995 ;
        RECT -68.165 -77.685 -67.835 -77.355 ;
        RECT -68.165 -79.045 -67.835 -78.715 ;
        RECT -68.165 -80.405 -67.835 -80.075 ;
        RECT -68.165 -81.765 -67.835 -81.435 ;
        RECT -68.165 -83.125 -67.835 -82.795 ;
        RECT -68.165 -84.485 -67.835 -84.155 ;
        RECT -68.165 -85.845 -67.835 -85.515 ;
        RECT -68.165 -87.205 -67.835 -86.875 ;
        RECT -68.165 -88.565 -67.835 -88.235 ;
        RECT -68.165 -89.925 -67.835 -89.595 ;
        RECT -68.165 -91.285 -67.835 -90.955 ;
        RECT -68.165 -92.645 -67.835 -92.315 ;
        RECT -68.165 -94.005 -67.835 -93.675 ;
        RECT -68.165 -95.365 -67.835 -95.035 ;
        RECT -68.165 -96.725 -67.835 -96.395 ;
        RECT -68.165 -98.085 -67.835 -97.755 ;
        RECT -68.165 -99.445 -67.835 -99.115 ;
        RECT -68.165 -100.805 -67.835 -100.475 ;
        RECT -68.165 -102.165 -67.835 -101.835 ;
        RECT -68.165 -103.525 -67.835 -103.195 ;
        RECT -68.165 -104.885 -67.835 -104.555 ;
        RECT -68.165 -106.245 -67.835 -105.915 ;
        RECT -68.165 -107.605 -67.835 -107.275 ;
        RECT -68.165 -108.965 -67.835 -108.635 ;
        RECT -68.165 -110.325 -67.835 -109.995 ;
        RECT -68.165 -111.685 -67.835 -111.355 ;
        RECT -68.165 -113.045 -67.835 -112.715 ;
        RECT -68.165 -114.405 -67.835 -114.075 ;
        RECT -68.165 -115.765 -67.835 -115.435 ;
        RECT -68.165 -117.125 -67.835 -116.795 ;
        RECT -68.165 -118.485 -67.835 -118.155 ;
        RECT -68.165 -119.845 -67.835 -119.515 ;
        RECT -68.165 -121.205 -67.835 -120.875 ;
        RECT -68.165 -122.565 -67.835 -122.235 ;
        RECT -68.165 -123.925 -67.835 -123.595 ;
        RECT -68.165 -125.285 -67.835 -124.955 ;
        RECT -68.165 -126.645 -67.835 -126.315 ;
        RECT -68.165 -128.005 -67.835 -127.675 ;
        RECT -68.165 -129.365 -67.835 -129.035 ;
        RECT -68.165 -130.725 -67.835 -130.395 ;
        RECT -68.165 -132.085 -67.835 -131.755 ;
        RECT -68.165 -133.445 -67.835 -133.115 ;
        RECT -68.165 -134.805 -67.835 -134.475 ;
        RECT -68.165 -136.165 -67.835 -135.835 ;
        RECT -68.165 -137.525 -67.835 -137.195 ;
        RECT -68.165 -138.885 -67.835 -138.555 ;
        RECT -68.165 -140.245 -67.835 -139.915 ;
        RECT -68.165 -141.605 -67.835 -141.275 ;
        RECT -68.165 -142.965 -67.835 -142.635 ;
        RECT -68.165 -144.325 -67.835 -143.995 ;
        RECT -68.165 -145.685 -67.835 -145.355 ;
        RECT -68.165 -147.045 -67.835 -146.715 ;
        RECT -68.165 -148.405 -67.835 -148.075 ;
        RECT -68.165 -149.765 -67.835 -149.435 ;
        RECT -68.165 -151.125 -67.835 -150.795 ;
        RECT -68.165 -152.485 -67.835 -152.155 ;
        RECT -68.165 -153.845 -67.835 -153.515 ;
        RECT -68.165 -155.205 -67.835 -154.875 ;
        RECT -68.165 -156.565 -67.835 -156.235 ;
        RECT -68.165 -157.925 -67.835 -157.595 ;
        RECT -68.165 -159.285 -67.835 -158.955 ;
        RECT -68.165 -160.645 -67.835 -160.315 ;
        RECT -68.165 -162.005 -67.835 -161.675 ;
        RECT -68.165 -163.365 -67.835 -163.035 ;
        RECT -68.165 -164.725 -67.835 -164.395 ;
        RECT -68.165 -166.085 -67.835 -165.755 ;
        RECT -68.165 -167.445 -67.835 -167.115 ;
        RECT -68.165 -170.165 -67.835 -169.835 ;
        RECT -68.165 -172.885 -67.835 -172.555 ;
        RECT -68.165 -174.245 -67.835 -173.915 ;
        RECT -68.165 -175.725 -67.835 -175.395 ;
        RECT -68.165 -176.965 -67.835 -176.635 ;
        RECT -68.165 -178.325 -67.835 -177.995 ;
        RECT -68.165 -180.57 -67.835 -179.44 ;
        RECT -68.16 -180.685 -67.84 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -66.805 241.32 -66.475 242.45 ;
        RECT -66.805 239.195 -66.475 239.525 ;
        RECT -66.805 237.835 -66.475 238.165 ;
        RECT -66.805 236.475 -66.475 236.805 ;
        RECT -66.805 235.115 -66.475 235.445 ;
        RECT -66.805 233.755 -66.475 234.085 ;
        RECT -66.805 232.395 -66.475 232.725 ;
        RECT -66.805 231.035 -66.475 231.365 ;
        RECT -66.805 229.675 -66.475 230.005 ;
        RECT -66.805 228.315 -66.475 228.645 ;
        RECT -66.805 226.955 -66.475 227.285 ;
        RECT -66.805 225.595 -66.475 225.925 ;
        RECT -66.805 224.235 -66.475 224.565 ;
        RECT -66.805 222.875 -66.475 223.205 ;
        RECT -66.805 221.515 -66.475 221.845 ;
        RECT -66.805 220.155 -66.475 220.485 ;
        RECT -66.805 218.795 -66.475 219.125 ;
        RECT -66.805 217.435 -66.475 217.765 ;
        RECT -66.805 216.075 -66.475 216.405 ;
        RECT -66.805 214.715 -66.475 215.045 ;
        RECT -66.805 213.355 -66.475 213.685 ;
        RECT -66.805 211.995 -66.475 212.325 ;
        RECT -66.805 210.635 -66.475 210.965 ;
        RECT -66.805 209.275 -66.475 209.605 ;
        RECT -66.805 207.915 -66.475 208.245 ;
        RECT -66.805 206.555 -66.475 206.885 ;
        RECT -66.805 205.195 -66.475 205.525 ;
        RECT -66.805 203.835 -66.475 204.165 ;
        RECT -66.805 202.475 -66.475 202.805 ;
        RECT -66.805 201.115 -66.475 201.445 ;
        RECT -66.805 199.755 -66.475 200.085 ;
        RECT -66.805 198.395 -66.475 198.725 ;
        RECT -66.805 197.035 -66.475 197.365 ;
        RECT -66.805 195.675 -66.475 196.005 ;
        RECT -66.805 194.315 -66.475 194.645 ;
        RECT -66.805 192.955 -66.475 193.285 ;
        RECT -66.805 191.595 -66.475 191.925 ;
        RECT -66.805 190.235 -66.475 190.565 ;
        RECT -66.805 188.875 -66.475 189.205 ;
        RECT -66.805 187.515 -66.475 187.845 ;
        RECT -66.805 186.155 -66.475 186.485 ;
        RECT -66.805 184.795 -66.475 185.125 ;
        RECT -66.805 183.435 -66.475 183.765 ;
        RECT -66.805 182.075 -66.475 182.405 ;
        RECT -66.805 180.715 -66.475 181.045 ;
        RECT -66.805 179.355 -66.475 179.685 ;
        RECT -66.805 177.995 -66.475 178.325 ;
        RECT -66.805 176.635 -66.475 176.965 ;
        RECT -66.805 175.275 -66.475 175.605 ;
        RECT -66.805 173.915 -66.475 174.245 ;
        RECT -66.805 172.555 -66.475 172.885 ;
        RECT -66.805 171.195 -66.475 171.525 ;
        RECT -66.805 169.835 -66.475 170.165 ;
        RECT -66.805 168.475 -66.475 168.805 ;
        RECT -66.805 167.115 -66.475 167.445 ;
        RECT -66.805 165.755 -66.475 166.085 ;
        RECT -66.805 164.395 -66.475 164.725 ;
        RECT -66.805 163.035 -66.475 163.365 ;
        RECT -66.805 161.675 -66.475 162.005 ;
        RECT -66.805 160.315 -66.475 160.645 ;
        RECT -66.805 158.955 -66.475 159.285 ;
        RECT -66.805 157.595 -66.475 157.925 ;
        RECT -66.805 156.235 -66.475 156.565 ;
        RECT -66.805 154.875 -66.475 155.205 ;
        RECT -66.805 153.515 -66.475 153.845 ;
        RECT -66.805 152.155 -66.475 152.485 ;
        RECT -66.805 150.795 -66.475 151.125 ;
        RECT -66.805 149.435 -66.475 149.765 ;
        RECT -66.805 148.075 -66.475 148.405 ;
        RECT -66.805 146.715 -66.475 147.045 ;
        RECT -66.805 145.355 -66.475 145.685 ;
        RECT -66.805 143.995 -66.475 144.325 ;
        RECT -66.805 142.635 -66.475 142.965 ;
        RECT -66.805 141.275 -66.475 141.605 ;
        RECT -66.805 139.915 -66.475 140.245 ;
        RECT -66.805 138.555 -66.475 138.885 ;
        RECT -66.805 137.195 -66.475 137.525 ;
        RECT -66.805 135.835 -66.475 136.165 ;
        RECT -66.805 134.475 -66.475 134.805 ;
        RECT -66.805 133.115 -66.475 133.445 ;
        RECT -66.805 131.755 -66.475 132.085 ;
        RECT -66.805 130.395 -66.475 130.725 ;
        RECT -66.805 129.035 -66.475 129.365 ;
        RECT -66.805 127.675 -66.475 128.005 ;
        RECT -66.805 126.315 -66.475 126.645 ;
        RECT -66.805 124.955 -66.475 125.285 ;
        RECT -66.805 123.595 -66.475 123.925 ;
        RECT -66.805 122.235 -66.475 122.565 ;
        RECT -66.805 120.875 -66.475 121.205 ;
        RECT -66.805 119.515 -66.475 119.845 ;
        RECT -66.805 118.155 -66.475 118.485 ;
        RECT -66.805 116.795 -66.475 117.125 ;
        RECT -66.805 115.435 -66.475 115.765 ;
        RECT -66.805 114.075 -66.475 114.405 ;
        RECT -66.805 112.715 -66.475 113.045 ;
        RECT -66.805 111.355 -66.475 111.685 ;
        RECT -66.805 109.995 -66.475 110.325 ;
        RECT -66.805 108.635 -66.475 108.965 ;
        RECT -66.805 107.275 -66.475 107.605 ;
        RECT -66.805 105.915 -66.475 106.245 ;
        RECT -66.805 104.555 -66.475 104.885 ;
        RECT -66.805 103.195 -66.475 103.525 ;
        RECT -66.805 101.835 -66.475 102.165 ;
        RECT -66.805 100.475 -66.475 100.805 ;
        RECT -66.805 99.115 -66.475 99.445 ;
        RECT -66.805 97.755 -66.475 98.085 ;
        RECT -66.805 96.395 -66.475 96.725 ;
        RECT -66.805 95.035 -66.475 95.365 ;
        RECT -66.805 93.675 -66.475 94.005 ;
        RECT -66.805 92.315 -66.475 92.645 ;
        RECT -66.805 90.955 -66.475 91.285 ;
        RECT -66.805 89.595 -66.475 89.925 ;
        RECT -66.805 88.235 -66.475 88.565 ;
        RECT -66.805 86.875 -66.475 87.205 ;
        RECT -66.805 85.515 -66.475 85.845 ;
        RECT -66.805 84.155 -66.475 84.485 ;
        RECT -66.805 82.795 -66.475 83.125 ;
        RECT -66.805 81.435 -66.475 81.765 ;
        RECT -66.805 80.075 -66.475 80.405 ;
        RECT -66.805 78.715 -66.475 79.045 ;
        RECT -66.805 77.355 -66.475 77.685 ;
        RECT -66.805 75.995 -66.475 76.325 ;
        RECT -66.805 74.635 -66.475 74.965 ;
        RECT -66.805 73.275 -66.475 73.605 ;
        RECT -66.805 71.915 -66.475 72.245 ;
        RECT -66.805 70.555 -66.475 70.885 ;
        RECT -66.805 69.195 -66.475 69.525 ;
        RECT -66.805 67.835 -66.475 68.165 ;
        RECT -66.805 66.475 -66.475 66.805 ;
        RECT -66.805 65.115 -66.475 65.445 ;
        RECT -66.805 63.755 -66.475 64.085 ;
        RECT -66.805 62.395 -66.475 62.725 ;
        RECT -66.805 61.035 -66.475 61.365 ;
        RECT -66.805 59.675 -66.475 60.005 ;
        RECT -66.805 58.315 -66.475 58.645 ;
        RECT -66.805 56.955 -66.475 57.285 ;
        RECT -66.805 55.595 -66.475 55.925 ;
        RECT -66.805 54.235 -66.475 54.565 ;
        RECT -66.805 52.875 -66.475 53.205 ;
        RECT -66.805 51.515 -66.475 51.845 ;
        RECT -66.805 50.155 -66.475 50.485 ;
        RECT -66.805 48.795 -66.475 49.125 ;
        RECT -66.805 47.435 -66.475 47.765 ;
        RECT -66.805 46.075 -66.475 46.405 ;
        RECT -66.805 44.715 -66.475 45.045 ;
        RECT -66.805 43.355 -66.475 43.685 ;
        RECT -66.805 41.995 -66.475 42.325 ;
        RECT -66.805 40.635 -66.475 40.965 ;
        RECT -66.805 39.275 -66.475 39.605 ;
        RECT -66.805 37.915 -66.475 38.245 ;
        RECT -66.805 36.555 -66.475 36.885 ;
        RECT -66.805 35.195 -66.475 35.525 ;
        RECT -66.805 33.835 -66.475 34.165 ;
        RECT -66.805 32.475 -66.475 32.805 ;
        RECT -66.805 31.115 -66.475 31.445 ;
        RECT -66.805 29.755 -66.475 30.085 ;
        RECT -66.805 28.395 -66.475 28.725 ;
        RECT -66.805 27.035 -66.475 27.365 ;
        RECT -66.805 25.675 -66.475 26.005 ;
        RECT -66.805 24.315 -66.475 24.645 ;
        RECT -66.805 22.955 -66.475 23.285 ;
        RECT -66.805 21.595 -66.475 21.925 ;
        RECT -66.805 20.235 -66.475 20.565 ;
        RECT -66.805 18.875 -66.475 19.205 ;
        RECT -66.805 17.515 -66.475 17.845 ;
        RECT -66.805 16.155 -66.475 16.485 ;
        RECT -66.805 14.795 -66.475 15.125 ;
        RECT -66.805 13.435 -66.475 13.765 ;
        RECT -66.805 12.075 -66.475 12.405 ;
        RECT -66.805 10.715 -66.475 11.045 ;
        RECT -66.805 9.355 -66.475 9.685 ;
        RECT -66.805 7.995 -66.475 8.325 ;
        RECT -66.805 6.635 -66.475 6.965 ;
        RECT -66.805 5.275 -66.475 5.605 ;
        RECT -66.805 3.915 -66.475 4.245 ;
        RECT -66.805 2.555 -66.475 2.885 ;
        RECT -66.805 1.195 -66.475 1.525 ;
        RECT -66.805 -0.165 -66.475 0.165 ;
        RECT -66.805 -1.525 -66.475 -1.195 ;
        RECT -66.805 -2.885 -66.475 -2.555 ;
        RECT -66.805 -4.245 -66.475 -3.915 ;
        RECT -66.805 -5.605 -66.475 -5.275 ;
        RECT -66.805 -6.965 -66.475 -6.635 ;
        RECT -66.805 -8.325 -66.475 -7.995 ;
        RECT -66.805 -9.685 -66.475 -9.355 ;
        RECT -66.805 -11.045 -66.475 -10.715 ;
        RECT -66.805 -12.405 -66.475 -12.075 ;
        RECT -66.805 -13.765 -66.475 -13.435 ;
        RECT -66.805 -15.125 -66.475 -14.795 ;
        RECT -66.805 -16.485 -66.475 -16.155 ;
        RECT -66.805 -17.845 -66.475 -17.515 ;
        RECT -66.805 -19.205 -66.475 -18.875 ;
        RECT -66.805 -20.565 -66.475 -20.235 ;
        RECT -66.805 -21.925 -66.475 -21.595 ;
        RECT -66.805 -23.285 -66.475 -22.955 ;
        RECT -66.805 -24.645 -66.475 -24.315 ;
        RECT -66.805 -26.005 -66.475 -25.675 ;
        RECT -66.805 -27.365 -66.475 -27.035 ;
        RECT -66.805 -28.725 -66.475 -28.395 ;
        RECT -66.805 -30.085 -66.475 -29.755 ;
        RECT -66.805 -31.445 -66.475 -31.115 ;
        RECT -66.805 -32.805 -66.475 -32.475 ;
        RECT -66.805 -34.165 -66.475 -33.835 ;
        RECT -66.805 -35.525 -66.475 -35.195 ;
        RECT -66.805 -36.885 -66.475 -36.555 ;
        RECT -66.805 -38.245 -66.475 -37.915 ;
        RECT -66.805 -39.605 -66.475 -39.275 ;
        RECT -66.805 -40.965 -66.475 -40.635 ;
        RECT -66.805 -42.325 -66.475 -41.995 ;
        RECT -66.805 -43.685 -66.475 -43.355 ;
        RECT -66.805 -45.045 -66.475 -44.715 ;
        RECT -66.805 -46.405 -66.475 -46.075 ;
        RECT -66.805 -47.765 -66.475 -47.435 ;
        RECT -66.805 -49.125 -66.475 -48.795 ;
        RECT -66.805 -50.485 -66.475 -50.155 ;
        RECT -66.805 -51.845 -66.475 -51.515 ;
        RECT -66.805 -53.205 -66.475 -52.875 ;
        RECT -66.805 -54.565 -66.475 -54.235 ;
        RECT -66.805 -55.925 -66.475 -55.595 ;
        RECT -66.805 -57.285 -66.475 -56.955 ;
        RECT -66.805 -58.645 -66.475 -58.315 ;
        RECT -66.805 -60.005 -66.475 -59.675 ;
        RECT -66.805 -61.365 -66.475 -61.035 ;
        RECT -66.805 -62.725 -66.475 -62.395 ;
        RECT -66.805 -64.085 -66.475 -63.755 ;
        RECT -66.805 -65.445 -66.475 -65.115 ;
        RECT -66.805 -66.805 -66.475 -66.475 ;
        RECT -66.805 -68.165 -66.475 -67.835 ;
        RECT -66.805 -69.525 -66.475 -69.195 ;
        RECT -66.805 -70.885 -66.475 -70.555 ;
        RECT -66.805 -72.245 -66.475 -71.915 ;
        RECT -66.805 -73.605 -66.475 -73.275 ;
        RECT -66.805 -74.965 -66.475 -74.635 ;
        RECT -66.805 -76.325 -66.475 -75.995 ;
        RECT -66.805 -77.685 -66.475 -77.355 ;
        RECT -66.805 -79.045 -66.475 -78.715 ;
        RECT -66.805 -80.405 -66.475 -80.075 ;
        RECT -66.805 -81.765 -66.475 -81.435 ;
        RECT -66.805 -83.125 -66.475 -82.795 ;
        RECT -66.805 -84.485 -66.475 -84.155 ;
        RECT -66.805 -85.845 -66.475 -85.515 ;
        RECT -66.805 -87.205 -66.475 -86.875 ;
        RECT -66.805 -88.565 -66.475 -88.235 ;
        RECT -66.805 -89.925 -66.475 -89.595 ;
        RECT -66.805 -91.285 -66.475 -90.955 ;
        RECT -66.805 -92.645 -66.475 -92.315 ;
        RECT -66.805 -94.005 -66.475 -93.675 ;
        RECT -66.805 -95.365 -66.475 -95.035 ;
        RECT -66.805 -96.725 -66.475 -96.395 ;
        RECT -66.805 -98.085 -66.475 -97.755 ;
        RECT -66.805 -99.445 -66.475 -99.115 ;
        RECT -66.805 -100.805 -66.475 -100.475 ;
        RECT -66.805 -102.165 -66.475 -101.835 ;
        RECT -66.805 -103.525 -66.475 -103.195 ;
        RECT -66.805 -104.885 -66.475 -104.555 ;
        RECT -66.805 -106.245 -66.475 -105.915 ;
        RECT -66.805 -107.605 -66.475 -107.275 ;
        RECT -66.805 -108.965 -66.475 -108.635 ;
        RECT -66.805 -110.325 -66.475 -109.995 ;
        RECT -66.805 -111.685 -66.475 -111.355 ;
        RECT -66.805 -113.045 -66.475 -112.715 ;
        RECT -66.805 -114.405 -66.475 -114.075 ;
        RECT -66.805 -115.765 -66.475 -115.435 ;
        RECT -66.805 -117.125 -66.475 -116.795 ;
        RECT -66.805 -118.485 -66.475 -118.155 ;
        RECT -66.805 -119.845 -66.475 -119.515 ;
        RECT -66.805 -121.205 -66.475 -120.875 ;
        RECT -66.805 -122.565 -66.475 -122.235 ;
        RECT -66.805 -123.925 -66.475 -123.595 ;
        RECT -66.805 -125.285 -66.475 -124.955 ;
        RECT -66.805 -126.645 -66.475 -126.315 ;
        RECT -66.805 -128.005 -66.475 -127.675 ;
        RECT -66.805 -129.365 -66.475 -129.035 ;
        RECT -66.805 -130.725 -66.475 -130.395 ;
        RECT -66.805 -132.085 -66.475 -131.755 ;
        RECT -66.805 -133.445 -66.475 -133.115 ;
        RECT -66.805 -134.805 -66.475 -134.475 ;
        RECT -66.805 -136.165 -66.475 -135.835 ;
        RECT -66.805 -137.525 -66.475 -137.195 ;
        RECT -66.805 -138.885 -66.475 -138.555 ;
        RECT -66.805 -140.245 -66.475 -139.915 ;
        RECT -66.805 -141.605 -66.475 -141.275 ;
        RECT -66.805 -142.965 -66.475 -142.635 ;
        RECT -66.805 -144.325 -66.475 -143.995 ;
        RECT -66.805 -145.685 -66.475 -145.355 ;
        RECT -66.805 -147.045 -66.475 -146.715 ;
        RECT -66.805 -148.405 -66.475 -148.075 ;
        RECT -66.805 -149.765 -66.475 -149.435 ;
        RECT -66.805 -151.125 -66.475 -150.795 ;
        RECT -66.805 -152.485 -66.475 -152.155 ;
        RECT -66.805 -153.845 -66.475 -153.515 ;
        RECT -66.805 -155.205 -66.475 -154.875 ;
        RECT -66.805 -156.565 -66.475 -156.235 ;
        RECT -66.805 -157.925 -66.475 -157.595 ;
        RECT -66.805 -159.285 -66.475 -158.955 ;
        RECT -66.805 -160.645 -66.475 -160.315 ;
        RECT -66.805 -162.005 -66.475 -161.675 ;
        RECT -66.805 -163.365 -66.475 -163.035 ;
        RECT -66.805 -164.725 -66.475 -164.395 ;
        RECT -66.805 -166.085 -66.475 -165.755 ;
        RECT -66.805 -167.445 -66.475 -167.115 ;
        RECT -66.805 -170.165 -66.475 -169.835 ;
        RECT -66.805 -174.245 -66.475 -173.915 ;
        RECT -66.805 -175.725 -66.475 -175.395 ;
        RECT -66.805 -176.965 -66.475 -176.635 ;
        RECT -66.805 -178.325 -66.475 -177.995 ;
        RECT -66.805 -180.57 -66.475 -179.44 ;
        RECT -66.8 -180.685 -66.48 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -65.445 -0.165 -65.115 0.165 ;
        RECT -65.445 -1.525 -65.115 -1.195 ;
        RECT -65.445 -2.885 -65.115 -2.555 ;
        RECT -65.445 -4.245 -65.115 -3.915 ;
        RECT -65.445 -5.605 -65.115 -5.275 ;
        RECT -65.445 -6.965 -65.115 -6.635 ;
        RECT -65.445 -8.325 -65.115 -7.995 ;
        RECT -65.445 -9.685 -65.115 -9.355 ;
        RECT -65.445 -11.045 -65.115 -10.715 ;
        RECT -65.445 -12.405 -65.115 -12.075 ;
        RECT -65.445 -13.765 -65.115 -13.435 ;
        RECT -65.445 -15.125 -65.115 -14.795 ;
        RECT -65.445 -16.485 -65.115 -16.155 ;
        RECT -65.445 -17.845 -65.115 -17.515 ;
        RECT -65.445 -19.205 -65.115 -18.875 ;
        RECT -65.445 -20.565 -65.115 -20.235 ;
        RECT -65.445 -21.925 -65.115 -21.595 ;
        RECT -65.445 -23.285 -65.115 -22.955 ;
        RECT -65.445 -24.645 -65.115 -24.315 ;
        RECT -65.445 -26.005 -65.115 -25.675 ;
        RECT -65.445 -27.365 -65.115 -27.035 ;
        RECT -65.445 -28.725 -65.115 -28.395 ;
        RECT -65.445 -30.085 -65.115 -29.755 ;
        RECT -65.445 -31.445 -65.115 -31.115 ;
        RECT -65.445 -32.805 -65.115 -32.475 ;
        RECT -65.445 -34.165 -65.115 -33.835 ;
        RECT -65.445 -35.525 -65.115 -35.195 ;
        RECT -65.445 -36.885 -65.115 -36.555 ;
        RECT -65.445 -38.245 -65.115 -37.915 ;
        RECT -65.445 -39.605 -65.115 -39.275 ;
        RECT -65.445 -40.965 -65.115 -40.635 ;
        RECT -65.445 -42.325 -65.115 -41.995 ;
        RECT -65.445 -43.685 -65.115 -43.355 ;
        RECT -65.445 -45.045 -65.115 -44.715 ;
        RECT -65.445 -46.405 -65.115 -46.075 ;
        RECT -65.445 -47.765 -65.115 -47.435 ;
        RECT -65.445 -49.125 -65.115 -48.795 ;
        RECT -65.445 -50.485 -65.115 -50.155 ;
        RECT -65.445 -51.845 -65.115 -51.515 ;
        RECT -65.445 -53.205 -65.115 -52.875 ;
        RECT -65.445 -54.565 -65.115 -54.235 ;
        RECT -65.445 -55.925 -65.115 -55.595 ;
        RECT -65.445 -57.285 -65.115 -56.955 ;
        RECT -65.445 -58.645 -65.115 -58.315 ;
        RECT -65.445 -60.005 -65.115 -59.675 ;
        RECT -65.445 -61.365 -65.115 -61.035 ;
        RECT -65.445 -62.725 -65.115 -62.395 ;
        RECT -65.445 -64.085 -65.115 -63.755 ;
        RECT -65.445 -65.445 -65.115 -65.115 ;
        RECT -65.445 -66.805 -65.115 -66.475 ;
        RECT -65.445 -68.165 -65.115 -67.835 ;
        RECT -65.445 -69.525 -65.115 -69.195 ;
        RECT -65.445 -70.885 -65.115 -70.555 ;
        RECT -65.445 -72.245 -65.115 -71.915 ;
        RECT -65.445 -73.605 -65.115 -73.275 ;
        RECT -65.445 -74.965 -65.115 -74.635 ;
        RECT -65.445 -76.325 -65.115 -75.995 ;
        RECT -65.445 -77.685 -65.115 -77.355 ;
        RECT -65.445 -79.045 -65.115 -78.715 ;
        RECT -65.445 -80.405 -65.115 -80.075 ;
        RECT -65.445 -81.765 -65.115 -81.435 ;
        RECT -65.445 -83.125 -65.115 -82.795 ;
        RECT -65.445 -84.485 -65.115 -84.155 ;
        RECT -65.445 -85.845 -65.115 -85.515 ;
        RECT -65.445 -87.205 -65.115 -86.875 ;
        RECT -65.445 -88.565 -65.115 -88.235 ;
        RECT -65.445 -89.925 -65.115 -89.595 ;
        RECT -65.445 -91.285 -65.115 -90.955 ;
        RECT -65.445 -92.645 -65.115 -92.315 ;
        RECT -65.445 -94.005 -65.115 -93.675 ;
        RECT -65.445 -95.365 -65.115 -95.035 ;
        RECT -65.445 -96.725 -65.115 -96.395 ;
        RECT -65.445 -98.085 -65.115 -97.755 ;
        RECT -65.445 -99.445 -65.115 -99.115 ;
        RECT -65.445 -100.805 -65.115 -100.475 ;
        RECT -65.445 -102.165 -65.115 -101.835 ;
        RECT -65.445 -103.525 -65.115 -103.195 ;
        RECT -65.445 -104.885 -65.115 -104.555 ;
        RECT -65.445 -106.245 -65.115 -105.915 ;
        RECT -65.445 -107.605 -65.115 -107.275 ;
        RECT -65.445 -108.965 -65.115 -108.635 ;
        RECT -65.445 -110.325 -65.115 -109.995 ;
        RECT -65.445 -111.685 -65.115 -111.355 ;
        RECT -65.445 -113.045 -65.115 -112.715 ;
        RECT -65.445 -114.405 -65.115 -114.075 ;
        RECT -65.445 -115.765 -65.115 -115.435 ;
        RECT -65.445 -117.125 -65.115 -116.795 ;
        RECT -65.445 -118.485 -65.115 -118.155 ;
        RECT -65.445 -119.845 -65.115 -119.515 ;
        RECT -65.445 -121.205 -65.115 -120.875 ;
        RECT -65.445 -122.565 -65.115 -122.235 ;
        RECT -65.445 -123.925 -65.115 -123.595 ;
        RECT -65.445 -125.285 -65.115 -124.955 ;
        RECT -65.445 -126.645 -65.115 -126.315 ;
        RECT -65.445 -128.005 -65.115 -127.675 ;
        RECT -65.445 -129.365 -65.115 -129.035 ;
        RECT -65.445 -130.725 -65.115 -130.395 ;
        RECT -65.445 -132.085 -65.115 -131.755 ;
        RECT -65.445 -133.445 -65.115 -133.115 ;
        RECT -65.445 -134.805 -65.115 -134.475 ;
        RECT -65.445 -136.165 -65.115 -135.835 ;
        RECT -65.445 -137.525 -65.115 -137.195 ;
        RECT -65.445 -138.885 -65.115 -138.555 ;
        RECT -65.445 -140.245 -65.115 -139.915 ;
        RECT -65.445 -141.605 -65.115 -141.275 ;
        RECT -65.445 -142.965 -65.115 -142.635 ;
        RECT -65.445 -144.325 -65.115 -143.995 ;
        RECT -65.445 -145.685 -65.115 -145.355 ;
        RECT -65.445 -147.045 -65.115 -146.715 ;
        RECT -65.445 -148.405 -65.115 -148.075 ;
        RECT -65.445 -149.765 -65.115 -149.435 ;
        RECT -65.445 -151.125 -65.115 -150.795 ;
        RECT -65.445 -152.485 -65.115 -152.155 ;
        RECT -65.445 -153.845 -65.115 -153.515 ;
        RECT -65.445 -155.205 -65.115 -154.875 ;
        RECT -65.445 -156.565 -65.115 -156.235 ;
        RECT -65.445 -157.925 -65.115 -157.595 ;
        RECT -65.445 -159.285 -65.115 -158.955 ;
        RECT -65.445 -160.645 -65.115 -160.315 ;
        RECT -65.445 -162.005 -65.115 -161.675 ;
        RECT -65.445 -163.365 -65.115 -163.035 ;
        RECT -65.445 -164.725 -65.115 -164.395 ;
        RECT -65.445 -166.085 -65.115 -165.755 ;
        RECT -65.445 -167.445 -65.115 -167.115 ;
        RECT -65.445 -170.165 -65.115 -169.835 ;
        RECT -65.445 -174.245 -65.115 -173.915 ;
        RECT -65.445 -175.725 -65.115 -175.395 ;
        RECT -65.445 -176.965 -65.115 -176.635 ;
        RECT -65.445 -178.325 -65.115 -177.995 ;
        RECT -65.445 -180.57 -65.115 -179.44 ;
        RECT -65.44 -180.685 -65.12 242.565 ;
        RECT -65.445 241.32 -65.115 242.45 ;
        RECT -65.445 239.195 -65.115 239.525 ;
        RECT -65.445 237.835 -65.115 238.165 ;
        RECT -65.445 236.475 -65.115 236.805 ;
        RECT -65.445 235.115 -65.115 235.445 ;
        RECT -65.445 233.755 -65.115 234.085 ;
        RECT -65.445 232.395 -65.115 232.725 ;
        RECT -65.445 231.035 -65.115 231.365 ;
        RECT -65.445 229.675 -65.115 230.005 ;
        RECT -65.445 228.315 -65.115 228.645 ;
        RECT -65.445 226.955 -65.115 227.285 ;
        RECT -65.445 225.595 -65.115 225.925 ;
        RECT -65.445 224.235 -65.115 224.565 ;
        RECT -65.445 222.875 -65.115 223.205 ;
        RECT -65.445 221.515 -65.115 221.845 ;
        RECT -65.445 220.155 -65.115 220.485 ;
        RECT -65.445 218.795 -65.115 219.125 ;
        RECT -65.445 217.435 -65.115 217.765 ;
        RECT -65.445 216.075 -65.115 216.405 ;
        RECT -65.445 214.715 -65.115 215.045 ;
        RECT -65.445 213.355 -65.115 213.685 ;
        RECT -65.445 211.995 -65.115 212.325 ;
        RECT -65.445 210.635 -65.115 210.965 ;
        RECT -65.445 209.275 -65.115 209.605 ;
        RECT -65.445 207.915 -65.115 208.245 ;
        RECT -65.445 206.555 -65.115 206.885 ;
        RECT -65.445 205.195 -65.115 205.525 ;
        RECT -65.445 203.835 -65.115 204.165 ;
        RECT -65.445 202.475 -65.115 202.805 ;
        RECT -65.445 201.115 -65.115 201.445 ;
        RECT -65.445 199.755 -65.115 200.085 ;
        RECT -65.445 198.395 -65.115 198.725 ;
        RECT -65.445 197.035 -65.115 197.365 ;
        RECT -65.445 195.675 -65.115 196.005 ;
        RECT -65.445 194.315 -65.115 194.645 ;
        RECT -65.445 192.955 -65.115 193.285 ;
        RECT -65.445 191.595 -65.115 191.925 ;
        RECT -65.445 190.235 -65.115 190.565 ;
        RECT -65.445 188.875 -65.115 189.205 ;
        RECT -65.445 187.515 -65.115 187.845 ;
        RECT -65.445 186.155 -65.115 186.485 ;
        RECT -65.445 184.795 -65.115 185.125 ;
        RECT -65.445 183.435 -65.115 183.765 ;
        RECT -65.445 182.075 -65.115 182.405 ;
        RECT -65.445 180.715 -65.115 181.045 ;
        RECT -65.445 179.355 -65.115 179.685 ;
        RECT -65.445 177.995 -65.115 178.325 ;
        RECT -65.445 176.635 -65.115 176.965 ;
        RECT -65.445 175.275 -65.115 175.605 ;
        RECT -65.445 173.915 -65.115 174.245 ;
        RECT -65.445 172.555 -65.115 172.885 ;
        RECT -65.445 171.195 -65.115 171.525 ;
        RECT -65.445 169.835 -65.115 170.165 ;
        RECT -65.445 168.475 -65.115 168.805 ;
        RECT -65.445 167.115 -65.115 167.445 ;
        RECT -65.445 165.755 -65.115 166.085 ;
        RECT -65.445 164.395 -65.115 164.725 ;
        RECT -65.445 163.035 -65.115 163.365 ;
        RECT -65.445 161.675 -65.115 162.005 ;
        RECT -65.445 160.315 -65.115 160.645 ;
        RECT -65.445 158.955 -65.115 159.285 ;
        RECT -65.445 157.595 -65.115 157.925 ;
        RECT -65.445 156.235 -65.115 156.565 ;
        RECT -65.445 154.875 -65.115 155.205 ;
        RECT -65.445 153.515 -65.115 153.845 ;
        RECT -65.445 152.155 -65.115 152.485 ;
        RECT -65.445 150.795 -65.115 151.125 ;
        RECT -65.445 149.435 -65.115 149.765 ;
        RECT -65.445 148.075 -65.115 148.405 ;
        RECT -65.445 146.715 -65.115 147.045 ;
        RECT -65.445 145.355 -65.115 145.685 ;
        RECT -65.445 143.995 -65.115 144.325 ;
        RECT -65.445 142.635 -65.115 142.965 ;
        RECT -65.445 141.275 -65.115 141.605 ;
        RECT -65.445 139.915 -65.115 140.245 ;
        RECT -65.445 138.555 -65.115 138.885 ;
        RECT -65.445 137.195 -65.115 137.525 ;
        RECT -65.445 135.835 -65.115 136.165 ;
        RECT -65.445 134.475 -65.115 134.805 ;
        RECT -65.445 133.115 -65.115 133.445 ;
        RECT -65.445 131.755 -65.115 132.085 ;
        RECT -65.445 130.395 -65.115 130.725 ;
        RECT -65.445 129.035 -65.115 129.365 ;
        RECT -65.445 127.675 -65.115 128.005 ;
        RECT -65.445 126.315 -65.115 126.645 ;
        RECT -65.445 124.955 -65.115 125.285 ;
        RECT -65.445 123.595 -65.115 123.925 ;
        RECT -65.445 122.235 -65.115 122.565 ;
        RECT -65.445 120.875 -65.115 121.205 ;
        RECT -65.445 119.515 -65.115 119.845 ;
        RECT -65.445 118.155 -65.115 118.485 ;
        RECT -65.445 116.795 -65.115 117.125 ;
        RECT -65.445 115.435 -65.115 115.765 ;
        RECT -65.445 114.075 -65.115 114.405 ;
        RECT -65.445 112.715 -65.115 113.045 ;
        RECT -65.445 111.355 -65.115 111.685 ;
        RECT -65.445 109.995 -65.115 110.325 ;
        RECT -65.445 108.635 -65.115 108.965 ;
        RECT -65.445 107.275 -65.115 107.605 ;
        RECT -65.445 105.915 -65.115 106.245 ;
        RECT -65.445 104.555 -65.115 104.885 ;
        RECT -65.445 103.195 -65.115 103.525 ;
        RECT -65.445 101.835 -65.115 102.165 ;
        RECT -65.445 100.475 -65.115 100.805 ;
        RECT -65.445 99.115 -65.115 99.445 ;
        RECT -65.445 97.755 -65.115 98.085 ;
        RECT -65.445 96.395 -65.115 96.725 ;
        RECT -65.445 95.035 -65.115 95.365 ;
        RECT -65.445 93.675 -65.115 94.005 ;
        RECT -65.445 92.315 -65.115 92.645 ;
        RECT -65.445 90.955 -65.115 91.285 ;
        RECT -65.445 89.595 -65.115 89.925 ;
        RECT -65.445 88.235 -65.115 88.565 ;
        RECT -65.445 86.875 -65.115 87.205 ;
        RECT -65.445 85.515 -65.115 85.845 ;
        RECT -65.445 84.155 -65.115 84.485 ;
        RECT -65.445 82.795 -65.115 83.125 ;
        RECT -65.445 81.435 -65.115 81.765 ;
        RECT -65.445 80.075 -65.115 80.405 ;
        RECT -65.445 78.715 -65.115 79.045 ;
        RECT -65.445 77.355 -65.115 77.685 ;
        RECT -65.445 75.995 -65.115 76.325 ;
        RECT -65.445 74.635 -65.115 74.965 ;
        RECT -65.445 73.275 -65.115 73.605 ;
        RECT -65.445 71.915 -65.115 72.245 ;
        RECT -65.445 70.555 -65.115 70.885 ;
        RECT -65.445 69.195 -65.115 69.525 ;
        RECT -65.445 67.835 -65.115 68.165 ;
        RECT -65.445 66.475 -65.115 66.805 ;
        RECT -65.445 65.115 -65.115 65.445 ;
        RECT -65.445 63.755 -65.115 64.085 ;
        RECT -65.445 62.395 -65.115 62.725 ;
        RECT -65.445 61.035 -65.115 61.365 ;
        RECT -65.445 59.675 -65.115 60.005 ;
        RECT -65.445 58.315 -65.115 58.645 ;
        RECT -65.445 56.955 -65.115 57.285 ;
        RECT -65.445 55.595 -65.115 55.925 ;
        RECT -65.445 54.235 -65.115 54.565 ;
        RECT -65.445 52.875 -65.115 53.205 ;
        RECT -65.445 51.515 -65.115 51.845 ;
        RECT -65.445 50.155 -65.115 50.485 ;
        RECT -65.445 48.795 -65.115 49.125 ;
        RECT -65.445 47.435 -65.115 47.765 ;
        RECT -65.445 46.075 -65.115 46.405 ;
        RECT -65.445 44.715 -65.115 45.045 ;
        RECT -65.445 43.355 -65.115 43.685 ;
        RECT -65.445 41.995 -65.115 42.325 ;
        RECT -65.445 40.635 -65.115 40.965 ;
        RECT -65.445 39.275 -65.115 39.605 ;
        RECT -65.445 37.915 -65.115 38.245 ;
        RECT -65.445 36.555 -65.115 36.885 ;
        RECT -65.445 35.195 -65.115 35.525 ;
        RECT -65.445 33.835 -65.115 34.165 ;
        RECT -65.445 32.475 -65.115 32.805 ;
        RECT -65.445 31.115 -65.115 31.445 ;
        RECT -65.445 29.755 -65.115 30.085 ;
        RECT -65.445 28.395 -65.115 28.725 ;
        RECT -65.445 27.035 -65.115 27.365 ;
        RECT -65.445 25.675 -65.115 26.005 ;
        RECT -65.445 24.315 -65.115 24.645 ;
        RECT -65.445 22.955 -65.115 23.285 ;
        RECT -65.445 21.595 -65.115 21.925 ;
        RECT -65.445 20.235 -65.115 20.565 ;
        RECT -65.445 18.875 -65.115 19.205 ;
        RECT -65.445 17.515 -65.115 17.845 ;
        RECT -65.445 16.155 -65.115 16.485 ;
        RECT -65.445 14.795 -65.115 15.125 ;
        RECT -65.445 13.435 -65.115 13.765 ;
        RECT -65.445 12.075 -65.115 12.405 ;
        RECT -65.445 10.715 -65.115 11.045 ;
        RECT -65.445 9.355 -65.115 9.685 ;
        RECT -65.445 7.995 -65.115 8.325 ;
        RECT -65.445 6.635 -65.115 6.965 ;
        RECT -65.445 5.275 -65.115 5.605 ;
        RECT -65.445 3.915 -65.115 4.245 ;
        RECT -65.445 2.555 -65.115 2.885 ;
        RECT -65.445 1.195 -65.115 1.525 ;
    END
    PORT
      LAYER met3 ;
        RECT -73.605 241.32 -73.275 242.45 ;
        RECT -73.605 239.195 -73.275 239.525 ;
        RECT -73.605 237.835 -73.275 238.165 ;
        RECT -73.605 236.475 -73.275 236.805 ;
        RECT -73.605 235.115 -73.275 235.445 ;
        RECT -73.605 233.755 -73.275 234.085 ;
        RECT -73.605 232.395 -73.275 232.725 ;
        RECT -73.605 231.035 -73.275 231.365 ;
        RECT -73.605 229.675 -73.275 230.005 ;
        RECT -73.605 228.315 -73.275 228.645 ;
        RECT -73.605 226.955 -73.275 227.285 ;
        RECT -73.605 225.595 -73.275 225.925 ;
        RECT -73.605 224.235 -73.275 224.565 ;
        RECT -73.605 222.875 -73.275 223.205 ;
        RECT -73.605 221.515 -73.275 221.845 ;
        RECT -73.605 220.155 -73.275 220.485 ;
        RECT -73.605 218.795 -73.275 219.125 ;
        RECT -73.605 217.435 -73.275 217.765 ;
        RECT -73.605 216.075 -73.275 216.405 ;
        RECT -73.605 214.715 -73.275 215.045 ;
        RECT -73.605 213.355 -73.275 213.685 ;
        RECT -73.605 211.995 -73.275 212.325 ;
        RECT -73.605 210.635 -73.275 210.965 ;
        RECT -73.605 209.275 -73.275 209.605 ;
        RECT -73.605 207.915 -73.275 208.245 ;
        RECT -73.605 206.555 -73.275 206.885 ;
        RECT -73.605 205.195 -73.275 205.525 ;
        RECT -73.605 203.835 -73.275 204.165 ;
        RECT -73.605 202.475 -73.275 202.805 ;
        RECT -73.605 201.115 -73.275 201.445 ;
        RECT -73.605 199.755 -73.275 200.085 ;
        RECT -73.605 198.395 -73.275 198.725 ;
        RECT -73.605 197.035 -73.275 197.365 ;
        RECT -73.605 195.675 -73.275 196.005 ;
        RECT -73.605 194.315 -73.275 194.645 ;
        RECT -73.605 192.955 -73.275 193.285 ;
        RECT -73.605 191.595 -73.275 191.925 ;
        RECT -73.605 190.235 -73.275 190.565 ;
        RECT -73.605 188.875 -73.275 189.205 ;
        RECT -73.605 187.515 -73.275 187.845 ;
        RECT -73.605 186.155 -73.275 186.485 ;
        RECT -73.605 184.795 -73.275 185.125 ;
        RECT -73.605 183.435 -73.275 183.765 ;
        RECT -73.605 182.075 -73.275 182.405 ;
        RECT -73.605 180.715 -73.275 181.045 ;
        RECT -73.605 179.355 -73.275 179.685 ;
        RECT -73.605 177.995 -73.275 178.325 ;
        RECT -73.605 176.635 -73.275 176.965 ;
        RECT -73.605 175.275 -73.275 175.605 ;
        RECT -73.605 173.915 -73.275 174.245 ;
        RECT -73.605 172.555 -73.275 172.885 ;
        RECT -73.605 171.195 -73.275 171.525 ;
        RECT -73.605 169.835 -73.275 170.165 ;
        RECT -73.605 168.475 -73.275 168.805 ;
        RECT -73.605 167.115 -73.275 167.445 ;
        RECT -73.605 165.755 -73.275 166.085 ;
        RECT -73.605 164.395 -73.275 164.725 ;
        RECT -73.605 163.035 -73.275 163.365 ;
        RECT -73.605 161.675 -73.275 162.005 ;
        RECT -73.605 160.315 -73.275 160.645 ;
        RECT -73.605 158.955 -73.275 159.285 ;
        RECT -73.605 157.595 -73.275 157.925 ;
        RECT -73.605 156.235 -73.275 156.565 ;
        RECT -73.605 154.875 -73.275 155.205 ;
        RECT -73.605 153.515 -73.275 153.845 ;
        RECT -73.605 152.155 -73.275 152.485 ;
        RECT -73.605 150.795 -73.275 151.125 ;
        RECT -73.605 149.435 -73.275 149.765 ;
        RECT -73.605 148.075 -73.275 148.405 ;
        RECT -73.605 146.715 -73.275 147.045 ;
        RECT -73.605 145.355 -73.275 145.685 ;
        RECT -73.605 143.995 -73.275 144.325 ;
        RECT -73.605 142.635 -73.275 142.965 ;
        RECT -73.605 141.275 -73.275 141.605 ;
        RECT -73.605 139.915 -73.275 140.245 ;
        RECT -73.605 138.555 -73.275 138.885 ;
        RECT -73.605 137.195 -73.275 137.525 ;
        RECT -73.605 135.835 -73.275 136.165 ;
        RECT -73.605 134.475 -73.275 134.805 ;
        RECT -73.605 133.115 -73.275 133.445 ;
        RECT -73.605 131.755 -73.275 132.085 ;
        RECT -73.605 130.395 -73.275 130.725 ;
        RECT -73.605 129.035 -73.275 129.365 ;
        RECT -73.605 127.675 -73.275 128.005 ;
        RECT -73.605 126.315 -73.275 126.645 ;
        RECT -73.605 124.955 -73.275 125.285 ;
        RECT -73.605 123.595 -73.275 123.925 ;
        RECT -73.605 122.235 -73.275 122.565 ;
        RECT -73.605 120.875 -73.275 121.205 ;
        RECT -73.605 119.515 -73.275 119.845 ;
        RECT -73.605 118.155 -73.275 118.485 ;
        RECT -73.605 116.795 -73.275 117.125 ;
        RECT -73.605 115.435 -73.275 115.765 ;
        RECT -73.605 114.075 -73.275 114.405 ;
        RECT -73.605 112.715 -73.275 113.045 ;
        RECT -73.605 111.355 -73.275 111.685 ;
        RECT -73.605 109.995 -73.275 110.325 ;
        RECT -73.605 108.635 -73.275 108.965 ;
        RECT -73.605 107.275 -73.275 107.605 ;
        RECT -73.605 105.915 -73.275 106.245 ;
        RECT -73.605 104.555 -73.275 104.885 ;
        RECT -73.605 103.195 -73.275 103.525 ;
        RECT -73.605 101.835 -73.275 102.165 ;
        RECT -73.605 100.475 -73.275 100.805 ;
        RECT -73.605 99.115 -73.275 99.445 ;
        RECT -73.605 97.755 -73.275 98.085 ;
        RECT -73.605 96.395 -73.275 96.725 ;
        RECT -73.605 95.035 -73.275 95.365 ;
        RECT -73.605 93.675 -73.275 94.005 ;
        RECT -73.605 92.315 -73.275 92.645 ;
        RECT -73.605 90.955 -73.275 91.285 ;
        RECT -73.605 89.595 -73.275 89.925 ;
        RECT -73.605 88.235 -73.275 88.565 ;
        RECT -73.605 86.875 -73.275 87.205 ;
        RECT -73.605 85.515 -73.275 85.845 ;
        RECT -73.605 84.155 -73.275 84.485 ;
        RECT -73.605 82.795 -73.275 83.125 ;
        RECT -73.605 81.435 -73.275 81.765 ;
        RECT -73.605 80.075 -73.275 80.405 ;
        RECT -73.605 78.715 -73.275 79.045 ;
        RECT -73.605 77.355 -73.275 77.685 ;
        RECT -73.605 75.995 -73.275 76.325 ;
        RECT -73.605 74.635 -73.275 74.965 ;
        RECT -73.605 73.275 -73.275 73.605 ;
        RECT -73.605 71.915 -73.275 72.245 ;
        RECT -73.605 70.555 -73.275 70.885 ;
        RECT -73.605 69.195 -73.275 69.525 ;
        RECT -73.605 67.835 -73.275 68.165 ;
        RECT -73.605 66.475 -73.275 66.805 ;
        RECT -73.605 65.115 -73.275 65.445 ;
        RECT -73.605 63.755 -73.275 64.085 ;
        RECT -73.605 62.395 -73.275 62.725 ;
        RECT -73.605 61.035 -73.275 61.365 ;
        RECT -73.605 59.675 -73.275 60.005 ;
        RECT -73.605 58.315 -73.275 58.645 ;
        RECT -73.605 56.955 -73.275 57.285 ;
        RECT -73.605 55.595 -73.275 55.925 ;
        RECT -73.605 54.235 -73.275 54.565 ;
        RECT -73.605 52.875 -73.275 53.205 ;
        RECT -73.605 51.515 -73.275 51.845 ;
        RECT -73.605 50.155 -73.275 50.485 ;
        RECT -73.605 48.795 -73.275 49.125 ;
        RECT -73.605 47.435 -73.275 47.765 ;
        RECT -73.605 46.075 -73.275 46.405 ;
        RECT -73.605 44.715 -73.275 45.045 ;
        RECT -73.605 43.355 -73.275 43.685 ;
        RECT -73.605 41.995 -73.275 42.325 ;
        RECT -73.605 40.635 -73.275 40.965 ;
        RECT -73.605 39.275 -73.275 39.605 ;
        RECT -73.605 37.915 -73.275 38.245 ;
        RECT -73.605 36.555 -73.275 36.885 ;
        RECT -73.605 35.195 -73.275 35.525 ;
        RECT -73.605 33.835 -73.275 34.165 ;
        RECT -73.605 32.475 -73.275 32.805 ;
        RECT -73.605 31.115 -73.275 31.445 ;
        RECT -73.605 29.755 -73.275 30.085 ;
        RECT -73.605 28.395 -73.275 28.725 ;
        RECT -73.605 27.035 -73.275 27.365 ;
        RECT -73.605 25.675 -73.275 26.005 ;
        RECT -73.605 24.315 -73.275 24.645 ;
        RECT -73.605 22.955 -73.275 23.285 ;
        RECT -73.605 21.595 -73.275 21.925 ;
        RECT -73.605 20.235 -73.275 20.565 ;
        RECT -73.605 18.875 -73.275 19.205 ;
        RECT -73.605 17.515 -73.275 17.845 ;
        RECT -73.605 16.155 -73.275 16.485 ;
        RECT -73.605 14.795 -73.275 15.125 ;
        RECT -73.605 13.435 -73.275 13.765 ;
        RECT -73.605 12.075 -73.275 12.405 ;
        RECT -73.605 10.715 -73.275 11.045 ;
        RECT -73.605 9.355 -73.275 9.685 ;
        RECT -73.605 7.995 -73.275 8.325 ;
        RECT -73.605 6.635 -73.275 6.965 ;
        RECT -73.605 5.275 -73.275 5.605 ;
        RECT -73.605 3.915 -73.275 4.245 ;
        RECT -73.605 2.555 -73.275 2.885 ;
        RECT -73.605 1.195 -73.275 1.525 ;
        RECT -73.605 -0.165 -73.275 0.165 ;
        RECT -73.605 -1.525 -73.275 -1.195 ;
        RECT -73.605 -2.885 -73.275 -2.555 ;
        RECT -73.605 -4.245 -73.275 -3.915 ;
        RECT -73.605 -5.605 -73.275 -5.275 ;
        RECT -73.605 -6.965 -73.275 -6.635 ;
        RECT -73.605 -8.325 -73.275 -7.995 ;
        RECT -73.605 -9.685 -73.275 -9.355 ;
        RECT -73.605 -11.045 -73.275 -10.715 ;
        RECT -73.605 -12.405 -73.275 -12.075 ;
        RECT -73.605 -13.765 -73.275 -13.435 ;
        RECT -73.605 -15.125 -73.275 -14.795 ;
        RECT -73.605 -16.485 -73.275 -16.155 ;
        RECT -73.605 -17.845 -73.275 -17.515 ;
        RECT -73.605 -19.205 -73.275 -18.875 ;
        RECT -73.605 -20.565 -73.275 -20.235 ;
        RECT -73.605 -21.925 -73.275 -21.595 ;
        RECT -73.605 -23.285 -73.275 -22.955 ;
        RECT -73.605 -24.645 -73.275 -24.315 ;
        RECT -73.605 -26.005 -73.275 -25.675 ;
        RECT -73.605 -27.365 -73.275 -27.035 ;
        RECT -73.605 -28.725 -73.275 -28.395 ;
        RECT -73.605 -30.085 -73.275 -29.755 ;
        RECT -73.605 -31.445 -73.275 -31.115 ;
        RECT -73.605 -32.805 -73.275 -32.475 ;
        RECT -73.605 -34.165 -73.275 -33.835 ;
        RECT -73.605 -35.525 -73.275 -35.195 ;
        RECT -73.605 -36.885 -73.275 -36.555 ;
        RECT -73.605 -38.245 -73.275 -37.915 ;
        RECT -73.605 -39.605 -73.275 -39.275 ;
        RECT -73.605 -40.965 -73.275 -40.635 ;
        RECT -73.605 -42.325 -73.275 -41.995 ;
        RECT -73.605 -43.685 -73.275 -43.355 ;
        RECT -73.605 -45.045 -73.275 -44.715 ;
        RECT -73.605 -46.405 -73.275 -46.075 ;
        RECT -73.605 -47.765 -73.275 -47.435 ;
        RECT -73.605 -49.125 -73.275 -48.795 ;
        RECT -73.605 -50.485 -73.275 -50.155 ;
        RECT -73.605 -51.845 -73.275 -51.515 ;
        RECT -73.605 -53.205 -73.275 -52.875 ;
        RECT -73.605 -54.565 -73.275 -54.235 ;
        RECT -73.605 -55.925 -73.275 -55.595 ;
        RECT -73.605 -57.285 -73.275 -56.955 ;
        RECT -73.605 -58.645 -73.275 -58.315 ;
        RECT -73.605 -60.005 -73.275 -59.675 ;
        RECT -73.605 -61.365 -73.275 -61.035 ;
        RECT -73.605 -62.725 -73.275 -62.395 ;
        RECT -73.605 -64.085 -73.275 -63.755 ;
        RECT -73.605 -65.445 -73.275 -65.115 ;
        RECT -73.605 -66.805 -73.275 -66.475 ;
        RECT -73.605 -68.165 -73.275 -67.835 ;
        RECT -73.605 -69.525 -73.275 -69.195 ;
        RECT -73.605 -70.885 -73.275 -70.555 ;
        RECT -73.605 -72.245 -73.275 -71.915 ;
        RECT -73.605 -73.605 -73.275 -73.275 ;
        RECT -73.605 -74.965 -73.275 -74.635 ;
        RECT -73.605 -76.325 -73.275 -75.995 ;
        RECT -73.605 -77.685 -73.275 -77.355 ;
        RECT -73.605 -79.045 -73.275 -78.715 ;
        RECT -73.605 -80.405 -73.275 -80.075 ;
        RECT -73.605 -81.765 -73.275 -81.435 ;
        RECT -73.605 -83.125 -73.275 -82.795 ;
        RECT -73.605 -84.485 -73.275 -84.155 ;
        RECT -73.605 -85.845 -73.275 -85.515 ;
        RECT -73.605 -87.205 -73.275 -86.875 ;
        RECT -73.605 -88.565 -73.275 -88.235 ;
        RECT -73.605 -89.925 -73.275 -89.595 ;
        RECT -73.605 -91.285 -73.275 -90.955 ;
        RECT -73.605 -92.645 -73.275 -92.315 ;
        RECT -73.605 -94.005 -73.275 -93.675 ;
        RECT -73.605 -95.365 -73.275 -95.035 ;
        RECT -73.605 -96.725 -73.275 -96.395 ;
        RECT -73.605 -98.085 -73.275 -97.755 ;
        RECT -73.605 -99.445 -73.275 -99.115 ;
        RECT -73.605 -100.805 -73.275 -100.475 ;
        RECT -73.605 -102.165 -73.275 -101.835 ;
        RECT -73.605 -103.525 -73.275 -103.195 ;
        RECT -73.605 -104.885 -73.275 -104.555 ;
        RECT -73.605 -106.245 -73.275 -105.915 ;
        RECT -73.605 -107.605 -73.275 -107.275 ;
        RECT -73.605 -108.965 -73.275 -108.635 ;
        RECT -73.605 -110.325 -73.275 -109.995 ;
        RECT -73.605 -111.685 -73.275 -111.355 ;
        RECT -73.605 -113.045 -73.275 -112.715 ;
        RECT -73.605 -114.405 -73.275 -114.075 ;
        RECT -73.605 -115.765 -73.275 -115.435 ;
        RECT -73.605 -117.125 -73.275 -116.795 ;
        RECT -73.605 -118.485 -73.275 -118.155 ;
        RECT -73.605 -119.845 -73.275 -119.515 ;
        RECT -73.605 -121.205 -73.275 -120.875 ;
        RECT -73.605 -122.565 -73.275 -122.235 ;
        RECT -73.605 -123.925 -73.275 -123.595 ;
        RECT -73.605 -125.285 -73.275 -124.955 ;
        RECT -73.605 -126.645 -73.275 -126.315 ;
        RECT -73.605 -128.005 -73.275 -127.675 ;
        RECT -73.605 -129.365 -73.275 -129.035 ;
        RECT -73.605 -130.725 -73.275 -130.395 ;
        RECT -73.605 -132.085 -73.275 -131.755 ;
        RECT -73.605 -133.445 -73.275 -133.115 ;
        RECT -73.605 -134.805 -73.275 -134.475 ;
        RECT -73.605 -136.165 -73.275 -135.835 ;
        RECT -73.605 -137.525 -73.275 -137.195 ;
        RECT -73.605 -138.885 -73.275 -138.555 ;
        RECT -73.605 -140.245 -73.275 -139.915 ;
        RECT -73.605 -141.605 -73.275 -141.275 ;
        RECT -73.605 -142.965 -73.275 -142.635 ;
        RECT -73.605 -144.325 -73.275 -143.995 ;
        RECT -73.605 -145.685 -73.275 -145.355 ;
        RECT -73.605 -147.045 -73.275 -146.715 ;
        RECT -73.605 -148.405 -73.275 -148.075 ;
        RECT -73.605 -149.765 -73.275 -149.435 ;
        RECT -73.605 -151.125 -73.275 -150.795 ;
        RECT -73.605 -152.485 -73.275 -152.155 ;
        RECT -73.605 -153.845 -73.275 -153.515 ;
        RECT -73.605 -155.205 -73.275 -154.875 ;
        RECT -73.605 -156.565 -73.275 -156.235 ;
        RECT -73.605 -157.925 -73.275 -157.595 ;
        RECT -73.605 -159.285 -73.275 -158.955 ;
        RECT -73.605 -160.645 -73.275 -160.315 ;
        RECT -73.605 -162.005 -73.275 -161.675 ;
        RECT -73.605 -163.365 -73.275 -163.035 ;
        RECT -73.605 -164.725 -73.275 -164.395 ;
        RECT -73.605 -166.085 -73.275 -165.755 ;
        RECT -73.605 -167.445 -73.275 -167.115 ;
        RECT -73.605 -168.805 -73.275 -168.475 ;
        RECT -73.605 -170.165 -73.275 -169.835 ;
        RECT -73.605 -171.525 -73.275 -171.195 ;
        RECT -73.605 -172.885 -73.275 -172.555 ;
        RECT -73.605 -174.245 -73.275 -173.915 ;
        RECT -73.605 -175.605 -73.275 -175.275 ;
        RECT -73.605 -176.965 -73.275 -176.635 ;
        RECT -73.605 -178.325 -73.275 -177.995 ;
        RECT -73.605 -180.57 -73.275 -179.44 ;
        RECT -73.6 -180.685 -73.28 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -72.245 241.32 -71.915 242.45 ;
        RECT -72.245 239.195 -71.915 239.525 ;
        RECT -72.245 237.835 -71.915 238.165 ;
        RECT -72.245 236.475 -71.915 236.805 ;
        RECT -72.245 235.115 -71.915 235.445 ;
        RECT -72.245 233.755 -71.915 234.085 ;
        RECT -72.245 232.395 -71.915 232.725 ;
        RECT -72.245 231.035 -71.915 231.365 ;
        RECT -72.245 229.675 -71.915 230.005 ;
        RECT -72.245 228.315 -71.915 228.645 ;
        RECT -72.245 226.955 -71.915 227.285 ;
        RECT -72.245 225.595 -71.915 225.925 ;
        RECT -72.245 224.235 -71.915 224.565 ;
        RECT -72.245 222.875 -71.915 223.205 ;
        RECT -72.245 221.515 -71.915 221.845 ;
        RECT -72.245 220.155 -71.915 220.485 ;
        RECT -72.245 218.795 -71.915 219.125 ;
        RECT -72.245 217.435 -71.915 217.765 ;
        RECT -72.245 216.075 -71.915 216.405 ;
        RECT -72.245 214.715 -71.915 215.045 ;
        RECT -72.245 213.355 -71.915 213.685 ;
        RECT -72.245 211.995 -71.915 212.325 ;
        RECT -72.245 210.635 -71.915 210.965 ;
        RECT -72.245 209.275 -71.915 209.605 ;
        RECT -72.245 207.915 -71.915 208.245 ;
        RECT -72.245 206.555 -71.915 206.885 ;
        RECT -72.245 205.195 -71.915 205.525 ;
        RECT -72.245 203.835 -71.915 204.165 ;
        RECT -72.245 202.475 -71.915 202.805 ;
        RECT -72.245 201.115 -71.915 201.445 ;
        RECT -72.245 199.755 -71.915 200.085 ;
        RECT -72.245 198.395 -71.915 198.725 ;
        RECT -72.245 197.035 -71.915 197.365 ;
        RECT -72.245 195.675 -71.915 196.005 ;
        RECT -72.245 194.315 -71.915 194.645 ;
        RECT -72.245 192.955 -71.915 193.285 ;
        RECT -72.245 191.595 -71.915 191.925 ;
        RECT -72.245 190.235 -71.915 190.565 ;
        RECT -72.245 188.875 -71.915 189.205 ;
        RECT -72.245 187.515 -71.915 187.845 ;
        RECT -72.245 186.155 -71.915 186.485 ;
        RECT -72.245 184.795 -71.915 185.125 ;
        RECT -72.245 183.435 -71.915 183.765 ;
        RECT -72.245 182.075 -71.915 182.405 ;
        RECT -72.245 180.715 -71.915 181.045 ;
        RECT -72.245 179.355 -71.915 179.685 ;
        RECT -72.245 177.995 -71.915 178.325 ;
        RECT -72.245 176.635 -71.915 176.965 ;
        RECT -72.245 175.275 -71.915 175.605 ;
        RECT -72.245 173.915 -71.915 174.245 ;
        RECT -72.245 172.555 -71.915 172.885 ;
        RECT -72.245 171.195 -71.915 171.525 ;
        RECT -72.245 169.835 -71.915 170.165 ;
        RECT -72.245 168.475 -71.915 168.805 ;
        RECT -72.245 167.115 -71.915 167.445 ;
        RECT -72.245 165.755 -71.915 166.085 ;
        RECT -72.245 164.395 -71.915 164.725 ;
        RECT -72.245 163.035 -71.915 163.365 ;
        RECT -72.245 161.675 -71.915 162.005 ;
        RECT -72.245 160.315 -71.915 160.645 ;
        RECT -72.245 158.955 -71.915 159.285 ;
        RECT -72.245 157.595 -71.915 157.925 ;
        RECT -72.245 156.235 -71.915 156.565 ;
        RECT -72.245 154.875 -71.915 155.205 ;
        RECT -72.245 153.515 -71.915 153.845 ;
        RECT -72.245 152.155 -71.915 152.485 ;
        RECT -72.245 150.795 -71.915 151.125 ;
        RECT -72.245 149.435 -71.915 149.765 ;
        RECT -72.245 148.075 -71.915 148.405 ;
        RECT -72.245 146.715 -71.915 147.045 ;
        RECT -72.245 145.355 -71.915 145.685 ;
        RECT -72.245 143.995 -71.915 144.325 ;
        RECT -72.245 142.635 -71.915 142.965 ;
        RECT -72.245 141.275 -71.915 141.605 ;
        RECT -72.245 139.915 -71.915 140.245 ;
        RECT -72.245 138.555 -71.915 138.885 ;
        RECT -72.245 137.195 -71.915 137.525 ;
        RECT -72.245 135.835 -71.915 136.165 ;
        RECT -72.245 134.475 -71.915 134.805 ;
        RECT -72.245 133.115 -71.915 133.445 ;
        RECT -72.245 131.755 -71.915 132.085 ;
        RECT -72.245 130.395 -71.915 130.725 ;
        RECT -72.245 129.035 -71.915 129.365 ;
        RECT -72.245 127.675 -71.915 128.005 ;
        RECT -72.245 126.315 -71.915 126.645 ;
        RECT -72.245 124.955 -71.915 125.285 ;
        RECT -72.245 123.595 -71.915 123.925 ;
        RECT -72.245 122.235 -71.915 122.565 ;
        RECT -72.245 120.875 -71.915 121.205 ;
        RECT -72.245 119.515 -71.915 119.845 ;
        RECT -72.245 118.155 -71.915 118.485 ;
        RECT -72.245 116.795 -71.915 117.125 ;
        RECT -72.245 115.435 -71.915 115.765 ;
        RECT -72.245 114.075 -71.915 114.405 ;
        RECT -72.245 112.715 -71.915 113.045 ;
        RECT -72.245 111.355 -71.915 111.685 ;
        RECT -72.245 109.995 -71.915 110.325 ;
        RECT -72.245 108.635 -71.915 108.965 ;
        RECT -72.245 107.275 -71.915 107.605 ;
        RECT -72.245 105.915 -71.915 106.245 ;
        RECT -72.245 104.555 -71.915 104.885 ;
        RECT -72.245 103.195 -71.915 103.525 ;
        RECT -72.245 101.835 -71.915 102.165 ;
        RECT -72.245 100.475 -71.915 100.805 ;
        RECT -72.245 99.115 -71.915 99.445 ;
        RECT -72.245 97.755 -71.915 98.085 ;
        RECT -72.245 96.395 -71.915 96.725 ;
        RECT -72.245 95.035 -71.915 95.365 ;
        RECT -72.245 93.675 -71.915 94.005 ;
        RECT -72.245 92.315 -71.915 92.645 ;
        RECT -72.245 90.955 -71.915 91.285 ;
        RECT -72.245 89.595 -71.915 89.925 ;
        RECT -72.245 88.235 -71.915 88.565 ;
        RECT -72.245 86.875 -71.915 87.205 ;
        RECT -72.245 85.515 -71.915 85.845 ;
        RECT -72.245 84.155 -71.915 84.485 ;
        RECT -72.245 82.795 -71.915 83.125 ;
        RECT -72.245 81.435 -71.915 81.765 ;
        RECT -72.245 80.075 -71.915 80.405 ;
        RECT -72.245 78.715 -71.915 79.045 ;
        RECT -72.245 77.355 -71.915 77.685 ;
        RECT -72.245 75.995 -71.915 76.325 ;
        RECT -72.245 74.635 -71.915 74.965 ;
        RECT -72.245 73.275 -71.915 73.605 ;
        RECT -72.245 71.915 -71.915 72.245 ;
        RECT -72.245 70.555 -71.915 70.885 ;
        RECT -72.245 69.195 -71.915 69.525 ;
        RECT -72.245 67.835 -71.915 68.165 ;
        RECT -72.245 66.475 -71.915 66.805 ;
        RECT -72.245 65.115 -71.915 65.445 ;
        RECT -72.245 63.755 -71.915 64.085 ;
        RECT -72.245 62.395 -71.915 62.725 ;
        RECT -72.245 61.035 -71.915 61.365 ;
        RECT -72.245 59.675 -71.915 60.005 ;
        RECT -72.245 58.315 -71.915 58.645 ;
        RECT -72.245 56.955 -71.915 57.285 ;
        RECT -72.245 55.595 -71.915 55.925 ;
        RECT -72.245 54.235 -71.915 54.565 ;
        RECT -72.245 52.875 -71.915 53.205 ;
        RECT -72.245 51.515 -71.915 51.845 ;
        RECT -72.245 50.155 -71.915 50.485 ;
        RECT -72.245 48.795 -71.915 49.125 ;
        RECT -72.245 47.435 -71.915 47.765 ;
        RECT -72.245 46.075 -71.915 46.405 ;
        RECT -72.245 44.715 -71.915 45.045 ;
        RECT -72.245 43.355 -71.915 43.685 ;
        RECT -72.245 41.995 -71.915 42.325 ;
        RECT -72.245 40.635 -71.915 40.965 ;
        RECT -72.245 39.275 -71.915 39.605 ;
        RECT -72.245 37.915 -71.915 38.245 ;
        RECT -72.245 36.555 -71.915 36.885 ;
        RECT -72.245 35.195 -71.915 35.525 ;
        RECT -72.245 33.835 -71.915 34.165 ;
        RECT -72.245 32.475 -71.915 32.805 ;
        RECT -72.245 31.115 -71.915 31.445 ;
        RECT -72.245 29.755 -71.915 30.085 ;
        RECT -72.245 28.395 -71.915 28.725 ;
        RECT -72.245 27.035 -71.915 27.365 ;
        RECT -72.245 25.675 -71.915 26.005 ;
        RECT -72.245 24.315 -71.915 24.645 ;
        RECT -72.245 22.955 -71.915 23.285 ;
        RECT -72.245 21.595 -71.915 21.925 ;
        RECT -72.245 20.235 -71.915 20.565 ;
        RECT -72.245 18.875 -71.915 19.205 ;
        RECT -72.245 17.515 -71.915 17.845 ;
        RECT -72.245 16.155 -71.915 16.485 ;
        RECT -72.245 14.795 -71.915 15.125 ;
        RECT -72.245 13.435 -71.915 13.765 ;
        RECT -72.245 12.075 -71.915 12.405 ;
        RECT -72.245 10.715 -71.915 11.045 ;
        RECT -72.245 9.355 -71.915 9.685 ;
        RECT -72.245 7.995 -71.915 8.325 ;
        RECT -72.245 6.635 -71.915 6.965 ;
        RECT -72.245 5.275 -71.915 5.605 ;
        RECT -72.245 3.915 -71.915 4.245 ;
        RECT -72.245 2.555 -71.915 2.885 ;
        RECT -72.245 1.195 -71.915 1.525 ;
        RECT -72.245 -0.165 -71.915 0.165 ;
        RECT -72.245 -1.525 -71.915 -1.195 ;
        RECT -72.245 -2.885 -71.915 -2.555 ;
        RECT -72.245 -4.245 -71.915 -3.915 ;
        RECT -72.245 -5.605 -71.915 -5.275 ;
        RECT -72.245 -6.965 -71.915 -6.635 ;
        RECT -72.245 -8.325 -71.915 -7.995 ;
        RECT -72.245 -9.685 -71.915 -9.355 ;
        RECT -72.245 -11.045 -71.915 -10.715 ;
        RECT -72.245 -12.405 -71.915 -12.075 ;
        RECT -72.245 -13.765 -71.915 -13.435 ;
        RECT -72.245 -15.125 -71.915 -14.795 ;
        RECT -72.245 -16.485 -71.915 -16.155 ;
        RECT -72.245 -17.845 -71.915 -17.515 ;
        RECT -72.245 -19.205 -71.915 -18.875 ;
        RECT -72.245 -20.565 -71.915 -20.235 ;
        RECT -72.245 -21.925 -71.915 -21.595 ;
        RECT -72.245 -23.285 -71.915 -22.955 ;
        RECT -72.245 -24.645 -71.915 -24.315 ;
        RECT -72.245 -26.005 -71.915 -25.675 ;
        RECT -72.245 -27.365 -71.915 -27.035 ;
        RECT -72.245 -28.725 -71.915 -28.395 ;
        RECT -72.245 -30.085 -71.915 -29.755 ;
        RECT -72.245 -31.445 -71.915 -31.115 ;
        RECT -72.245 -32.805 -71.915 -32.475 ;
        RECT -72.245 -34.165 -71.915 -33.835 ;
        RECT -72.245 -35.525 -71.915 -35.195 ;
        RECT -72.245 -36.885 -71.915 -36.555 ;
        RECT -72.245 -38.245 -71.915 -37.915 ;
        RECT -72.245 -39.605 -71.915 -39.275 ;
        RECT -72.245 -40.965 -71.915 -40.635 ;
        RECT -72.245 -42.325 -71.915 -41.995 ;
        RECT -72.245 -43.685 -71.915 -43.355 ;
        RECT -72.245 -45.045 -71.915 -44.715 ;
        RECT -72.245 -46.405 -71.915 -46.075 ;
        RECT -72.245 -47.765 -71.915 -47.435 ;
        RECT -72.245 -49.125 -71.915 -48.795 ;
        RECT -72.245 -50.485 -71.915 -50.155 ;
        RECT -72.245 -51.845 -71.915 -51.515 ;
        RECT -72.245 -53.205 -71.915 -52.875 ;
        RECT -72.245 -54.565 -71.915 -54.235 ;
        RECT -72.245 -55.925 -71.915 -55.595 ;
        RECT -72.245 -57.285 -71.915 -56.955 ;
        RECT -72.245 -58.645 -71.915 -58.315 ;
        RECT -72.245 -60.005 -71.915 -59.675 ;
        RECT -72.245 -61.365 -71.915 -61.035 ;
        RECT -72.245 -62.725 -71.915 -62.395 ;
        RECT -72.245 -64.085 -71.915 -63.755 ;
        RECT -72.245 -65.445 -71.915 -65.115 ;
        RECT -72.245 -66.805 -71.915 -66.475 ;
        RECT -72.245 -68.165 -71.915 -67.835 ;
        RECT -72.245 -69.525 -71.915 -69.195 ;
        RECT -72.245 -70.885 -71.915 -70.555 ;
        RECT -72.245 -72.245 -71.915 -71.915 ;
        RECT -72.245 -73.605 -71.915 -73.275 ;
        RECT -72.245 -74.965 -71.915 -74.635 ;
        RECT -72.245 -76.325 -71.915 -75.995 ;
        RECT -72.245 -77.685 -71.915 -77.355 ;
        RECT -72.245 -79.045 -71.915 -78.715 ;
        RECT -72.245 -80.405 -71.915 -80.075 ;
        RECT -72.245 -81.765 -71.915 -81.435 ;
        RECT -72.245 -83.125 -71.915 -82.795 ;
        RECT -72.245 -84.485 -71.915 -84.155 ;
        RECT -72.245 -85.845 -71.915 -85.515 ;
        RECT -72.245 -87.205 -71.915 -86.875 ;
        RECT -72.245 -88.565 -71.915 -88.235 ;
        RECT -72.245 -89.925 -71.915 -89.595 ;
        RECT -72.245 -91.285 -71.915 -90.955 ;
        RECT -72.245 -92.645 -71.915 -92.315 ;
        RECT -72.245 -94.005 -71.915 -93.675 ;
        RECT -72.245 -95.365 -71.915 -95.035 ;
        RECT -72.245 -96.725 -71.915 -96.395 ;
        RECT -72.245 -98.085 -71.915 -97.755 ;
        RECT -72.245 -99.445 -71.915 -99.115 ;
        RECT -72.245 -100.805 -71.915 -100.475 ;
        RECT -72.245 -102.165 -71.915 -101.835 ;
        RECT -72.245 -103.525 -71.915 -103.195 ;
        RECT -72.245 -104.885 -71.915 -104.555 ;
        RECT -72.245 -106.245 -71.915 -105.915 ;
        RECT -72.245 -107.605 -71.915 -107.275 ;
        RECT -72.245 -108.965 -71.915 -108.635 ;
        RECT -72.245 -110.325 -71.915 -109.995 ;
        RECT -72.245 -111.685 -71.915 -111.355 ;
        RECT -72.245 -113.045 -71.915 -112.715 ;
        RECT -72.245 -114.405 -71.915 -114.075 ;
        RECT -72.245 -115.765 -71.915 -115.435 ;
        RECT -72.245 -117.125 -71.915 -116.795 ;
        RECT -72.245 -118.485 -71.915 -118.155 ;
        RECT -72.245 -119.845 -71.915 -119.515 ;
        RECT -72.245 -121.205 -71.915 -120.875 ;
        RECT -72.245 -122.565 -71.915 -122.235 ;
        RECT -72.245 -123.925 -71.915 -123.595 ;
        RECT -72.245 -125.285 -71.915 -124.955 ;
        RECT -72.245 -126.645 -71.915 -126.315 ;
        RECT -72.245 -128.005 -71.915 -127.675 ;
        RECT -72.245 -129.365 -71.915 -129.035 ;
        RECT -72.245 -130.725 -71.915 -130.395 ;
        RECT -72.245 -132.085 -71.915 -131.755 ;
        RECT -72.245 -133.445 -71.915 -133.115 ;
        RECT -72.245 -134.805 -71.915 -134.475 ;
        RECT -72.245 -136.165 -71.915 -135.835 ;
        RECT -72.245 -137.525 -71.915 -137.195 ;
        RECT -72.245 -138.885 -71.915 -138.555 ;
        RECT -72.245 -140.245 -71.915 -139.915 ;
        RECT -72.245 -141.605 -71.915 -141.275 ;
        RECT -72.245 -142.965 -71.915 -142.635 ;
        RECT -72.245 -144.325 -71.915 -143.995 ;
        RECT -72.245 -145.685 -71.915 -145.355 ;
        RECT -72.245 -147.045 -71.915 -146.715 ;
        RECT -72.245 -148.405 -71.915 -148.075 ;
        RECT -72.245 -149.765 -71.915 -149.435 ;
        RECT -72.245 -151.125 -71.915 -150.795 ;
        RECT -72.245 -152.485 -71.915 -152.155 ;
        RECT -72.245 -153.845 -71.915 -153.515 ;
        RECT -72.245 -155.205 -71.915 -154.875 ;
        RECT -72.245 -156.565 -71.915 -156.235 ;
        RECT -72.245 -157.925 -71.915 -157.595 ;
        RECT -72.245 -159.285 -71.915 -158.955 ;
        RECT -72.245 -160.645 -71.915 -160.315 ;
        RECT -72.245 -162.005 -71.915 -161.675 ;
        RECT -72.245 -163.365 -71.915 -163.035 ;
        RECT -72.245 -164.725 -71.915 -164.395 ;
        RECT -72.245 -166.085 -71.915 -165.755 ;
        RECT -72.245 -167.445 -71.915 -167.115 ;
        RECT -72.245 -170.165 -71.915 -169.835 ;
        RECT -72.245 -171.525 -71.915 -171.195 ;
        RECT -72.245 -172.885 -71.915 -172.555 ;
        RECT -72.245 -174.245 -71.915 -173.915 ;
        RECT -72.245 -176.965 -71.915 -176.635 ;
        RECT -72.245 -178.325 -71.915 -177.995 ;
        RECT -72.245 -180.57 -71.915 -179.44 ;
        RECT -72.24 -180.685 -71.92 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -70.885 241.32 -70.555 242.45 ;
        RECT -70.885 239.195 -70.555 239.525 ;
        RECT -70.885 237.835 -70.555 238.165 ;
        RECT -70.885 236.475 -70.555 236.805 ;
        RECT -70.885 235.115 -70.555 235.445 ;
        RECT -70.885 233.755 -70.555 234.085 ;
        RECT -70.885 232.395 -70.555 232.725 ;
        RECT -70.885 231.035 -70.555 231.365 ;
        RECT -70.885 229.675 -70.555 230.005 ;
        RECT -70.885 228.315 -70.555 228.645 ;
        RECT -70.885 226.955 -70.555 227.285 ;
        RECT -70.885 225.595 -70.555 225.925 ;
        RECT -70.885 224.235 -70.555 224.565 ;
        RECT -70.885 222.875 -70.555 223.205 ;
        RECT -70.885 221.515 -70.555 221.845 ;
        RECT -70.885 220.155 -70.555 220.485 ;
        RECT -70.885 218.795 -70.555 219.125 ;
        RECT -70.885 217.435 -70.555 217.765 ;
        RECT -70.885 216.075 -70.555 216.405 ;
        RECT -70.885 214.715 -70.555 215.045 ;
        RECT -70.885 213.355 -70.555 213.685 ;
        RECT -70.885 211.995 -70.555 212.325 ;
        RECT -70.885 210.635 -70.555 210.965 ;
        RECT -70.885 209.275 -70.555 209.605 ;
        RECT -70.885 207.915 -70.555 208.245 ;
        RECT -70.885 206.555 -70.555 206.885 ;
        RECT -70.885 205.195 -70.555 205.525 ;
        RECT -70.885 203.835 -70.555 204.165 ;
        RECT -70.885 202.475 -70.555 202.805 ;
        RECT -70.885 201.115 -70.555 201.445 ;
        RECT -70.885 199.755 -70.555 200.085 ;
        RECT -70.885 198.395 -70.555 198.725 ;
        RECT -70.885 197.035 -70.555 197.365 ;
        RECT -70.885 195.675 -70.555 196.005 ;
        RECT -70.885 194.315 -70.555 194.645 ;
        RECT -70.885 192.955 -70.555 193.285 ;
        RECT -70.885 191.595 -70.555 191.925 ;
        RECT -70.885 190.235 -70.555 190.565 ;
        RECT -70.885 188.875 -70.555 189.205 ;
        RECT -70.885 187.515 -70.555 187.845 ;
        RECT -70.885 186.155 -70.555 186.485 ;
        RECT -70.885 184.795 -70.555 185.125 ;
        RECT -70.885 183.435 -70.555 183.765 ;
        RECT -70.885 182.075 -70.555 182.405 ;
        RECT -70.885 180.715 -70.555 181.045 ;
        RECT -70.885 179.355 -70.555 179.685 ;
        RECT -70.885 177.995 -70.555 178.325 ;
        RECT -70.885 176.635 -70.555 176.965 ;
        RECT -70.885 175.275 -70.555 175.605 ;
        RECT -70.885 173.915 -70.555 174.245 ;
        RECT -70.885 172.555 -70.555 172.885 ;
        RECT -70.885 171.195 -70.555 171.525 ;
        RECT -70.885 169.835 -70.555 170.165 ;
        RECT -70.885 168.475 -70.555 168.805 ;
        RECT -70.885 167.115 -70.555 167.445 ;
        RECT -70.885 165.755 -70.555 166.085 ;
        RECT -70.885 164.395 -70.555 164.725 ;
        RECT -70.885 163.035 -70.555 163.365 ;
        RECT -70.885 161.675 -70.555 162.005 ;
        RECT -70.885 160.315 -70.555 160.645 ;
        RECT -70.885 158.955 -70.555 159.285 ;
        RECT -70.885 157.595 -70.555 157.925 ;
        RECT -70.885 156.235 -70.555 156.565 ;
        RECT -70.885 154.875 -70.555 155.205 ;
        RECT -70.885 153.515 -70.555 153.845 ;
        RECT -70.885 152.155 -70.555 152.485 ;
        RECT -70.885 150.795 -70.555 151.125 ;
        RECT -70.885 149.435 -70.555 149.765 ;
        RECT -70.885 148.075 -70.555 148.405 ;
        RECT -70.885 146.715 -70.555 147.045 ;
        RECT -70.885 145.355 -70.555 145.685 ;
        RECT -70.885 143.995 -70.555 144.325 ;
        RECT -70.885 142.635 -70.555 142.965 ;
        RECT -70.885 141.275 -70.555 141.605 ;
        RECT -70.885 139.915 -70.555 140.245 ;
        RECT -70.885 138.555 -70.555 138.885 ;
        RECT -70.885 137.195 -70.555 137.525 ;
        RECT -70.885 135.835 -70.555 136.165 ;
        RECT -70.885 134.475 -70.555 134.805 ;
        RECT -70.885 133.115 -70.555 133.445 ;
        RECT -70.885 131.755 -70.555 132.085 ;
        RECT -70.885 130.395 -70.555 130.725 ;
        RECT -70.885 129.035 -70.555 129.365 ;
        RECT -70.885 127.675 -70.555 128.005 ;
        RECT -70.885 126.315 -70.555 126.645 ;
        RECT -70.885 124.955 -70.555 125.285 ;
        RECT -70.885 123.595 -70.555 123.925 ;
        RECT -70.885 122.235 -70.555 122.565 ;
        RECT -70.885 120.875 -70.555 121.205 ;
        RECT -70.885 119.515 -70.555 119.845 ;
        RECT -70.885 118.155 -70.555 118.485 ;
        RECT -70.885 116.795 -70.555 117.125 ;
        RECT -70.885 115.435 -70.555 115.765 ;
        RECT -70.885 114.075 -70.555 114.405 ;
        RECT -70.885 112.715 -70.555 113.045 ;
        RECT -70.885 111.355 -70.555 111.685 ;
        RECT -70.885 109.995 -70.555 110.325 ;
        RECT -70.885 108.635 -70.555 108.965 ;
        RECT -70.885 107.275 -70.555 107.605 ;
        RECT -70.885 105.915 -70.555 106.245 ;
        RECT -70.885 104.555 -70.555 104.885 ;
        RECT -70.885 103.195 -70.555 103.525 ;
        RECT -70.885 101.835 -70.555 102.165 ;
        RECT -70.885 100.475 -70.555 100.805 ;
        RECT -70.885 99.115 -70.555 99.445 ;
        RECT -70.885 97.755 -70.555 98.085 ;
        RECT -70.885 96.395 -70.555 96.725 ;
        RECT -70.885 95.035 -70.555 95.365 ;
        RECT -70.885 93.675 -70.555 94.005 ;
        RECT -70.885 92.315 -70.555 92.645 ;
        RECT -70.885 90.955 -70.555 91.285 ;
        RECT -70.885 89.595 -70.555 89.925 ;
        RECT -70.885 88.235 -70.555 88.565 ;
        RECT -70.885 86.875 -70.555 87.205 ;
        RECT -70.885 85.515 -70.555 85.845 ;
        RECT -70.885 84.155 -70.555 84.485 ;
        RECT -70.885 82.795 -70.555 83.125 ;
        RECT -70.885 81.435 -70.555 81.765 ;
        RECT -70.885 80.075 -70.555 80.405 ;
        RECT -70.885 78.715 -70.555 79.045 ;
        RECT -70.885 77.355 -70.555 77.685 ;
        RECT -70.885 75.995 -70.555 76.325 ;
        RECT -70.885 74.635 -70.555 74.965 ;
        RECT -70.885 73.275 -70.555 73.605 ;
        RECT -70.885 71.915 -70.555 72.245 ;
        RECT -70.885 70.555 -70.555 70.885 ;
        RECT -70.885 69.195 -70.555 69.525 ;
        RECT -70.885 67.835 -70.555 68.165 ;
        RECT -70.885 66.475 -70.555 66.805 ;
        RECT -70.885 65.115 -70.555 65.445 ;
        RECT -70.885 63.755 -70.555 64.085 ;
        RECT -70.885 62.395 -70.555 62.725 ;
        RECT -70.885 61.035 -70.555 61.365 ;
        RECT -70.885 59.675 -70.555 60.005 ;
        RECT -70.885 58.315 -70.555 58.645 ;
        RECT -70.885 56.955 -70.555 57.285 ;
        RECT -70.885 55.595 -70.555 55.925 ;
        RECT -70.885 54.235 -70.555 54.565 ;
        RECT -70.885 52.875 -70.555 53.205 ;
        RECT -70.885 51.515 -70.555 51.845 ;
        RECT -70.885 50.155 -70.555 50.485 ;
        RECT -70.885 48.795 -70.555 49.125 ;
        RECT -70.885 47.435 -70.555 47.765 ;
        RECT -70.885 46.075 -70.555 46.405 ;
        RECT -70.885 44.715 -70.555 45.045 ;
        RECT -70.885 43.355 -70.555 43.685 ;
        RECT -70.885 41.995 -70.555 42.325 ;
        RECT -70.885 40.635 -70.555 40.965 ;
        RECT -70.885 39.275 -70.555 39.605 ;
        RECT -70.885 37.915 -70.555 38.245 ;
        RECT -70.885 36.555 -70.555 36.885 ;
        RECT -70.885 35.195 -70.555 35.525 ;
        RECT -70.885 33.835 -70.555 34.165 ;
        RECT -70.885 32.475 -70.555 32.805 ;
        RECT -70.885 31.115 -70.555 31.445 ;
        RECT -70.885 29.755 -70.555 30.085 ;
        RECT -70.885 28.395 -70.555 28.725 ;
        RECT -70.885 27.035 -70.555 27.365 ;
        RECT -70.885 25.675 -70.555 26.005 ;
        RECT -70.885 24.315 -70.555 24.645 ;
        RECT -70.885 22.955 -70.555 23.285 ;
        RECT -70.885 21.595 -70.555 21.925 ;
        RECT -70.885 20.235 -70.555 20.565 ;
        RECT -70.885 18.875 -70.555 19.205 ;
        RECT -70.885 17.515 -70.555 17.845 ;
        RECT -70.885 16.155 -70.555 16.485 ;
        RECT -70.885 14.795 -70.555 15.125 ;
        RECT -70.885 13.435 -70.555 13.765 ;
        RECT -70.885 12.075 -70.555 12.405 ;
        RECT -70.885 10.715 -70.555 11.045 ;
        RECT -70.885 9.355 -70.555 9.685 ;
        RECT -70.885 7.995 -70.555 8.325 ;
        RECT -70.885 6.635 -70.555 6.965 ;
        RECT -70.885 5.275 -70.555 5.605 ;
        RECT -70.885 3.915 -70.555 4.245 ;
        RECT -70.885 2.555 -70.555 2.885 ;
        RECT -70.885 1.195 -70.555 1.525 ;
        RECT -70.885 -0.165 -70.555 0.165 ;
        RECT -70.885 -1.525 -70.555 -1.195 ;
        RECT -70.885 -2.885 -70.555 -2.555 ;
        RECT -70.885 -4.245 -70.555 -3.915 ;
        RECT -70.885 -5.605 -70.555 -5.275 ;
        RECT -70.885 -6.965 -70.555 -6.635 ;
        RECT -70.885 -8.325 -70.555 -7.995 ;
        RECT -70.885 -9.685 -70.555 -9.355 ;
        RECT -70.885 -11.045 -70.555 -10.715 ;
        RECT -70.885 -12.405 -70.555 -12.075 ;
        RECT -70.885 -13.765 -70.555 -13.435 ;
        RECT -70.885 -15.125 -70.555 -14.795 ;
        RECT -70.885 -16.485 -70.555 -16.155 ;
        RECT -70.885 -17.845 -70.555 -17.515 ;
        RECT -70.885 -19.205 -70.555 -18.875 ;
        RECT -70.885 -20.565 -70.555 -20.235 ;
        RECT -70.885 -21.925 -70.555 -21.595 ;
        RECT -70.885 -23.285 -70.555 -22.955 ;
        RECT -70.885 -24.645 -70.555 -24.315 ;
        RECT -70.885 -26.005 -70.555 -25.675 ;
        RECT -70.885 -27.365 -70.555 -27.035 ;
        RECT -70.885 -28.725 -70.555 -28.395 ;
        RECT -70.885 -30.085 -70.555 -29.755 ;
        RECT -70.885 -31.445 -70.555 -31.115 ;
        RECT -70.885 -32.805 -70.555 -32.475 ;
        RECT -70.885 -34.165 -70.555 -33.835 ;
        RECT -70.885 -35.525 -70.555 -35.195 ;
        RECT -70.885 -36.885 -70.555 -36.555 ;
        RECT -70.885 -38.245 -70.555 -37.915 ;
        RECT -70.885 -39.605 -70.555 -39.275 ;
        RECT -70.885 -40.965 -70.555 -40.635 ;
        RECT -70.885 -42.325 -70.555 -41.995 ;
        RECT -70.885 -43.685 -70.555 -43.355 ;
        RECT -70.885 -45.045 -70.555 -44.715 ;
        RECT -70.885 -46.405 -70.555 -46.075 ;
        RECT -70.885 -47.765 -70.555 -47.435 ;
        RECT -70.885 -49.125 -70.555 -48.795 ;
        RECT -70.885 -50.485 -70.555 -50.155 ;
        RECT -70.885 -51.845 -70.555 -51.515 ;
        RECT -70.885 -53.205 -70.555 -52.875 ;
        RECT -70.885 -54.565 -70.555 -54.235 ;
        RECT -70.885 -55.925 -70.555 -55.595 ;
        RECT -70.885 -57.285 -70.555 -56.955 ;
        RECT -70.885 -58.645 -70.555 -58.315 ;
        RECT -70.885 -60.005 -70.555 -59.675 ;
        RECT -70.885 -61.365 -70.555 -61.035 ;
        RECT -70.885 -62.725 -70.555 -62.395 ;
        RECT -70.885 -64.085 -70.555 -63.755 ;
        RECT -70.885 -65.445 -70.555 -65.115 ;
        RECT -70.885 -66.805 -70.555 -66.475 ;
        RECT -70.885 -68.165 -70.555 -67.835 ;
        RECT -70.885 -69.525 -70.555 -69.195 ;
        RECT -70.885 -70.885 -70.555 -70.555 ;
        RECT -70.885 -72.245 -70.555 -71.915 ;
        RECT -70.885 -73.605 -70.555 -73.275 ;
        RECT -70.885 -74.965 -70.555 -74.635 ;
        RECT -70.885 -76.325 -70.555 -75.995 ;
        RECT -70.885 -77.685 -70.555 -77.355 ;
        RECT -70.885 -79.045 -70.555 -78.715 ;
        RECT -70.885 -80.405 -70.555 -80.075 ;
        RECT -70.885 -81.765 -70.555 -81.435 ;
        RECT -70.885 -83.125 -70.555 -82.795 ;
        RECT -70.885 -84.485 -70.555 -84.155 ;
        RECT -70.885 -85.845 -70.555 -85.515 ;
        RECT -70.885 -87.205 -70.555 -86.875 ;
        RECT -70.885 -88.565 -70.555 -88.235 ;
        RECT -70.885 -89.925 -70.555 -89.595 ;
        RECT -70.885 -91.285 -70.555 -90.955 ;
        RECT -70.885 -92.645 -70.555 -92.315 ;
        RECT -70.885 -94.005 -70.555 -93.675 ;
        RECT -70.885 -95.365 -70.555 -95.035 ;
        RECT -70.885 -96.725 -70.555 -96.395 ;
        RECT -70.885 -98.085 -70.555 -97.755 ;
        RECT -70.885 -99.445 -70.555 -99.115 ;
        RECT -70.885 -100.805 -70.555 -100.475 ;
        RECT -70.885 -102.165 -70.555 -101.835 ;
        RECT -70.885 -103.525 -70.555 -103.195 ;
        RECT -70.885 -104.885 -70.555 -104.555 ;
        RECT -70.885 -106.245 -70.555 -105.915 ;
        RECT -70.885 -107.605 -70.555 -107.275 ;
        RECT -70.885 -108.965 -70.555 -108.635 ;
        RECT -70.885 -110.325 -70.555 -109.995 ;
        RECT -70.885 -111.685 -70.555 -111.355 ;
        RECT -70.885 -113.045 -70.555 -112.715 ;
        RECT -70.885 -114.405 -70.555 -114.075 ;
        RECT -70.885 -115.765 -70.555 -115.435 ;
        RECT -70.885 -117.125 -70.555 -116.795 ;
        RECT -70.885 -118.485 -70.555 -118.155 ;
        RECT -70.885 -119.845 -70.555 -119.515 ;
        RECT -70.885 -121.205 -70.555 -120.875 ;
        RECT -70.885 -122.565 -70.555 -122.235 ;
        RECT -70.885 -123.925 -70.555 -123.595 ;
        RECT -70.885 -125.285 -70.555 -124.955 ;
        RECT -70.885 -126.645 -70.555 -126.315 ;
        RECT -70.885 -128.005 -70.555 -127.675 ;
        RECT -70.885 -129.365 -70.555 -129.035 ;
        RECT -70.885 -130.725 -70.555 -130.395 ;
        RECT -70.885 -132.085 -70.555 -131.755 ;
        RECT -70.885 -133.445 -70.555 -133.115 ;
        RECT -70.885 -134.805 -70.555 -134.475 ;
        RECT -70.885 -136.165 -70.555 -135.835 ;
        RECT -70.885 -137.525 -70.555 -137.195 ;
        RECT -70.885 -138.885 -70.555 -138.555 ;
        RECT -70.885 -140.245 -70.555 -139.915 ;
        RECT -70.885 -141.605 -70.555 -141.275 ;
        RECT -70.885 -142.965 -70.555 -142.635 ;
        RECT -70.885 -144.325 -70.555 -143.995 ;
        RECT -70.885 -145.685 -70.555 -145.355 ;
        RECT -70.885 -147.045 -70.555 -146.715 ;
        RECT -70.885 -148.405 -70.555 -148.075 ;
        RECT -70.885 -149.765 -70.555 -149.435 ;
        RECT -70.885 -151.125 -70.555 -150.795 ;
        RECT -70.885 -152.485 -70.555 -152.155 ;
        RECT -70.885 -153.845 -70.555 -153.515 ;
        RECT -70.885 -155.205 -70.555 -154.875 ;
        RECT -70.885 -156.565 -70.555 -156.235 ;
        RECT -70.885 -157.925 -70.555 -157.595 ;
        RECT -70.885 -159.285 -70.555 -158.955 ;
        RECT -70.885 -160.645 -70.555 -160.315 ;
        RECT -70.885 -162.005 -70.555 -161.675 ;
        RECT -70.885 -163.365 -70.555 -163.035 ;
        RECT -70.885 -164.725 -70.555 -164.395 ;
        RECT -70.885 -166.085 -70.555 -165.755 ;
        RECT -70.885 -167.445 -70.555 -167.115 ;
        RECT -70.885 -170.165 -70.555 -169.835 ;
        RECT -70.885 -171.525 -70.555 -171.195 ;
        RECT -70.88 -172.2 -70.56 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -69.525 -102.165 -69.195 -101.835 ;
        RECT -69.525 -103.525 -69.195 -103.195 ;
        RECT -69.525 -104.885 -69.195 -104.555 ;
        RECT -69.525 -106.245 -69.195 -105.915 ;
        RECT -69.525 -107.605 -69.195 -107.275 ;
        RECT -69.525 -108.965 -69.195 -108.635 ;
        RECT -69.525 -110.325 -69.195 -109.995 ;
        RECT -69.525 -111.685 -69.195 -111.355 ;
        RECT -69.525 -113.045 -69.195 -112.715 ;
        RECT -69.525 -114.405 -69.195 -114.075 ;
        RECT -69.525 -115.765 -69.195 -115.435 ;
        RECT -69.525 -117.125 -69.195 -116.795 ;
        RECT -69.525 -118.485 -69.195 -118.155 ;
        RECT -69.525 -119.845 -69.195 -119.515 ;
        RECT -69.525 -121.205 -69.195 -120.875 ;
        RECT -69.525 -122.565 -69.195 -122.235 ;
        RECT -69.525 -123.925 -69.195 -123.595 ;
        RECT -69.525 -125.285 -69.195 -124.955 ;
        RECT -69.525 -126.645 -69.195 -126.315 ;
        RECT -69.525 -128.005 -69.195 -127.675 ;
        RECT -69.525 -129.365 -69.195 -129.035 ;
        RECT -69.525 -130.725 -69.195 -130.395 ;
        RECT -69.525 -132.085 -69.195 -131.755 ;
        RECT -69.525 -133.445 -69.195 -133.115 ;
        RECT -69.525 -134.805 -69.195 -134.475 ;
        RECT -69.525 -136.165 -69.195 -135.835 ;
        RECT -69.525 -137.525 -69.195 -137.195 ;
        RECT -69.525 -138.885 -69.195 -138.555 ;
        RECT -69.525 -140.245 -69.195 -139.915 ;
        RECT -69.525 -141.605 -69.195 -141.275 ;
        RECT -69.525 -142.965 -69.195 -142.635 ;
        RECT -69.525 -144.325 -69.195 -143.995 ;
        RECT -69.525 -145.685 -69.195 -145.355 ;
        RECT -69.525 -147.045 -69.195 -146.715 ;
        RECT -69.525 -148.405 -69.195 -148.075 ;
        RECT -69.525 -149.765 -69.195 -149.435 ;
        RECT -69.525 -151.125 -69.195 -150.795 ;
        RECT -69.525 -152.485 -69.195 -152.155 ;
        RECT -69.525 -153.845 -69.195 -153.515 ;
        RECT -69.525 -155.205 -69.195 -154.875 ;
        RECT -69.525 -156.565 -69.195 -156.235 ;
        RECT -69.525 -157.925 -69.195 -157.595 ;
        RECT -69.525 -159.285 -69.195 -158.955 ;
        RECT -69.525 -160.645 -69.195 -160.315 ;
        RECT -69.525 -162.005 -69.195 -161.675 ;
        RECT -69.525 -163.365 -69.195 -163.035 ;
        RECT -69.525 -164.725 -69.195 -164.395 ;
        RECT -69.525 -166.085 -69.195 -165.755 ;
        RECT -69.525 -167.445 -69.195 -167.115 ;
        RECT -69.525 -170.165 -69.195 -169.835 ;
        RECT -69.525 -172.885 -69.195 -172.555 ;
        RECT -69.525 -174.245 -69.195 -173.915 ;
        RECT -69.525 -175.725 -69.195 -175.395 ;
        RECT -69.525 -176.965 -69.195 -176.635 ;
        RECT -69.525 -178.325 -69.195 -177.995 ;
        RECT -69.525 -180.57 -69.195 -179.44 ;
        RECT -69.52 -180.685 -69.2 242.565 ;
        RECT -69.525 241.32 -69.195 242.45 ;
        RECT -69.525 239.195 -69.195 239.525 ;
        RECT -69.525 237.835 -69.195 238.165 ;
        RECT -69.525 236.475 -69.195 236.805 ;
        RECT -69.525 235.115 -69.195 235.445 ;
        RECT -69.525 233.755 -69.195 234.085 ;
        RECT -69.525 232.395 -69.195 232.725 ;
        RECT -69.525 231.035 -69.195 231.365 ;
        RECT -69.525 229.675 -69.195 230.005 ;
        RECT -69.525 228.315 -69.195 228.645 ;
        RECT -69.525 226.955 -69.195 227.285 ;
        RECT -69.525 225.595 -69.195 225.925 ;
        RECT -69.525 224.235 -69.195 224.565 ;
        RECT -69.525 222.875 -69.195 223.205 ;
        RECT -69.525 221.515 -69.195 221.845 ;
        RECT -69.525 220.155 -69.195 220.485 ;
        RECT -69.525 218.795 -69.195 219.125 ;
        RECT -69.525 217.435 -69.195 217.765 ;
        RECT -69.525 216.075 -69.195 216.405 ;
        RECT -69.525 214.715 -69.195 215.045 ;
        RECT -69.525 213.355 -69.195 213.685 ;
        RECT -69.525 211.995 -69.195 212.325 ;
        RECT -69.525 210.635 -69.195 210.965 ;
        RECT -69.525 209.275 -69.195 209.605 ;
        RECT -69.525 207.915 -69.195 208.245 ;
        RECT -69.525 206.555 -69.195 206.885 ;
        RECT -69.525 205.195 -69.195 205.525 ;
        RECT -69.525 203.835 -69.195 204.165 ;
        RECT -69.525 202.475 -69.195 202.805 ;
        RECT -69.525 201.115 -69.195 201.445 ;
        RECT -69.525 199.755 -69.195 200.085 ;
        RECT -69.525 198.395 -69.195 198.725 ;
        RECT -69.525 197.035 -69.195 197.365 ;
        RECT -69.525 195.675 -69.195 196.005 ;
        RECT -69.525 194.315 -69.195 194.645 ;
        RECT -69.525 192.955 -69.195 193.285 ;
        RECT -69.525 191.595 -69.195 191.925 ;
        RECT -69.525 190.235 -69.195 190.565 ;
        RECT -69.525 188.875 -69.195 189.205 ;
        RECT -69.525 187.515 -69.195 187.845 ;
        RECT -69.525 186.155 -69.195 186.485 ;
        RECT -69.525 184.795 -69.195 185.125 ;
        RECT -69.525 183.435 -69.195 183.765 ;
        RECT -69.525 182.075 -69.195 182.405 ;
        RECT -69.525 180.715 -69.195 181.045 ;
        RECT -69.525 179.355 -69.195 179.685 ;
        RECT -69.525 177.995 -69.195 178.325 ;
        RECT -69.525 176.635 -69.195 176.965 ;
        RECT -69.525 175.275 -69.195 175.605 ;
        RECT -69.525 173.915 -69.195 174.245 ;
        RECT -69.525 172.555 -69.195 172.885 ;
        RECT -69.525 171.195 -69.195 171.525 ;
        RECT -69.525 169.835 -69.195 170.165 ;
        RECT -69.525 168.475 -69.195 168.805 ;
        RECT -69.525 167.115 -69.195 167.445 ;
        RECT -69.525 165.755 -69.195 166.085 ;
        RECT -69.525 164.395 -69.195 164.725 ;
        RECT -69.525 163.035 -69.195 163.365 ;
        RECT -69.525 161.675 -69.195 162.005 ;
        RECT -69.525 160.315 -69.195 160.645 ;
        RECT -69.525 158.955 -69.195 159.285 ;
        RECT -69.525 157.595 -69.195 157.925 ;
        RECT -69.525 156.235 -69.195 156.565 ;
        RECT -69.525 154.875 -69.195 155.205 ;
        RECT -69.525 153.515 -69.195 153.845 ;
        RECT -69.525 152.155 -69.195 152.485 ;
        RECT -69.525 150.795 -69.195 151.125 ;
        RECT -69.525 149.435 -69.195 149.765 ;
        RECT -69.525 148.075 -69.195 148.405 ;
        RECT -69.525 146.715 -69.195 147.045 ;
        RECT -69.525 145.355 -69.195 145.685 ;
        RECT -69.525 143.995 -69.195 144.325 ;
        RECT -69.525 142.635 -69.195 142.965 ;
        RECT -69.525 141.275 -69.195 141.605 ;
        RECT -69.525 139.915 -69.195 140.245 ;
        RECT -69.525 138.555 -69.195 138.885 ;
        RECT -69.525 137.195 -69.195 137.525 ;
        RECT -69.525 135.835 -69.195 136.165 ;
        RECT -69.525 134.475 -69.195 134.805 ;
        RECT -69.525 133.115 -69.195 133.445 ;
        RECT -69.525 131.755 -69.195 132.085 ;
        RECT -69.525 130.395 -69.195 130.725 ;
        RECT -69.525 129.035 -69.195 129.365 ;
        RECT -69.525 127.675 -69.195 128.005 ;
        RECT -69.525 126.315 -69.195 126.645 ;
        RECT -69.525 124.955 -69.195 125.285 ;
        RECT -69.525 123.595 -69.195 123.925 ;
        RECT -69.525 122.235 -69.195 122.565 ;
        RECT -69.525 120.875 -69.195 121.205 ;
        RECT -69.525 119.515 -69.195 119.845 ;
        RECT -69.525 118.155 -69.195 118.485 ;
        RECT -69.525 116.795 -69.195 117.125 ;
        RECT -69.525 115.435 -69.195 115.765 ;
        RECT -69.525 114.075 -69.195 114.405 ;
        RECT -69.525 112.715 -69.195 113.045 ;
        RECT -69.525 111.355 -69.195 111.685 ;
        RECT -69.525 109.995 -69.195 110.325 ;
        RECT -69.525 108.635 -69.195 108.965 ;
        RECT -69.525 107.275 -69.195 107.605 ;
        RECT -69.525 105.915 -69.195 106.245 ;
        RECT -69.525 104.555 -69.195 104.885 ;
        RECT -69.525 103.195 -69.195 103.525 ;
        RECT -69.525 101.835 -69.195 102.165 ;
        RECT -69.525 100.475 -69.195 100.805 ;
        RECT -69.525 99.115 -69.195 99.445 ;
        RECT -69.525 97.755 -69.195 98.085 ;
        RECT -69.525 96.395 -69.195 96.725 ;
        RECT -69.525 95.035 -69.195 95.365 ;
        RECT -69.525 93.675 -69.195 94.005 ;
        RECT -69.525 92.315 -69.195 92.645 ;
        RECT -69.525 90.955 -69.195 91.285 ;
        RECT -69.525 89.595 -69.195 89.925 ;
        RECT -69.525 88.235 -69.195 88.565 ;
        RECT -69.525 86.875 -69.195 87.205 ;
        RECT -69.525 85.515 -69.195 85.845 ;
        RECT -69.525 84.155 -69.195 84.485 ;
        RECT -69.525 82.795 -69.195 83.125 ;
        RECT -69.525 81.435 -69.195 81.765 ;
        RECT -69.525 80.075 -69.195 80.405 ;
        RECT -69.525 78.715 -69.195 79.045 ;
        RECT -69.525 77.355 -69.195 77.685 ;
        RECT -69.525 75.995 -69.195 76.325 ;
        RECT -69.525 74.635 -69.195 74.965 ;
        RECT -69.525 73.275 -69.195 73.605 ;
        RECT -69.525 71.915 -69.195 72.245 ;
        RECT -69.525 70.555 -69.195 70.885 ;
        RECT -69.525 69.195 -69.195 69.525 ;
        RECT -69.525 67.835 -69.195 68.165 ;
        RECT -69.525 66.475 -69.195 66.805 ;
        RECT -69.525 65.115 -69.195 65.445 ;
        RECT -69.525 63.755 -69.195 64.085 ;
        RECT -69.525 62.395 -69.195 62.725 ;
        RECT -69.525 61.035 -69.195 61.365 ;
        RECT -69.525 59.675 -69.195 60.005 ;
        RECT -69.525 58.315 -69.195 58.645 ;
        RECT -69.525 56.955 -69.195 57.285 ;
        RECT -69.525 55.595 -69.195 55.925 ;
        RECT -69.525 54.235 -69.195 54.565 ;
        RECT -69.525 52.875 -69.195 53.205 ;
        RECT -69.525 51.515 -69.195 51.845 ;
        RECT -69.525 50.155 -69.195 50.485 ;
        RECT -69.525 48.795 -69.195 49.125 ;
        RECT -69.525 47.435 -69.195 47.765 ;
        RECT -69.525 46.075 -69.195 46.405 ;
        RECT -69.525 44.715 -69.195 45.045 ;
        RECT -69.525 43.355 -69.195 43.685 ;
        RECT -69.525 41.995 -69.195 42.325 ;
        RECT -69.525 40.635 -69.195 40.965 ;
        RECT -69.525 39.275 -69.195 39.605 ;
        RECT -69.525 37.915 -69.195 38.245 ;
        RECT -69.525 36.555 -69.195 36.885 ;
        RECT -69.525 35.195 -69.195 35.525 ;
        RECT -69.525 33.835 -69.195 34.165 ;
        RECT -69.525 32.475 -69.195 32.805 ;
        RECT -69.525 31.115 -69.195 31.445 ;
        RECT -69.525 29.755 -69.195 30.085 ;
        RECT -69.525 28.395 -69.195 28.725 ;
        RECT -69.525 27.035 -69.195 27.365 ;
        RECT -69.525 25.675 -69.195 26.005 ;
        RECT -69.525 24.315 -69.195 24.645 ;
        RECT -69.525 22.955 -69.195 23.285 ;
        RECT -69.525 21.595 -69.195 21.925 ;
        RECT -69.525 20.235 -69.195 20.565 ;
        RECT -69.525 18.875 -69.195 19.205 ;
        RECT -69.525 17.515 -69.195 17.845 ;
        RECT -69.525 16.155 -69.195 16.485 ;
        RECT -69.525 14.795 -69.195 15.125 ;
        RECT -69.525 13.435 -69.195 13.765 ;
        RECT -69.525 12.075 -69.195 12.405 ;
        RECT -69.525 10.715 -69.195 11.045 ;
        RECT -69.525 9.355 -69.195 9.685 ;
        RECT -69.525 7.995 -69.195 8.325 ;
        RECT -69.525 6.635 -69.195 6.965 ;
        RECT -69.525 5.275 -69.195 5.605 ;
        RECT -69.525 3.915 -69.195 4.245 ;
        RECT -69.525 2.555 -69.195 2.885 ;
        RECT -69.525 1.195 -69.195 1.525 ;
        RECT -69.525 -0.165 -69.195 0.165 ;
        RECT -69.525 -1.525 -69.195 -1.195 ;
        RECT -69.525 -2.885 -69.195 -2.555 ;
        RECT -69.525 -4.245 -69.195 -3.915 ;
        RECT -69.525 -5.605 -69.195 -5.275 ;
        RECT -69.525 -6.965 -69.195 -6.635 ;
        RECT -69.525 -8.325 -69.195 -7.995 ;
        RECT -69.525 -9.685 -69.195 -9.355 ;
        RECT -69.525 -11.045 -69.195 -10.715 ;
        RECT -69.525 -12.405 -69.195 -12.075 ;
        RECT -69.525 -13.765 -69.195 -13.435 ;
        RECT -69.525 -15.125 -69.195 -14.795 ;
        RECT -69.525 -16.485 -69.195 -16.155 ;
        RECT -69.525 -17.845 -69.195 -17.515 ;
        RECT -69.525 -19.205 -69.195 -18.875 ;
        RECT -69.525 -20.565 -69.195 -20.235 ;
        RECT -69.525 -21.925 -69.195 -21.595 ;
        RECT -69.525 -23.285 -69.195 -22.955 ;
        RECT -69.525 -24.645 -69.195 -24.315 ;
        RECT -69.525 -26.005 -69.195 -25.675 ;
        RECT -69.525 -27.365 -69.195 -27.035 ;
        RECT -69.525 -28.725 -69.195 -28.395 ;
        RECT -69.525 -30.085 -69.195 -29.755 ;
        RECT -69.525 -31.445 -69.195 -31.115 ;
        RECT -69.525 -32.805 -69.195 -32.475 ;
        RECT -69.525 -34.165 -69.195 -33.835 ;
        RECT -69.525 -35.525 -69.195 -35.195 ;
        RECT -69.525 -36.885 -69.195 -36.555 ;
        RECT -69.525 -38.245 -69.195 -37.915 ;
        RECT -69.525 -39.605 -69.195 -39.275 ;
        RECT -69.525 -40.965 -69.195 -40.635 ;
        RECT -69.525 -42.325 -69.195 -41.995 ;
        RECT -69.525 -43.685 -69.195 -43.355 ;
        RECT -69.525 -45.045 -69.195 -44.715 ;
        RECT -69.525 -46.405 -69.195 -46.075 ;
        RECT -69.525 -47.765 -69.195 -47.435 ;
        RECT -69.525 -49.125 -69.195 -48.795 ;
        RECT -69.525 -50.485 -69.195 -50.155 ;
        RECT -69.525 -51.845 -69.195 -51.515 ;
        RECT -69.525 -53.205 -69.195 -52.875 ;
        RECT -69.525 -54.565 -69.195 -54.235 ;
        RECT -69.525 -55.925 -69.195 -55.595 ;
        RECT -69.525 -57.285 -69.195 -56.955 ;
        RECT -69.525 -58.645 -69.195 -58.315 ;
        RECT -69.525 -60.005 -69.195 -59.675 ;
        RECT -69.525 -61.365 -69.195 -61.035 ;
        RECT -69.525 -62.725 -69.195 -62.395 ;
        RECT -69.525 -64.085 -69.195 -63.755 ;
        RECT -69.525 -65.445 -69.195 -65.115 ;
        RECT -69.525 -66.805 -69.195 -66.475 ;
        RECT -69.525 -68.165 -69.195 -67.835 ;
        RECT -69.525 -69.525 -69.195 -69.195 ;
        RECT -69.525 -70.885 -69.195 -70.555 ;
        RECT -69.525 -72.245 -69.195 -71.915 ;
        RECT -69.525 -73.605 -69.195 -73.275 ;
        RECT -69.525 -74.965 -69.195 -74.635 ;
        RECT -69.525 -76.325 -69.195 -75.995 ;
        RECT -69.525 -77.685 -69.195 -77.355 ;
        RECT -69.525 -79.045 -69.195 -78.715 ;
        RECT -69.525 -80.405 -69.195 -80.075 ;
        RECT -69.525 -81.765 -69.195 -81.435 ;
        RECT -69.525 -83.125 -69.195 -82.795 ;
        RECT -69.525 -84.485 -69.195 -84.155 ;
        RECT -69.525 -85.845 -69.195 -85.515 ;
        RECT -69.525 -87.205 -69.195 -86.875 ;
        RECT -69.525 -88.565 -69.195 -88.235 ;
        RECT -69.525 -89.925 -69.195 -89.595 ;
        RECT -69.525 -91.285 -69.195 -90.955 ;
        RECT -69.525 -92.645 -69.195 -92.315 ;
        RECT -69.525 -94.005 -69.195 -93.675 ;
        RECT -69.525 -95.365 -69.195 -95.035 ;
        RECT -69.525 -96.725 -69.195 -96.395 ;
        RECT -69.525 -98.085 -69.195 -97.755 ;
        RECT -69.525 -99.445 -69.195 -99.115 ;
        RECT -69.525 -100.805 -69.195 -100.475 ;
    END
    PORT
      LAYER met3 ;
        RECT -74.965 214.715 -74.635 215.045 ;
        RECT -74.965 213.355 -74.635 213.685 ;
        RECT -74.965 211.995 -74.635 212.325 ;
        RECT -74.965 210.635 -74.635 210.965 ;
        RECT -74.965 209.275 -74.635 209.605 ;
        RECT -74.965 207.915 -74.635 208.245 ;
        RECT -74.965 206.555 -74.635 206.885 ;
        RECT -74.965 205.195 -74.635 205.525 ;
        RECT -74.965 203.835 -74.635 204.165 ;
        RECT -74.965 202.475 -74.635 202.805 ;
        RECT -74.965 201.115 -74.635 201.445 ;
        RECT -74.965 199.755 -74.635 200.085 ;
        RECT -74.965 198.395 -74.635 198.725 ;
        RECT -74.965 197.035 -74.635 197.365 ;
        RECT -74.965 195.675 -74.635 196.005 ;
        RECT -74.965 194.315 -74.635 194.645 ;
        RECT -74.965 192.955 -74.635 193.285 ;
        RECT -74.965 191.595 -74.635 191.925 ;
        RECT -74.965 190.235 -74.635 190.565 ;
        RECT -74.965 188.875 -74.635 189.205 ;
        RECT -74.965 187.515 -74.635 187.845 ;
        RECT -74.965 186.155 -74.635 186.485 ;
        RECT -74.965 184.795 -74.635 185.125 ;
        RECT -74.965 183.435 -74.635 183.765 ;
        RECT -74.965 182.075 -74.635 182.405 ;
        RECT -74.965 180.715 -74.635 181.045 ;
        RECT -74.965 179.355 -74.635 179.685 ;
        RECT -74.965 177.995 -74.635 178.325 ;
        RECT -74.965 176.635 -74.635 176.965 ;
        RECT -74.965 175.275 -74.635 175.605 ;
        RECT -74.965 173.915 -74.635 174.245 ;
        RECT -74.965 172.555 -74.635 172.885 ;
        RECT -74.965 171.195 -74.635 171.525 ;
        RECT -74.965 169.835 -74.635 170.165 ;
        RECT -74.965 168.475 -74.635 168.805 ;
        RECT -74.965 167.115 -74.635 167.445 ;
        RECT -74.965 165.755 -74.635 166.085 ;
        RECT -74.965 164.395 -74.635 164.725 ;
        RECT -74.965 163.035 -74.635 163.365 ;
        RECT -74.965 161.675 -74.635 162.005 ;
        RECT -74.965 160.315 -74.635 160.645 ;
        RECT -74.965 158.955 -74.635 159.285 ;
        RECT -74.965 157.595 -74.635 157.925 ;
        RECT -74.965 156.235 -74.635 156.565 ;
        RECT -74.965 154.875 -74.635 155.205 ;
        RECT -74.965 153.515 -74.635 153.845 ;
        RECT -74.965 152.155 -74.635 152.485 ;
        RECT -74.965 150.795 -74.635 151.125 ;
        RECT -74.965 149.435 -74.635 149.765 ;
        RECT -74.965 148.075 -74.635 148.405 ;
        RECT -74.965 146.715 -74.635 147.045 ;
        RECT -74.965 145.355 -74.635 145.685 ;
        RECT -74.965 143.995 -74.635 144.325 ;
        RECT -74.965 142.635 -74.635 142.965 ;
        RECT -74.965 141.275 -74.635 141.605 ;
        RECT -74.965 139.915 -74.635 140.245 ;
        RECT -74.965 138.555 -74.635 138.885 ;
        RECT -74.965 137.195 -74.635 137.525 ;
        RECT -74.965 135.835 -74.635 136.165 ;
        RECT -74.965 134.475 -74.635 134.805 ;
        RECT -74.965 133.115 -74.635 133.445 ;
        RECT -74.965 131.755 -74.635 132.085 ;
        RECT -74.965 130.395 -74.635 130.725 ;
        RECT -74.965 129.035 -74.635 129.365 ;
        RECT -74.965 127.675 -74.635 128.005 ;
        RECT -74.965 126.315 -74.635 126.645 ;
        RECT -74.965 124.955 -74.635 125.285 ;
        RECT -74.965 123.595 -74.635 123.925 ;
        RECT -74.965 122.235 -74.635 122.565 ;
        RECT -74.965 120.875 -74.635 121.205 ;
        RECT -74.965 119.515 -74.635 119.845 ;
        RECT -74.965 118.155 -74.635 118.485 ;
        RECT -74.965 116.795 -74.635 117.125 ;
        RECT -74.965 115.435 -74.635 115.765 ;
        RECT -74.965 114.075 -74.635 114.405 ;
        RECT -74.965 112.715 -74.635 113.045 ;
        RECT -74.965 111.355 -74.635 111.685 ;
        RECT -74.965 109.995 -74.635 110.325 ;
        RECT -74.965 108.635 -74.635 108.965 ;
        RECT -74.965 107.275 -74.635 107.605 ;
        RECT -74.965 105.915 -74.635 106.245 ;
        RECT -74.965 104.555 -74.635 104.885 ;
        RECT -74.965 103.195 -74.635 103.525 ;
        RECT -74.965 101.835 -74.635 102.165 ;
        RECT -74.965 100.475 -74.635 100.805 ;
        RECT -74.965 99.115 -74.635 99.445 ;
        RECT -74.965 97.755 -74.635 98.085 ;
        RECT -74.965 96.395 -74.635 96.725 ;
        RECT -74.965 95.035 -74.635 95.365 ;
        RECT -74.965 93.675 -74.635 94.005 ;
        RECT -74.965 92.315 -74.635 92.645 ;
        RECT -74.965 90.955 -74.635 91.285 ;
        RECT -74.965 89.595 -74.635 89.925 ;
        RECT -74.965 88.235 -74.635 88.565 ;
        RECT -74.965 86.875 -74.635 87.205 ;
        RECT -74.965 85.515 -74.635 85.845 ;
        RECT -74.965 84.155 -74.635 84.485 ;
        RECT -74.965 82.795 -74.635 83.125 ;
        RECT -74.965 81.435 -74.635 81.765 ;
        RECT -74.965 80.075 -74.635 80.405 ;
        RECT -74.965 78.715 -74.635 79.045 ;
        RECT -74.965 77.355 -74.635 77.685 ;
        RECT -74.965 75.995 -74.635 76.325 ;
        RECT -74.965 74.635 -74.635 74.965 ;
        RECT -74.965 73.275 -74.635 73.605 ;
        RECT -74.965 71.915 -74.635 72.245 ;
        RECT -74.965 70.555 -74.635 70.885 ;
        RECT -74.965 69.195 -74.635 69.525 ;
        RECT -74.965 67.835 -74.635 68.165 ;
        RECT -74.965 66.475 -74.635 66.805 ;
        RECT -74.965 65.115 -74.635 65.445 ;
        RECT -74.965 63.755 -74.635 64.085 ;
        RECT -74.965 62.395 -74.635 62.725 ;
        RECT -74.965 61.035 -74.635 61.365 ;
        RECT -74.965 59.675 -74.635 60.005 ;
        RECT -74.965 58.315 -74.635 58.645 ;
        RECT -74.965 56.955 -74.635 57.285 ;
        RECT -74.965 55.595 -74.635 55.925 ;
        RECT -74.965 54.235 -74.635 54.565 ;
        RECT -74.965 52.875 -74.635 53.205 ;
        RECT -74.965 51.515 -74.635 51.845 ;
        RECT -74.965 50.155 -74.635 50.485 ;
        RECT -74.965 48.795 -74.635 49.125 ;
        RECT -74.965 47.435 -74.635 47.765 ;
        RECT -74.965 46.075 -74.635 46.405 ;
        RECT -74.965 44.715 -74.635 45.045 ;
        RECT -74.965 43.355 -74.635 43.685 ;
        RECT -74.965 41.995 -74.635 42.325 ;
        RECT -74.965 40.635 -74.635 40.965 ;
        RECT -74.965 39.275 -74.635 39.605 ;
        RECT -74.965 37.915 -74.635 38.245 ;
        RECT -74.965 36.555 -74.635 36.885 ;
        RECT -74.965 35.195 -74.635 35.525 ;
        RECT -74.965 33.835 -74.635 34.165 ;
        RECT -74.965 32.475 -74.635 32.805 ;
        RECT -74.965 31.115 -74.635 31.445 ;
        RECT -74.965 29.755 -74.635 30.085 ;
        RECT -74.965 28.395 -74.635 28.725 ;
        RECT -74.965 27.035 -74.635 27.365 ;
        RECT -74.965 25.675 -74.635 26.005 ;
        RECT -74.965 24.315 -74.635 24.645 ;
        RECT -74.965 22.955 -74.635 23.285 ;
        RECT -74.965 21.595 -74.635 21.925 ;
        RECT -74.965 20.235 -74.635 20.565 ;
        RECT -74.965 18.875 -74.635 19.205 ;
        RECT -74.965 17.515 -74.635 17.845 ;
        RECT -74.965 16.155 -74.635 16.485 ;
        RECT -74.965 14.795 -74.635 15.125 ;
        RECT -74.965 13.435 -74.635 13.765 ;
        RECT -74.965 12.075 -74.635 12.405 ;
        RECT -74.965 10.715 -74.635 11.045 ;
        RECT -74.965 9.355 -74.635 9.685 ;
        RECT -74.965 7.995 -74.635 8.325 ;
        RECT -74.965 6.635 -74.635 6.965 ;
        RECT -74.965 5.275 -74.635 5.605 ;
        RECT -74.965 3.915 -74.635 4.245 ;
        RECT -74.965 2.555 -74.635 2.885 ;
        RECT -74.965 1.195 -74.635 1.525 ;
        RECT -74.965 -0.165 -74.635 0.165 ;
        RECT -74.965 -1.525 -74.635 -1.195 ;
        RECT -74.965 -2.885 -74.635 -2.555 ;
        RECT -74.965 -4.245 -74.635 -3.915 ;
        RECT -74.965 -5.605 -74.635 -5.275 ;
        RECT -74.965 -6.965 -74.635 -6.635 ;
        RECT -74.965 -8.325 -74.635 -7.995 ;
        RECT -74.965 -9.685 -74.635 -9.355 ;
        RECT -74.965 -11.045 -74.635 -10.715 ;
        RECT -74.965 -12.405 -74.635 -12.075 ;
        RECT -74.965 -13.765 -74.635 -13.435 ;
        RECT -74.965 -15.125 -74.635 -14.795 ;
        RECT -74.965 -16.485 -74.635 -16.155 ;
        RECT -74.965 -17.845 -74.635 -17.515 ;
        RECT -74.965 -19.205 -74.635 -18.875 ;
        RECT -74.965 -20.565 -74.635 -20.235 ;
        RECT -74.965 -21.925 -74.635 -21.595 ;
        RECT -74.965 -23.285 -74.635 -22.955 ;
        RECT -74.965 -24.645 -74.635 -24.315 ;
        RECT -74.965 -26.005 -74.635 -25.675 ;
        RECT -74.965 -27.365 -74.635 -27.035 ;
        RECT -74.965 -28.725 -74.635 -28.395 ;
        RECT -74.965 -30.085 -74.635 -29.755 ;
        RECT -74.965 -31.445 -74.635 -31.115 ;
        RECT -74.965 -32.805 -74.635 -32.475 ;
        RECT -74.965 -34.165 -74.635 -33.835 ;
        RECT -74.965 -35.525 -74.635 -35.195 ;
        RECT -74.965 -36.885 -74.635 -36.555 ;
        RECT -74.965 -38.245 -74.635 -37.915 ;
        RECT -74.965 -39.605 -74.635 -39.275 ;
        RECT -74.965 -40.965 -74.635 -40.635 ;
        RECT -74.965 -42.325 -74.635 -41.995 ;
        RECT -74.965 -43.685 -74.635 -43.355 ;
        RECT -74.965 -45.045 -74.635 -44.715 ;
        RECT -74.965 -46.405 -74.635 -46.075 ;
        RECT -74.965 -47.765 -74.635 -47.435 ;
        RECT -74.965 -49.125 -74.635 -48.795 ;
        RECT -74.965 -50.485 -74.635 -50.155 ;
        RECT -74.965 -51.845 -74.635 -51.515 ;
        RECT -74.965 -53.205 -74.635 -52.875 ;
        RECT -74.965 -54.565 -74.635 -54.235 ;
        RECT -74.965 -55.925 -74.635 -55.595 ;
        RECT -74.965 -57.285 -74.635 -56.955 ;
        RECT -74.965 -58.645 -74.635 -58.315 ;
        RECT -74.965 -60.005 -74.635 -59.675 ;
        RECT -74.965 -61.365 -74.635 -61.035 ;
        RECT -74.965 -62.725 -74.635 -62.395 ;
        RECT -74.965 -64.085 -74.635 -63.755 ;
        RECT -74.965 -65.445 -74.635 -65.115 ;
        RECT -74.965 -66.805 -74.635 -66.475 ;
        RECT -74.965 -68.165 -74.635 -67.835 ;
        RECT -74.965 -69.525 -74.635 -69.195 ;
        RECT -74.965 -70.885 -74.635 -70.555 ;
        RECT -74.965 -72.245 -74.635 -71.915 ;
        RECT -74.965 -73.605 -74.635 -73.275 ;
        RECT -74.965 -74.965 -74.635 -74.635 ;
        RECT -74.965 -76.325 -74.635 -75.995 ;
        RECT -74.965 -77.685 -74.635 -77.355 ;
        RECT -74.965 -79.045 -74.635 -78.715 ;
        RECT -74.965 -80.405 -74.635 -80.075 ;
        RECT -74.965 -81.765 -74.635 -81.435 ;
        RECT -74.965 -83.125 -74.635 -82.795 ;
        RECT -74.965 -84.485 -74.635 -84.155 ;
        RECT -74.965 -85.845 -74.635 -85.515 ;
        RECT -74.965 -87.205 -74.635 -86.875 ;
        RECT -74.965 -88.565 -74.635 -88.235 ;
        RECT -74.965 -89.925 -74.635 -89.595 ;
        RECT -74.965 -91.285 -74.635 -90.955 ;
        RECT -74.965 -92.645 -74.635 -92.315 ;
        RECT -74.965 -94.005 -74.635 -93.675 ;
        RECT -74.965 -95.365 -74.635 -95.035 ;
        RECT -74.965 -96.725 -74.635 -96.395 ;
        RECT -74.965 -98.085 -74.635 -97.755 ;
        RECT -74.965 -99.445 -74.635 -99.115 ;
        RECT -74.965 -100.805 -74.635 -100.475 ;
        RECT -74.965 -102.165 -74.635 -101.835 ;
        RECT -74.965 -103.525 -74.635 -103.195 ;
        RECT -74.965 -104.885 -74.635 -104.555 ;
        RECT -74.965 -106.245 -74.635 -105.915 ;
        RECT -74.965 -107.605 -74.635 -107.275 ;
        RECT -74.965 -108.965 -74.635 -108.635 ;
        RECT -74.965 -110.325 -74.635 -109.995 ;
        RECT -74.965 -111.685 -74.635 -111.355 ;
        RECT -74.965 -113.045 -74.635 -112.715 ;
        RECT -74.965 -114.405 -74.635 -114.075 ;
        RECT -74.965 -115.765 -74.635 -115.435 ;
        RECT -74.965 -117.125 -74.635 -116.795 ;
        RECT -74.965 -118.485 -74.635 -118.155 ;
        RECT -74.965 -119.845 -74.635 -119.515 ;
        RECT -74.965 -121.205 -74.635 -120.875 ;
        RECT -74.965 -122.565 -74.635 -122.235 ;
        RECT -74.965 -123.925 -74.635 -123.595 ;
        RECT -74.965 -125.285 -74.635 -124.955 ;
        RECT -74.965 -126.645 -74.635 -126.315 ;
        RECT -74.965 -128.005 -74.635 -127.675 ;
        RECT -74.965 -129.365 -74.635 -129.035 ;
        RECT -74.965 -130.725 -74.635 -130.395 ;
        RECT -74.965 -132.085 -74.635 -131.755 ;
        RECT -74.965 -133.445 -74.635 -133.115 ;
        RECT -74.965 -134.805 -74.635 -134.475 ;
        RECT -74.965 -136.165 -74.635 -135.835 ;
        RECT -74.965 -137.525 -74.635 -137.195 ;
        RECT -74.965 -138.885 -74.635 -138.555 ;
        RECT -74.965 -140.245 -74.635 -139.915 ;
        RECT -74.965 -141.605 -74.635 -141.275 ;
        RECT -74.965 -142.965 -74.635 -142.635 ;
        RECT -74.965 -144.325 -74.635 -143.995 ;
        RECT -74.965 -145.685 -74.635 -145.355 ;
        RECT -74.965 -147.045 -74.635 -146.715 ;
        RECT -74.965 -148.405 -74.635 -148.075 ;
        RECT -74.965 -149.765 -74.635 -149.435 ;
        RECT -74.965 -151.125 -74.635 -150.795 ;
        RECT -74.965 -152.485 -74.635 -152.155 ;
        RECT -74.965 -153.845 -74.635 -153.515 ;
        RECT -74.965 -155.205 -74.635 -154.875 ;
        RECT -74.965 -156.565 -74.635 -156.235 ;
        RECT -74.965 -157.925 -74.635 -157.595 ;
        RECT -74.965 -159.285 -74.635 -158.955 ;
        RECT -74.965 -160.645 -74.635 -160.315 ;
        RECT -74.965 -162.005 -74.635 -161.675 ;
        RECT -74.965 -163.365 -74.635 -163.035 ;
        RECT -74.965 -164.725 -74.635 -164.395 ;
        RECT -74.965 -166.085 -74.635 -165.755 ;
        RECT -74.965 -167.445 -74.635 -167.115 ;
        RECT -74.965 -168.805 -74.635 -168.475 ;
        RECT -74.965 -170.165 -74.635 -169.835 ;
        RECT -74.965 -171.525 -74.635 -171.195 ;
        RECT -74.965 -172.885 -74.635 -172.555 ;
        RECT -74.965 -174.245 -74.635 -173.915 ;
        RECT -74.965 -175.605 -74.635 -175.275 ;
        RECT -74.965 -176.965 -74.635 -176.635 ;
        RECT -74.965 -178.325 -74.635 -177.995 ;
        RECT -74.965 -180.57 -74.635 -179.44 ;
        RECT -74.96 -180.685 -74.64 242.565 ;
        RECT -74.965 241.32 -74.635 242.45 ;
        RECT -74.965 239.195 -74.635 239.525 ;
        RECT -74.965 237.835 -74.635 238.165 ;
        RECT -74.965 236.475 -74.635 236.805 ;
        RECT -74.965 235.115 -74.635 235.445 ;
        RECT -74.965 233.755 -74.635 234.085 ;
        RECT -74.965 232.395 -74.635 232.725 ;
        RECT -74.965 231.035 -74.635 231.365 ;
        RECT -74.965 229.675 -74.635 230.005 ;
        RECT -74.965 228.315 -74.635 228.645 ;
        RECT -74.965 226.955 -74.635 227.285 ;
        RECT -74.965 225.595 -74.635 225.925 ;
        RECT -74.965 224.235 -74.635 224.565 ;
        RECT -74.965 222.875 -74.635 223.205 ;
        RECT -74.965 221.515 -74.635 221.845 ;
        RECT -74.965 220.155 -74.635 220.485 ;
        RECT -74.965 218.795 -74.635 219.125 ;
        RECT -74.965 217.435 -74.635 217.765 ;
        RECT -74.965 216.075 -74.635 216.405 ;
    END
  END vss
  PIN addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -21.24 -183.565 -20.92 -183.245 ;
    END
  END addr[0]
  PIN addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -28.04 -183.565 -27.72 -183.245 ;
    END
  END addr[1]
  PIN addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -34.16 -183.565 -33.84 -183.245 ;
    END
  END addr[2]
  PIN addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -40.28 -183.565 -39.96 -183.245 ;
    END
  END addr[3]
  PIN addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -46.4 -183.565 -46.08 -183.245 ;
    END
  END addr[4]
  PIN addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -52.52 -183.565 -52.2 -183.245 ;
    END
  END addr[5]
  PIN addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -58.64 -183.565 -58.32 -183.245 ;
    END
  END addr[6]
  PIN addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -64.76 -183.565 -64.44 -183.245 ;
    END
  END addr[7]
  PIN addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -70.88 -183.565 -70.56 -183.245 ;
    END
  END addr[8]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -9.68 -183.565 -9.36 -183.245 ;
    END
  END clk
  PIN din[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 5.6 -183.565 6 -183.165 ;
    END
  END din[0]
  PIN din[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 66.6 -183.565 67 -183.165 ;
    END
  END din[10]
  PIN din[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 72.7 -183.565 73.1 -183.165 ;
    END
  END din[11]
  PIN din[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 78.8 -183.565 79.2 -183.165 ;
    END
  END din[12]
  PIN din[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 84.9 -183.565 85.3 -183.165 ;
    END
  END din[13]
  PIN din[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 91 -183.565 91.4 -183.165 ;
    END
  END din[14]
  PIN din[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 97.1 -183.565 97.5 -183.165 ;
    END
  END din[15]
  PIN din[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.2 -183.565 103.6 -183.165 ;
    END
  END din[16]
  PIN din[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 109.3 -183.565 109.7 -183.165 ;
    END
  END din[17]
  PIN din[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 115.4 -183.565 115.8 -183.165 ;
    END
  END din[18]
  PIN din[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 121.5 -183.565 121.9 -183.165 ;
    END
  END din[19]
  PIN din[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 11.7 -183.565 12.1 -183.165 ;
    END
  END din[1]
  PIN din[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 127.6 -183.565 128 -183.165 ;
    END
  END din[20]
  PIN din[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 133.7 -183.565 134.1 -183.165 ;
    END
  END din[21]
  PIN din[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 139.8 -183.565 140.2 -183.165 ;
    END
  END din[22]
  PIN din[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 145.9 -183.565 146.3 -183.165 ;
    END
  END din[23]
  PIN din[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 152 -183.565 152.4 -183.165 ;
    END
  END din[24]
  PIN din[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 158.1 -183.565 158.5 -183.165 ;
    END
  END din[25]
  PIN din[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 164.2 -183.565 164.6 -183.165 ;
    END
  END din[26]
  PIN din[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 170.3 -183.565 170.7 -183.165 ;
    END
  END din[27]
  PIN din[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 176.4 -183.565 176.8 -183.165 ;
    END
  END din[28]
  PIN din[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 182.5 -183.565 182.9 -183.165 ;
    END
  END din[29]
  PIN din[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 17.8 -183.565 18.2 -183.165 ;
    END
  END din[2]
  PIN din[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 188.6 -183.565 189 -183.165 ;
    END
  END din[30]
  PIN din[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 194.7 -183.565 195.1 -183.165 ;
    END
  END din[31]
  PIN din[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 200.8 -183.565 201.2 -183.165 ;
    END
  END din[32]
  PIN din[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 206.9 -183.565 207.3 -183.165 ;
    END
  END din[33]
  PIN din[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 213 -183.565 213.4 -183.165 ;
    END
  END din[34]
  PIN din[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 219.1 -183.565 219.5 -183.165 ;
    END
  END din[35]
  PIN din[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 225.2 -183.565 225.6 -183.165 ;
    END
  END din[36]
  PIN din[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 231.3 -183.565 231.7 -183.165 ;
    END
  END din[37]
  PIN din[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 237.4 -183.565 237.8 -183.165 ;
    END
  END din[38]
  PIN din[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 243.5 -183.565 243.9 -183.165 ;
    END
  END din[39]
  PIN din[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 23.9 -183.565 24.3 -183.165 ;
    END
  END din[3]
  PIN din[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 249.6 -183.565 250 -183.165 ;
    END
  END din[40]
  PIN din[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 255.7 -183.565 256.1 -183.165 ;
    END
  END din[41]
  PIN din[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 261.8 -183.565 262.2 -183.165 ;
    END
  END din[42]
  PIN din[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 267.9 -183.565 268.3 -183.165 ;
    END
  END din[43]
  PIN din[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 274 -183.565 274.4 -183.165 ;
    END
  END din[44]
  PIN din[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 280.1 -183.565 280.5 -183.165 ;
    END
  END din[45]
  PIN din[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 286.2 -183.565 286.6 -183.165 ;
    END
  END din[46]
  PIN din[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 292.3 -183.565 292.7 -183.165 ;
    END
  END din[47]
  PIN din[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 298.4 -183.565 298.8 -183.165 ;
    END
  END din[48]
  PIN din[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 304.5 -183.565 304.9 -183.165 ;
    END
  END din[49]
  PIN din[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 30 -183.565 30.4 -183.165 ;
    END
  END din[4]
  PIN din[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 310.6 -183.565 311 -183.165 ;
    END
  END din[50]
  PIN din[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 316.7 -183.565 317.1 -183.165 ;
    END
  END din[51]
  PIN din[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 322.8 -183.565 323.2 -183.165 ;
    END
  END din[52]
  PIN din[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 328.9 -183.565 329.3 -183.165 ;
    END
  END din[53]
  PIN din[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 335 -183.565 335.4 -183.165 ;
    END
  END din[54]
  PIN din[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 341.1 -183.565 341.5 -183.165 ;
    END
  END din[55]
  PIN din[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 347.2 -183.565 347.6 -183.165 ;
    END
  END din[56]
  PIN din[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 353.3 -183.565 353.7 -183.165 ;
    END
  END din[57]
  PIN din[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 359.4 -183.565 359.8 -183.165 ;
    END
  END din[58]
  PIN din[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 365.5 -183.565 365.9 -183.165 ;
    END
  END din[59]
  PIN din[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.1 -183.565 36.5 -183.165 ;
    END
  END din[5]
  PIN din[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 371.6 -183.565 372 -183.165 ;
    END
  END din[60]
  PIN din[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 377.7 -183.565 378.1 -183.165 ;
    END
  END din[61]
  PIN din[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 383.8 -183.565 384.2 -183.165 ;
    END
  END din[62]
  PIN din[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 389.9 -183.565 390.3 -183.165 ;
    END
  END din[63]
  PIN din[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 42.2 -183.565 42.6 -183.165 ;
    END
  END din[6]
  PIN din[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 48.3 -183.565 48.7 -183.165 ;
    END
  END din[7]
  PIN din[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 54.4 -183.565 54.8 -183.165 ;
    END
  END din[8]
  PIN din[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 60.5 -183.565 60.9 -183.165 ;
    END
  END din[9]
  PIN dout[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 4 -183.565 4.4 -183.165 ;
    END
  END dout[0]
  PIN dout[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 65 -183.565 65.4 -183.165 ;
    END
  END dout[10]
  PIN dout[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71.1 -183.565 71.5 -183.165 ;
    END
  END dout[11]
  PIN dout[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 77.2 -183.565 77.6 -183.165 ;
    END
  END dout[12]
  PIN dout[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 83.3 -183.565 83.7 -183.165 ;
    END
  END dout[13]
  PIN dout[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 89.4 -183.565 89.8 -183.165 ;
    END
  END dout[14]
  PIN dout[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 95.5 -183.565 95.9 -183.165 ;
    END
  END dout[15]
  PIN dout[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 101.6 -183.565 102 -183.165 ;
    END
  END dout[16]
  PIN dout[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 107.7 -183.565 108.1 -183.165 ;
    END
  END dout[17]
  PIN dout[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 113.8 -183.565 114.2 -183.165 ;
    END
  END dout[18]
  PIN dout[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 119.9 -183.565 120.3 -183.165 ;
    END
  END dout[19]
  PIN dout[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 10.1 -183.565 10.5 -183.165 ;
    END
  END dout[1]
  PIN dout[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 126 -183.565 126.4 -183.165 ;
    END
  END dout[20]
  PIN dout[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 132.1 -183.565 132.5 -183.165 ;
    END
  END dout[21]
  PIN dout[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 138.2 -183.565 138.6 -183.165 ;
    END
  END dout[22]
  PIN dout[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 144.3 -183.565 144.7 -183.165 ;
    END
  END dout[23]
  PIN dout[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 150.4 -183.565 150.8 -183.165 ;
    END
  END dout[24]
  PIN dout[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.5 -183.565 156.9 -183.165 ;
    END
  END dout[25]
  PIN dout[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 162.6 -183.565 163 -183.165 ;
    END
  END dout[26]
  PIN dout[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 168.7 -183.565 169.1 -183.165 ;
    END
  END dout[27]
  PIN dout[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 174.8 -183.565 175.2 -183.165 ;
    END
  END dout[28]
  PIN dout[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 180.9 -183.565 181.3 -183.165 ;
    END
  END dout[29]
  PIN dout[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 16.2 -183.565 16.6 -183.165 ;
    END
  END dout[2]
  PIN dout[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 187 -183.565 187.4 -183.165 ;
    END
  END dout[30]
  PIN dout[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 193.1 -183.565 193.5 -183.165 ;
    END
  END dout[31]
  PIN dout[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 199.2 -183.565 199.6 -183.165 ;
    END
  END dout[32]
  PIN dout[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 205.3 -183.565 205.7 -183.165 ;
    END
  END dout[33]
  PIN dout[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 211.4 -183.565 211.8 -183.165 ;
    END
  END dout[34]
  PIN dout[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 217.5 -183.565 217.9 -183.165 ;
    END
  END dout[35]
  PIN dout[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 223.6 -183.565 224 -183.165 ;
    END
  END dout[36]
  PIN dout[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 229.7 -183.565 230.1 -183.165 ;
    END
  END dout[37]
  PIN dout[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 235.8 -183.565 236.2 -183.165 ;
    END
  END dout[38]
  PIN dout[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 241.9 -183.565 242.3 -183.165 ;
    END
  END dout[39]
  PIN dout[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 22.3 -183.565 22.7 -183.165 ;
    END
  END dout[3]
  PIN dout[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 248 -183.565 248.4 -183.165 ;
    END
  END dout[40]
  PIN dout[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 254.1 -183.565 254.5 -183.165 ;
    END
  END dout[41]
  PIN dout[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 260.2 -183.565 260.6 -183.165 ;
    END
  END dout[42]
  PIN dout[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 266.3 -183.565 266.7 -183.165 ;
    END
  END dout[43]
  PIN dout[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 272.4 -183.565 272.8 -183.165 ;
    END
  END dout[44]
  PIN dout[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 278.5 -183.565 278.9 -183.165 ;
    END
  END dout[45]
  PIN dout[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 284.6 -183.565 285 -183.165 ;
    END
  END dout[46]
  PIN dout[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 290.7 -183.565 291.1 -183.165 ;
    END
  END dout[47]
  PIN dout[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 296.8 -183.565 297.2 -183.165 ;
    END
  END dout[48]
  PIN dout[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 302.9 -183.565 303.3 -183.165 ;
    END
  END dout[49]
  PIN dout[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 28.4 -183.565 28.8 -183.165 ;
    END
  END dout[4]
  PIN dout[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 309 -183.565 309.4 -183.165 ;
    END
  END dout[50]
  PIN dout[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 315.1 -183.565 315.5 -183.165 ;
    END
  END dout[51]
  PIN dout[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 321.2 -183.565 321.6 -183.165 ;
    END
  END dout[52]
  PIN dout[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 327.3 -183.565 327.7 -183.165 ;
    END
  END dout[53]
  PIN dout[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 333.4 -183.565 333.8 -183.165 ;
    END
  END dout[54]
  PIN dout[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 339.5 -183.565 339.9 -183.165 ;
    END
  END dout[55]
  PIN dout[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 345.6 -183.565 346 -183.165 ;
    END
  END dout[56]
  PIN dout[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 351.7 -183.565 352.1 -183.165 ;
    END
  END dout[57]
  PIN dout[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 357.8 -183.565 358.2 -183.165 ;
    END
  END dout[58]
  PIN dout[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 363.9 -183.565 364.3 -183.165 ;
    END
  END dout[59]
  PIN dout[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 34.5 -183.565 34.9 -183.165 ;
    END
  END dout[5]
  PIN dout[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 370 -183.565 370.4 -183.165 ;
    END
  END dout[60]
  PIN dout[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 376.1 -183.565 376.5 -183.165 ;
    END
  END dout[61]
  PIN dout[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 382.2 -183.565 382.6 -183.165 ;
    END
  END dout[62]
  PIN dout[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 388.3 -183.565 388.7 -183.165 ;
    END
  END dout[63]
  PIN dout[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 40.6 -183.565 41 -183.165 ;
    END
  END dout[6]
  PIN dout[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 46.7 -183.565 47.1 -183.165 ;
    END
  END dout[7]
  PIN dout[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 52.8 -183.565 53.2 -183.165 ;
    END
  END dout[8]
  PIN dout[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 58.9 -183.565 59.3 -183.165 ;
    END
  END dout[9]
  PIN we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -15.12 -183.565 -14.8 -183.245 ;
    END
  END we
  PIN wmask[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 6.4 -183.565 6.8 -183.165 ;
    END
  END wmask[0]
  PIN wmask[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 55.2 -183.565 55.6 -183.165 ;
    END
  END wmask[1]
  PIN wmask[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 104 -183.565 104.4 -183.165 ;
    END
  END wmask[2]
  PIN wmask[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 152.8 -183.565 153.2 -183.165 ;
    END
  END wmask[3]
  PIN wmask[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 201.6 -183.565 202 -183.165 ;
    END
  END wmask[4]
  PIN wmask[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 250.4 -183.565 250.8 -183.165 ;
    END
  END wmask[5]
  PIN wmask[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 299.2 -183.565 299.6 -183.165 ;
    END
  END wmask[6]
  PIN wmask[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 348 -183.565 348.4 -183.165 ;
    END
  END wmask[7]
  OBS
    LAYER met1 SPACING 0.14 ;
      RECT -80.225 -183.565 407.985 245.445 ;
    LAYER met2 SPACING 0.14 ;
      RECT -80.225 -183.565 407.985 245.445 ;
    LAYER met3 SPACING 0.3 ;
      RECT 0.515 -34.845 0.845 -34.515 ;
      RECT 0.52 -49.805 0.84 -34.515 ;
      RECT 0.515 -49.805 0.845 -49.475 ;
      RECT -0.165 -34.165 0.165 -33.835 ;
      RECT -0.16 -34.845 0.16 -33.835 ;
      RECT -0.165 -34.845 0.165 -34.515 ;
      RECT -8.325 -1.525 -7.995 -1.195 ;
      RECT -8.32 -121.205 -8 -1.195 ;
      RECT -8.325 -11.045 -7.995 -10.715 ;
      RECT -8.325 -121.205 -7.995 -120.875 ;
      RECT -9.005 -19.885 -8.675 -19.555 ;
      RECT -9 -108.965 -8.68 -19.555 ;
      RECT -9.005 -108.965 -8.675 -108.635 ;
      RECT -9.685 -86.525 -9.355 -86.195 ;
      RECT -9.68 -182.755 -9.36 -86.195 ;
      RECT -9.685 -157.925 -9.355 -157.595 ;
      RECT -9.685 -171.525 -9.355 -171.195 ;
      RECT -10.365 -167.445 -10.035 -167.115 ;
      RECT -10.36 -172.885 -10.04 -167.115 ;
      RECT -10.365 -172.885 -10.035 -172.555 ;
      RECT -12.405 -13.765 -12.075 -13.435 ;
      RECT -12.4 -26.005 -12.08 -13.435 ;
      RECT -12.405 -26.005 -12.075 -25.675 ;
      RECT -13.085 -18.525 -12.755 -18.195 ;
      RECT -13.08 -108.285 -12.76 -18.195 ;
      RECT -13.085 -108.285 -12.755 -107.955 ;
      RECT -14.445 -110.13 -14.115 -109.8 ;
      RECT -14.44 -112.365 -14.12 -109.8 ;
      RECT -14.445 -112.365 -14.115 -112.035 ;
      RECT -15.125 -172.885 -14.795 -172.555 ;
      RECT -15.12 -182.755 -14.8 -172.555 ;
      RECT -15.125 -110.61 -14.795 -110.28 ;
      RECT -15.12 -113.045 -14.8 -110.28 ;
      RECT -15.125 -113.045 -14.795 -112.715 ;
      RECT -15.805 -111.09 -15.475 -110.76 ;
      RECT -15.8 -113.725 -15.48 -110.76 ;
      RECT -15.805 -113.725 -15.475 -113.395 ;
      RECT -15.805 -20.565 -15.475 -20.235 ;
      RECT -15.8 -101.485 -15.48 -20.235 ;
      RECT -15.805 -101.485 -15.475 -101.155 ;
      RECT -16.485 -111.57 -16.155 -111.24 ;
      RECT -16.48 -173.565 -16.16 -111.24 ;
      RECT -16.485 -173.565 -16.155 -173.235 ;
      RECT -16.485 -13.085 -16.155 -12.755 ;
      RECT -16.48 -26.005 -16.16 -12.755 ;
      RECT -16.485 -26.005 -16.155 -25.675 ;
      RECT -17.165 -113.725 -16.835 -113.395 ;
      RECT -17.16 -172.205 -16.84 -113.395 ;
      RECT -17.165 -172.205 -16.835 -171.875 ;
      RECT -17.165 -12.405 -16.835 -12.075 ;
      RECT -17.16 -26.005 -16.84 -12.075 ;
      RECT -17.165 -26.005 -16.835 -25.675 ;
      RECT -17.845 -11.725 -17.515 -11.395 ;
      RECT -17.84 -26.005 -17.52 -11.395 ;
      RECT -17.845 -26.005 -17.515 -25.675 ;
      RECT -18.525 -113.045 -18.195 -112.715 ;
      RECT -18.52 -173.565 -18.2 -112.715 ;
      RECT -18.525 -173.565 -18.195 -173.235 ;
      RECT -18.525 -22.49 -18.195 -22.16 ;
      RECT -18.52 -26.005 -18.2 -22.16 ;
      RECT -18.525 -26.005 -18.195 -25.675 ;
      RECT -19.205 -22.97 -18.875 -22.64 ;
      RECT -19.2 -26.685 -18.88 -22.64 ;
      RECT -19.205 -26.685 -18.875 -26.355 ;
      RECT -19.885 -23.45 -19.555 -23.12 ;
      RECT -19.88 -27.365 -19.56 -23.12 ;
      RECT -19.885 -27.365 -19.555 -27.035 ;
      RECT -20.565 -23.93 -20.235 -23.6 ;
      RECT -20.56 -28.045 -20.24 -23.6 ;
      RECT -20.565 -28.045 -20.235 -27.715 ;
      RECT -21.245 -172.885 -20.915 -172.555 ;
      RECT -21.24 -182.755 -20.92 -172.555 ;
      RECT -21.245 -88.565 -20.915 -88.235 ;
      RECT -21.24 -119.165 -20.92 -88.235 ;
      RECT -21.245 -119.165 -20.915 -118.835 ;
      RECT -21.245 -24.41 -20.915 -24.08 ;
      RECT -21.24 -62.725 -20.92 -24.08 ;
      RECT -21.245 -62.725 -20.915 -62.395 ;
      RECT -21.925 -24.89 -21.595 -24.56 ;
      RECT -21.92 -63.405 -21.6 -24.56 ;
      RECT -21.925 -63.405 -21.595 -63.075 ;
      RECT -23.285 -112.365 -22.955 -112.035 ;
      RECT -23.28 -172.205 -22.96 -112.035 ;
      RECT -23.285 -172.205 -22.955 -171.875 ;
      RECT -28.045 -172.885 -27.715 -172.555 ;
      RECT -28.04 -182.755 -27.72 -172.555 ;
      RECT -28.725 -64.33 -28.395 -64 ;
      RECT -28.72 -66.805 -28.4 -64 ;
      RECT -28.725 -66.805 -28.395 -66.475 ;
      RECT -29.405 -112.365 -29.075 -112.035 ;
      RECT -29.4 -173.565 -29.08 -112.035 ;
      RECT -29.405 -173.565 -29.075 -173.235 ;
      RECT -29.405 -64.81 -29.075 -64.48 ;
      RECT -29.4 -67.485 -29.08 -64.48 ;
      RECT -29.405 -67.485 -29.075 -67.155 ;
      RECT -30.085 -112.365 -29.755 -112.035 ;
      RECT -30.08 -172.205 -29.76 -112.035 ;
      RECT -30.085 -172.205 -29.755 -171.875 ;
      RECT -30.085 -65.29 -29.755 -64.96 ;
      RECT -30.08 -68.165 -29.76 -64.96 ;
      RECT -30.085 -68.165 -29.755 -67.835 ;
      RECT -30.765 -65.77 -30.435 -65.44 ;
      RECT -30.76 -68.845 -30.44 -65.44 ;
      RECT -30.765 -68.845 -30.435 -68.515 ;
      RECT -34.165 -172.885 -33.835 -172.555 ;
      RECT -34.16 -182.755 -33.84 -172.555 ;
      RECT -34.845 -113.045 -34.515 -112.715 ;
      RECT -34.84 -173.565 -34.52 -112.715 ;
      RECT -34.845 -173.565 -34.515 -173.235 ;
      RECT -35.525 -112.365 -35.195 -112.035 ;
      RECT -35.52 -172.205 -35.2 -112.035 ;
      RECT -35.525 -172.205 -35.195 -171.875 ;
      RECT -40.285 -172.885 -39.955 -172.555 ;
      RECT -40.28 -182.755 -39.96 -172.555 ;
      RECT -41.645 -112.365 -41.315 -112.035 ;
      RECT -41.64 -172.205 -41.32 -112.035 ;
      RECT -41.645 -172.205 -41.315 -171.875 ;
      RECT -42.325 -113.045 -41.995 -112.715 ;
      RECT -42.32 -173.565 -42 -112.715 ;
      RECT -42.325 -173.565 -41.995 -173.235 ;
      RECT -43.005 -64.33 -42.675 -64 ;
      RECT -43 -66.805 -42.68 -64 ;
      RECT -43.005 -66.805 -42.675 -66.475 ;
      RECT -43.685 -64.81 -43.355 -64.48 ;
      RECT -43.68 -67.485 -43.36 -64.48 ;
      RECT -43.685 -67.485 -43.355 -67.155 ;
      RECT -44.365 -65.29 -44.035 -64.96 ;
      RECT -44.36 -68.165 -44.04 -64.96 ;
      RECT -44.365 -68.165 -44.035 -67.835 ;
      RECT -45.045 -65.77 -44.715 -65.44 ;
      RECT -45.04 -68.845 -44.72 -65.44 ;
      RECT -45.045 -68.845 -44.715 -68.515 ;
      RECT -46.405 -172.885 -46.075 -172.555 ;
      RECT -46.4 -182.755 -46.08 -172.555 ;
      RECT -46.405 -112.365 -46.075 -112.035 ;
      RECT -46.4 -172.205 -46.08 -112.035 ;
      RECT -46.405 -172.205 -46.075 -171.875 ;
      RECT -46.405 -2.205 -46.075 -1.875 ;
      RECT -46.4 -28.725 -46.08 -1.875 ;
      RECT -46.405 -28.725 -46.075 -28.395 ;
      RECT -47.085 -2.205 -46.755 -1.875 ;
      RECT -47.08 -29.405 -46.76 -1.875 ;
      RECT -47.085 -29.405 -46.755 -29.075 ;
      RECT -48.445 -113.725 -48.115 -113.395 ;
      RECT -48.44 -173.565 -48.12 -113.395 ;
      RECT -48.445 -173.565 -48.115 -173.235 ;
      RECT -52.525 -172.885 -52.195 -172.555 ;
      RECT -52.52 -182.755 -52.2 -172.555 ;
      RECT -52.525 -112.365 -52.195 -112.035 ;
      RECT -52.52 -172.205 -52.2 -112.035 ;
      RECT -52.525 -172.205 -52.195 -171.875 ;
      RECT -53.48 116.48 -52.2 117.12 ;
      RECT -52.52 -110.325 -52.2 117.12 ;
      RECT -52.525 -110.325 -52.195 -109.995 ;
      RECT -54.565 -113.045 -54.235 -112.715 ;
      RECT -54.56 -173.565 -54.24 -112.715 ;
      RECT -54.565 -173.565 -54.235 -173.235 ;
      RECT -58.645 -172.885 -58.315 -172.555 ;
      RECT -58.64 -182.755 -58.32 -172.555 ;
      RECT -58.645 -113.725 -58.315 -113.395 ;
      RECT -58.64 -172.205 -58.32 -113.395 ;
      RECT -58.645 -172.205 -58.315 -171.875 ;
      RECT -59.325 86.875 -58.995 87.205 ;
      RECT -59.32 -1.525 -59 87.205 ;
      RECT -59.325 -1.525 -58.995 -1.195 ;
      RECT -60.005 86.195 -59.675 86.525 ;
      RECT -60 -121.205 -59.68 86.525 ;
      RECT -60.005 -121.205 -59.675 -120.875 ;
      RECT -60.685 -114.405 -60.355 -114.075 ;
      RECT -60.68 -173.565 -60.36 -114.075 ;
      RECT -60.685 -173.565 -60.355 -173.235 ;
      RECT -61.365 -113.045 -61.035 -112.715 ;
      RECT -61.36 -173.565 -61.04 -112.715 ;
      RECT -61.365 -173.565 -61.035 -173.235 ;
      RECT -62.045 -111.685 -61.715 -111.355 ;
      RECT -62.04 -119.845 -61.72 -111.355 ;
      RECT -62.045 -119.845 -61.715 -119.515 ;
      RECT -64.765 -172.885 -64.435 -172.555 ;
      RECT -64.76 -182.755 -64.44 -172.555 ;
      RECT -64.765 -112.365 -64.435 -112.035 ;
      RECT -64.76 -172.205 -64.44 -112.035 ;
      RECT -64.765 -172.205 -64.435 -171.875 ;
      RECT -70.885 -172.885 -70.555 -172.555 ;
      RECT -70.88 -182.755 -70.56 -172.555 ;
      RECT 391.5 -80.215 391.9 -20.12 ;
      RECT 390.7 -79.355 391.1 -20.12 ;
      RECT 389.9 -182.675 390.3 -79.445 ;
      RECT 389.1 -63.5 389.5 -48.905 ;
      RECT 389.1 -45.08 389.5 -15.74 ;
      RECT 388.3 -182.675 388.7 -73.605 ;
      RECT 388.3 -64 388.7 -49.36 ;
      RECT 388.3 -45.51 388.7 -12.47 ;
      RECT 385.4 -80.215 385.8 -20.12 ;
      RECT 384.6 -79.355 385 -20.12 ;
      RECT 383.8 -182.675 384.2 -79.445 ;
      RECT 383 -63.5 383.4 -48.905 ;
      RECT 383 -45.08 383.4 -15.74 ;
      RECT 382.2 -182.675 382.6 -73.605 ;
      RECT 382.2 -64 382.6 -49.36 ;
      RECT 382.2 -45.51 382.6 -12.47 ;
      RECT 379.3 -80.215 379.7 -20.12 ;
      RECT 378.5 -79.355 378.9 -20.12 ;
      RECT 377.7 -182.675 378.1 -79.445 ;
      RECT 376.9 -63.5 377.3 -48.905 ;
      RECT 376.9 -45.08 377.3 -15.74 ;
      RECT 376.1 -182.675 376.5 -73.605 ;
      RECT 376.1 -64 376.5 -49.36 ;
      RECT 376.1 -45.51 376.5 -12.47 ;
      RECT 373.2 -80.215 373.6 -20.12 ;
      RECT 372.4 -79.355 372.8 -20.12 ;
      RECT 371.6 -182.675 372 -79.445 ;
      RECT 370.8 -63.5 371.2 -48.905 ;
      RECT 370.8 -45.08 371.2 -15.74 ;
      RECT 370 -182.675 370.4 -73.605 ;
      RECT 370 -64 370.4 -49.36 ;
      RECT 370 -45.51 370.4 -12.47 ;
      RECT 367.1 -80.215 367.5 -20.12 ;
      RECT 366.3 -79.355 366.7 -20.12 ;
      RECT 365.5 -182.675 365.9 -79.445 ;
      RECT 364.7 -63.5 365.1 -48.905 ;
      RECT 364.7 -45.08 365.1 -15.74 ;
      RECT 363.9 -182.675 364.3 -73.605 ;
      RECT 363.9 -64 364.3 -49.36 ;
      RECT 363.9 -45.51 364.3 -12.47 ;
      RECT 361 -80.215 361.4 -20.12 ;
      RECT 360.2 -79.355 360.6 -20.12 ;
      RECT 359.4 -182.675 359.8 -79.445 ;
      RECT 358.6 -63.5 359 -48.905 ;
      RECT 358.6 -45.08 359 -15.74 ;
      RECT 357.8 -182.675 358.2 -73.605 ;
      RECT 357.8 -64 358.2 -49.36 ;
      RECT 357.8 -45.51 358.2 -12.47 ;
      RECT 354.9 -80.215 355.3 -20.12 ;
      RECT 354.1 -79.355 354.5 -20.12 ;
      RECT 353.3 -182.675 353.7 -79.445 ;
      RECT 352.5 -63.5 352.9 -48.905 ;
      RECT 352.5 -45.08 352.9 -15.74 ;
      RECT 351.7 -182.675 352.1 -73.605 ;
      RECT 351.7 -64 352.1 -49.36 ;
      RECT 351.7 -45.51 352.1 -12.47 ;
      RECT 349.6 -87.06 350 -20.12 ;
      RECT 348.8 -80.215 349.2 -20.12 ;
      RECT 348 -182.675 348.4 -87.15 ;
      RECT 348 -79.355 348.4 -20.12 ;
      RECT 347.2 -182.675 347.6 -79.445 ;
      RECT 346.4 -63.5 346.8 -48.905 ;
      RECT 346.4 -45.08 346.8 -15.74 ;
      RECT 345.6 -182.675 346 -73.605 ;
      RECT 345.6 -64 346 -49.36 ;
      RECT 345.6 -45.51 346 -12.47 ;
      RECT 342.7 -80.215 343.1 -20.12 ;
      RECT 341.9 -79.355 342.3 -20.12 ;
      RECT 341.1 -182.675 341.5 -79.445 ;
      RECT 340.3 -63.5 340.7 -48.905 ;
      RECT 340.3 -45.08 340.7 -15.74 ;
      RECT 339.5 -182.675 339.9 -73.605 ;
      RECT 339.5 -64 339.9 -49.36 ;
      RECT 339.5 -45.51 339.9 -12.47 ;
      RECT 336.6 -80.215 337 -20.12 ;
      RECT 335.8 -79.355 336.2 -20.12 ;
      RECT 335 -182.675 335.4 -79.445 ;
      RECT 334.2 -63.5 334.6 -48.905 ;
      RECT 334.2 -45.08 334.6 -15.74 ;
      RECT 333.4 -182.675 333.8 -73.605 ;
      RECT 333.4 -64 333.8 -49.36 ;
      RECT 333.4 -45.51 333.8 -12.47 ;
      RECT 330.5 -80.215 330.9 -20.12 ;
      RECT 329.7 -79.355 330.1 -20.12 ;
      RECT 328.9 -182.675 329.3 -79.445 ;
      RECT 328.1 -63.5 328.5 -48.905 ;
      RECT 328.1 -45.08 328.5 -15.74 ;
      RECT 327.3 -182.675 327.7 -73.605 ;
      RECT 327.3 -64 327.7 -49.36 ;
      RECT 327.3 -45.51 327.7 -12.47 ;
      RECT 324.4 -80.215 324.8 -20.12 ;
      RECT 323.6 -79.355 324 -20.12 ;
      RECT 322.8 -182.675 323.2 -79.445 ;
      RECT 322 -63.5 322.4 -48.905 ;
      RECT 322 -45.08 322.4 -15.74 ;
      RECT 321.2 -182.675 321.6 -73.605 ;
      RECT 321.2 -64 321.6 -49.36 ;
      RECT 321.2 -45.51 321.6 -12.47 ;
      RECT 318.3 -80.215 318.7 -20.12 ;
      RECT 317.5 -79.355 317.9 -20.12 ;
      RECT 316.7 -182.675 317.1 -79.445 ;
      RECT 315.9 -63.5 316.3 -48.905 ;
      RECT 315.9 -45.08 316.3 -15.74 ;
      RECT 315.1 -182.675 315.5 -73.605 ;
      RECT 315.1 -64 315.5 -49.36 ;
      RECT 315.1 -45.51 315.5 -12.47 ;
      RECT 312.2 -80.215 312.6 -20.12 ;
      RECT 311.4 -79.355 311.8 -20.12 ;
      RECT 310.6 -182.675 311 -79.445 ;
      RECT 309.8 -63.5 310.2 -48.905 ;
      RECT 309.8 -45.08 310.2 -15.74 ;
      RECT 309 -182.675 309.4 -73.605 ;
      RECT 309 -64 309.4 -49.36 ;
      RECT 309 -45.51 309.4 -12.47 ;
      RECT 306.1 -80.215 306.5 -20.12 ;
      RECT 305.3 -79.355 305.7 -20.12 ;
      RECT 304.5 -182.675 304.9 -79.445 ;
      RECT 303.7 -63.5 304.1 -48.905 ;
      RECT 303.7 -45.08 304.1 -15.74 ;
      RECT 302.9 -182.675 303.3 -73.605 ;
      RECT 302.9 -64 303.3 -49.36 ;
      RECT 302.9 -45.51 303.3 -12.47 ;
      RECT 300.8 -87.06 301.2 -20.12 ;
      RECT 300 -80.215 300.4 -20.12 ;
      RECT 299.2 -182.675 299.6 -87.15 ;
      RECT 299.2 -79.355 299.6 -20.12 ;
      RECT 298.4 -182.675 298.8 -79.445 ;
      RECT 297.6 -63.5 298 -48.905 ;
      RECT 297.6 -45.08 298 -15.74 ;
      RECT 296.8 -182.675 297.2 -73.605 ;
      RECT 296.8 -64 297.2 -49.36 ;
      RECT 296.8 -45.51 297.2 -12.47 ;
      RECT 293.9 -80.215 294.3 -20.12 ;
      RECT 293.1 -79.355 293.5 -20.12 ;
      RECT 292.3 -182.675 292.7 -79.445 ;
      RECT 291.5 -63.5 291.9 -48.905 ;
      RECT 291.5 -45.08 291.9 -15.74 ;
      RECT 290.7 -182.675 291.1 -73.605 ;
      RECT 290.7 -64 291.1 -49.36 ;
      RECT 290.7 -45.51 291.1 -12.47 ;
      RECT 287.8 -80.215 288.2 -20.12 ;
      RECT 287 -79.355 287.4 -20.12 ;
      RECT 286.2 -182.675 286.6 -79.445 ;
      RECT 285.4 -63.5 285.8 -48.905 ;
      RECT 285.4 -45.08 285.8 -15.74 ;
      RECT 284.6 -182.675 285 -73.605 ;
      RECT 284.6 -64 285 -49.36 ;
      RECT 284.6 -45.51 285 -12.47 ;
      RECT 281.7 -80.215 282.1 -20.12 ;
      RECT 280.9 -79.355 281.3 -20.12 ;
      RECT 280.1 -182.675 280.5 -79.445 ;
      RECT 279.3 -63.5 279.7 -48.905 ;
      RECT 279.3 -45.08 279.7 -15.74 ;
      RECT 278.5 -182.675 278.9 -73.605 ;
      RECT 278.5 -64 278.9 -49.36 ;
      RECT 278.5 -45.51 278.9 -12.47 ;
      RECT 275.6 -80.215 276 -20.12 ;
      RECT 274.8 -79.355 275.2 -20.12 ;
      RECT 274 -182.675 274.4 -79.445 ;
      RECT 273.2 -63.5 273.6 -48.905 ;
      RECT 273.2 -45.08 273.6 -15.74 ;
      RECT 272.4 -182.675 272.8 -73.605 ;
      RECT 272.4 -64 272.8 -49.36 ;
      RECT 272.4 -45.51 272.8 -12.47 ;
      RECT 269.5 -80.215 269.9 -20.12 ;
      RECT 268.7 -79.355 269.1 -20.12 ;
      RECT 267.9 -182.675 268.3 -79.445 ;
      RECT 267.1 -63.5 267.5 -48.905 ;
      RECT 267.1 -45.08 267.5 -15.74 ;
      RECT 266.3 -182.675 266.7 -73.605 ;
      RECT 266.3 -64 266.7 -49.36 ;
      RECT 266.3 -45.51 266.7 -12.47 ;
      RECT 263.4 -80.215 263.8 -20.12 ;
      RECT 262.6 -79.355 263 -20.12 ;
      RECT 261.8 -182.675 262.2 -79.445 ;
      RECT 261 -63.5 261.4 -48.905 ;
      RECT 261 -45.08 261.4 -15.74 ;
      RECT 260.2 -182.675 260.6 -73.605 ;
      RECT 260.2 -64 260.6 -49.36 ;
      RECT 260.2 -45.51 260.6 -12.47 ;
      RECT 257.3 -80.215 257.7 -20.12 ;
      RECT 256.5 -79.355 256.9 -20.12 ;
      RECT 255.7 -182.675 256.1 -79.445 ;
      RECT 254.9 -63.5 255.3 -48.905 ;
      RECT 254.9 -45.08 255.3 -15.74 ;
      RECT 254.1 -182.675 254.5 -73.605 ;
      RECT 254.1 -64 254.5 -49.36 ;
      RECT 254.1 -45.51 254.5 -12.47 ;
      RECT 252 -87.06 252.4 -20.12 ;
      RECT 251.2 -80.215 251.6 -20.12 ;
      RECT 250.4 -182.675 250.8 -87.15 ;
      RECT 250.4 -79.355 250.8 -20.12 ;
      RECT 249.6 -182.675 250 -79.445 ;
      RECT 248.8 -63.5 249.2 -48.905 ;
      RECT 248.8 -45.08 249.2 -15.74 ;
      RECT 248 -182.675 248.4 -73.605 ;
      RECT 248 -64 248.4 -49.36 ;
      RECT 248 -45.51 248.4 -12.47 ;
      RECT 245.1 -80.215 245.5 -20.12 ;
      RECT 244.3 -79.355 244.7 -20.12 ;
      RECT 243.5 -182.675 243.9 -79.445 ;
      RECT 242.7 -63.5 243.1 -48.905 ;
      RECT 242.7 -45.08 243.1 -15.74 ;
      RECT 241.9 -182.675 242.3 -73.605 ;
      RECT 241.9 -64 242.3 -49.36 ;
      RECT 241.9 -45.51 242.3 -12.47 ;
      RECT 239 -80.215 239.4 -20.12 ;
      RECT 238.2 -79.355 238.6 -20.12 ;
      RECT 237.4 -182.675 237.8 -79.445 ;
      RECT 236.6 -63.5 237 -48.905 ;
      RECT 236.6 -45.08 237 -15.74 ;
      RECT 235.8 -182.675 236.2 -73.605 ;
      RECT 235.8 -64 236.2 -49.36 ;
      RECT 235.8 -45.51 236.2 -12.47 ;
      RECT 232.9 -80.215 233.3 -20.12 ;
      RECT 232.1 -79.355 232.5 -20.12 ;
      RECT 231.3 -182.675 231.7 -79.445 ;
      RECT 230.5 -63.5 230.9 -48.905 ;
      RECT 230.5 -45.08 230.9 -15.74 ;
      RECT 229.7 -182.675 230.1 -73.605 ;
      RECT 229.7 -64 230.1 -49.36 ;
      RECT 229.7 -45.51 230.1 -12.47 ;
      RECT 226.8 -80.215 227.2 -20.12 ;
      RECT 226 -79.355 226.4 -20.12 ;
      RECT 225.2 -182.675 225.6 -79.445 ;
      RECT 224.4 -63.5 224.8 -48.905 ;
      RECT 224.4 -45.08 224.8 -15.74 ;
      RECT 223.6 -182.675 224 -73.605 ;
      RECT 223.6 -64 224 -49.36 ;
      RECT 223.6 -45.51 224 -12.47 ;
      RECT 220.7 -80.215 221.1 -20.12 ;
      RECT 219.9 -79.355 220.3 -20.12 ;
      RECT 219.1 -182.675 219.5 -79.445 ;
      RECT 218.3 -63.5 218.7 -48.905 ;
      RECT 218.3 -45.08 218.7 -15.74 ;
      RECT 217.5 -182.675 217.9 -73.605 ;
      RECT 217.5 -64 217.9 -49.36 ;
      RECT 217.5 -45.51 217.9 -12.47 ;
      RECT 214.6 -80.215 215 -20.12 ;
      RECT 213.8 -79.355 214.2 -20.12 ;
      RECT 213 -182.675 213.4 -79.445 ;
      RECT 212.2 -63.5 212.6 -48.905 ;
      RECT 212.2 -45.08 212.6 -15.74 ;
      RECT 211.4 -182.675 211.8 -73.605 ;
      RECT 211.4 -64 211.8 -49.36 ;
      RECT 211.4 -45.51 211.8 -12.47 ;
      RECT 208.5 -80.215 208.9 -20.12 ;
      RECT 207.7 -79.355 208.1 -20.12 ;
      RECT 206.9 -182.675 207.3 -79.445 ;
      RECT 206.1 -63.5 206.5 -48.905 ;
      RECT 206.1 -45.08 206.5 -15.74 ;
      RECT 205.3 -182.675 205.7 -73.605 ;
      RECT 205.3 -64 205.7 -49.36 ;
      RECT 205.3 -45.51 205.7 -12.47 ;
      RECT 203.2 -87.06 203.6 -20.12 ;
      RECT 202.4 -80.215 202.8 -20.12 ;
      RECT 201.6 -182.675 202 -87.15 ;
      RECT 201.6 -79.355 202 -20.12 ;
      RECT 200.8 -182.675 201.2 -79.445 ;
      RECT 200 -63.5 200.4 -48.905 ;
      RECT 200 -45.08 200.4 -15.74 ;
      RECT 199.2 -182.675 199.6 -73.605 ;
      RECT 199.2 -64 199.6 -49.36 ;
      RECT 199.2 -45.51 199.6 -12.47 ;
      RECT 196.3 -80.215 196.7 -20.12 ;
      RECT 195.5 -79.355 195.9 -20.12 ;
      RECT 194.7 -182.675 195.1 -79.445 ;
      RECT 193.9 -63.5 194.3 -48.905 ;
      RECT 193.9 -45.08 194.3 -15.74 ;
      RECT 193.1 -182.675 193.5 -73.605 ;
      RECT 193.1 -64 193.5 -49.36 ;
      RECT 193.1 -45.51 193.5 -12.47 ;
      RECT 190.2 -80.215 190.6 -20.12 ;
      RECT 189.4 -79.355 189.8 -20.12 ;
      RECT 188.6 -182.675 189 -79.445 ;
      RECT 187.8 -63.5 188.2 -48.905 ;
      RECT 187.8 -45.08 188.2 -15.74 ;
      RECT 187 -182.675 187.4 -73.605 ;
      RECT 187 -64 187.4 -49.36 ;
      RECT 187 -45.51 187.4 -12.47 ;
      RECT 184.1 -80.215 184.5 -20.12 ;
      RECT 183.3 -79.355 183.7 -20.12 ;
      RECT 182.5 -182.675 182.9 -79.445 ;
      RECT 181.7 -63.5 182.1 -48.905 ;
      RECT 181.7 -45.08 182.1 -15.74 ;
      RECT 180.9 -182.675 181.3 -73.605 ;
      RECT 180.9 -64 181.3 -49.36 ;
      RECT 180.9 -45.51 181.3 -12.47 ;
      RECT 178 -80.215 178.4 -20.12 ;
      RECT 177.2 -79.355 177.6 -20.12 ;
      RECT 176.4 -182.675 176.8 -79.445 ;
      RECT 175.6 -63.5 176 -48.905 ;
      RECT 175.6 -45.08 176 -15.74 ;
      RECT 174.8 -182.675 175.2 -73.605 ;
      RECT 174.8 -64 175.2 -49.36 ;
      RECT 174.8 -45.51 175.2 -12.47 ;
      RECT 171.9 -80.215 172.3 -20.12 ;
      RECT 171.1 -79.355 171.5 -20.12 ;
      RECT 170.3 -182.675 170.7 -79.445 ;
      RECT 169.5 -63.5 169.9 -48.905 ;
      RECT 169.5 -45.08 169.9 -15.74 ;
      RECT 168.7 -182.675 169.1 -73.605 ;
      RECT 168.7 -64 169.1 -49.36 ;
      RECT 168.7 -45.51 169.1 -12.47 ;
      RECT 165.8 -80.215 166.2 -20.12 ;
      RECT 165 -79.355 165.4 -20.12 ;
      RECT 164.2 -182.675 164.6 -79.445 ;
      RECT 163.4 -63.5 163.8 -48.905 ;
      RECT 163.4 -45.08 163.8 -15.74 ;
      RECT 162.6 -182.675 163 -73.605 ;
      RECT 162.6 -64 163 -49.36 ;
      RECT 162.6 -45.51 163 -12.47 ;
      RECT 159.7 -80.215 160.1 -20.12 ;
      RECT 158.9 -79.355 159.3 -20.12 ;
      RECT 158.1 -182.675 158.5 -79.445 ;
      RECT 157.3 -63.5 157.7 -48.905 ;
      RECT 157.3 -45.08 157.7 -15.74 ;
      RECT 156.5 -182.675 156.9 -73.605 ;
      RECT 156.5 -64 156.9 -49.36 ;
      RECT 156.5 -45.51 156.9 -12.47 ;
      RECT 154.4 -87.06 154.8 -20.12 ;
      RECT 153.6 -80.215 154 -20.12 ;
      RECT 152.8 -182.675 153.2 -87.15 ;
      RECT 152.8 -79.355 153.2 -20.12 ;
      RECT 152 -182.675 152.4 -79.445 ;
      RECT 151.2 -63.5 151.6 -48.905 ;
      RECT 151.2 -45.08 151.6 -15.74 ;
      RECT 150.4 -182.675 150.8 -73.605 ;
      RECT 150.4 -64 150.8 -49.36 ;
      RECT 150.4 -45.51 150.8 -12.47 ;
      RECT 147.5 -80.215 147.9 -20.12 ;
      RECT 146.7 -79.355 147.1 -20.12 ;
      RECT 145.9 -182.675 146.3 -79.445 ;
      RECT 145.1 -63.5 145.5 -48.905 ;
      RECT 145.1 -45.08 145.5 -15.74 ;
      RECT 144.3 -182.675 144.7 -73.605 ;
      RECT 144.3 -64 144.7 -49.36 ;
      RECT 144.3 -45.51 144.7 -12.47 ;
      RECT 141.4 -80.215 141.8 -20.12 ;
      RECT 140.6 -79.355 141 -20.12 ;
      RECT 139.8 -182.675 140.2 -79.445 ;
      RECT 139 -63.5 139.4 -48.905 ;
      RECT 139 -45.08 139.4 -15.74 ;
      RECT 138.2 -182.675 138.6 -73.605 ;
      RECT 138.2 -64 138.6 -49.36 ;
      RECT 138.2 -45.51 138.6 -12.47 ;
      RECT 135.3 -80.215 135.7 -20.12 ;
      RECT 134.5 -79.355 134.9 -20.12 ;
      RECT 133.7 -182.675 134.1 -79.445 ;
      RECT 132.9 -63.5 133.3 -48.905 ;
      RECT 132.9 -45.08 133.3 -15.74 ;
      RECT 132.1 -182.675 132.5 -73.605 ;
      RECT 132.1 -64 132.5 -49.36 ;
      RECT 132.1 -45.51 132.5 -12.47 ;
      RECT 129.2 -80.215 129.6 -20.12 ;
      RECT 128.4 -79.355 128.8 -20.12 ;
      RECT 127.6 -182.675 128 -79.445 ;
      RECT 126.8 -63.5 127.2 -48.905 ;
      RECT 126.8 -45.08 127.2 -15.74 ;
      RECT 126 -182.675 126.4 -73.605 ;
      RECT 126 -64 126.4 -49.36 ;
      RECT 126 -45.51 126.4 -12.47 ;
      RECT 123.1 -80.215 123.5 -20.12 ;
      RECT 122.3 -79.355 122.7 -20.12 ;
      RECT 121.5 -182.675 121.9 -79.445 ;
      RECT 120.7 -63.5 121.1 -48.905 ;
      RECT 120.7 -45.08 121.1 -15.74 ;
      RECT 119.9 -182.675 120.3 -73.605 ;
      RECT 119.9 -64 120.3 -49.36 ;
      RECT 119.9 -45.51 120.3 -12.47 ;
      RECT 117 -80.215 117.4 -20.12 ;
      RECT 116.2 -79.355 116.6 -20.12 ;
      RECT 115.4 -182.675 115.8 -79.445 ;
      RECT 114.6 -63.5 115 -48.905 ;
      RECT 114.6 -45.08 115 -15.74 ;
      RECT 113.8 -182.675 114.2 -73.605 ;
      RECT 113.8 -64 114.2 -49.36 ;
      RECT 113.8 -45.51 114.2 -12.47 ;
      RECT 110.9 -80.215 111.3 -20.12 ;
      RECT 110.1 -79.355 110.5 -20.12 ;
      RECT 109.3 -182.675 109.7 -79.445 ;
      RECT 108.5 -63.5 108.9 -48.905 ;
      RECT 108.5 -45.08 108.9 -15.74 ;
      RECT 107.7 -182.675 108.1 -73.605 ;
      RECT 107.7 -64 108.1 -49.36 ;
      RECT 107.7 -45.51 108.1 -12.47 ;
      RECT 105.6 -87.06 106 -20.12 ;
      RECT 104.8 -80.215 105.2 -20.12 ;
      RECT 104 -182.675 104.4 -87.15 ;
      RECT 104 -79.355 104.4 -20.12 ;
      RECT 103.2 -182.675 103.6 -79.445 ;
      RECT 102.4 -63.5 102.8 -48.905 ;
      RECT 102.4 -45.08 102.8 -15.74 ;
      RECT 101.6 -182.675 102 -73.605 ;
      RECT 101.6 -64 102 -49.36 ;
      RECT 101.6 -45.51 102 -12.47 ;
      RECT 98.7 -80.215 99.1 -20.12 ;
      RECT 97.9 -79.355 98.3 -20.12 ;
      RECT 97.1 -182.675 97.5 -79.445 ;
      RECT 96.3 -63.5 96.7 -48.905 ;
      RECT 96.3 -45.08 96.7 -15.74 ;
      RECT 95.5 -182.675 95.9 -73.605 ;
      RECT 95.5 -64 95.9 -49.36 ;
      RECT 95.5 -45.51 95.9 -12.47 ;
      RECT 92.6 -80.215 93 -20.12 ;
      RECT 91.8 -79.355 92.2 -20.12 ;
      RECT 91 -182.675 91.4 -79.445 ;
      RECT 90.2 -63.5 90.6 -48.905 ;
      RECT 90.2 -45.08 90.6 -15.74 ;
      RECT 89.4 -182.675 89.8 -73.605 ;
      RECT 89.4 -64 89.8 -49.36 ;
      RECT 89.4 -45.51 89.8 -12.47 ;
      RECT 86.5 -80.215 86.9 -20.12 ;
      RECT 85.7 -79.355 86.1 -20.12 ;
      RECT 84.9 -182.675 85.3 -79.445 ;
      RECT 84.1 -63.5 84.5 -48.905 ;
      RECT 84.1 -45.08 84.5 -15.74 ;
      RECT 83.3 -182.675 83.7 -73.605 ;
      RECT 83.3 -64 83.7 -49.36 ;
      RECT 83.3 -45.51 83.7 -12.47 ;
      RECT 80.4 -80.215 80.8 -20.12 ;
      RECT 79.6 -79.355 80 -20.12 ;
      RECT 78.8 -182.675 79.2 -79.445 ;
      RECT 78 -63.5 78.4 -48.905 ;
      RECT 78 -45.08 78.4 -15.74 ;
      RECT 77.2 -182.675 77.6 -73.605 ;
      RECT 77.2 -64 77.6 -49.36 ;
      RECT 77.2 -45.51 77.6 -12.47 ;
      RECT 74.3 -80.215 74.7 -20.12 ;
      RECT 73.5 -79.355 73.9 -20.12 ;
      RECT 72.7 -182.675 73.1 -79.445 ;
      RECT 71.9 -63.5 72.3 -48.905 ;
      RECT 71.9 -45.08 72.3 -15.74 ;
      RECT 71.1 -182.675 71.5 -73.605 ;
      RECT 71.1 -64 71.5 -49.36 ;
      RECT 71.1 -45.51 71.5 -12.47 ;
      RECT 68.2 -80.215 68.6 -20.12 ;
      RECT 67.4 -79.355 67.8 -20.12 ;
      RECT 66.6 -182.675 67 -79.445 ;
      RECT 65.8 -63.5 66.2 -48.905 ;
      RECT 65.8 -45.08 66.2 -15.74 ;
      RECT 65 -182.675 65.4 -73.605 ;
      RECT 65 -64 65.4 -49.36 ;
      RECT 65 -45.51 65.4 -12.47 ;
      RECT 62.1 -80.215 62.5 -20.12 ;
      RECT 61.3 -79.355 61.7 -20.12 ;
      RECT 60.5 -182.675 60.9 -79.445 ;
      RECT 59.7 -63.5 60.1 -48.905 ;
      RECT 59.7 -45.08 60.1 -15.74 ;
      RECT 58.9 -182.675 59.3 -73.605 ;
      RECT 58.9 -64 59.3 -49.36 ;
      RECT 58.9 -45.51 59.3 -12.47 ;
      RECT 56.8 -87.06 57.2 -20.12 ;
      RECT 56 -80.215 56.4 -20.12 ;
      RECT 55.2 -182.675 55.6 -87.15 ;
      RECT 55.2 -79.355 55.6 -20.12 ;
      RECT 54.4 -182.675 54.8 -79.445 ;
      RECT 53.6 -63.5 54 -48.905 ;
      RECT 53.6 -45.08 54 -15.74 ;
      RECT 52.8 -182.675 53.2 -73.605 ;
      RECT 52.8 -64 53.2 -49.36 ;
      RECT 52.8 -45.51 53.2 -12.47 ;
      RECT 49.9 -80.215 50.3 -20.12 ;
      RECT 49.1 -79.355 49.5 -20.12 ;
      RECT 48.3 -182.675 48.7 -79.445 ;
      RECT 47.5 -63.5 47.9 -48.905 ;
      RECT 47.5 -45.08 47.9 -15.74 ;
      RECT 46.7 -182.675 47.1 -73.605 ;
      RECT 46.7 -64 47.1 -49.36 ;
      RECT 46.7 -45.51 47.1 -12.47 ;
      RECT 43.8 -80.215 44.2 -20.12 ;
      RECT 43 -79.355 43.4 -20.12 ;
      RECT 42.2 -182.675 42.6 -79.445 ;
      RECT 41.4 -63.5 41.8 -48.905 ;
      RECT 41.4 -45.08 41.8 -15.74 ;
      RECT 40.6 -182.675 41 -73.605 ;
      RECT 40.6 -64 41 -49.36 ;
      RECT 40.6 -45.51 41 -12.47 ;
      RECT 37.7 -80.215 38.1 -20.12 ;
      RECT 36.9 -79.355 37.3 -20.12 ;
      RECT 36.1 -182.675 36.5 -79.445 ;
      RECT 35.3 -63.5 35.7 -48.905 ;
      RECT 35.3 -45.08 35.7 -15.74 ;
      RECT 34.5 -182.675 34.9 -73.605 ;
      RECT 34.5 -64 34.9 -49.36 ;
      RECT 34.5 -45.51 34.9 -12.47 ;
      RECT 31.6 -80.215 32 -20.12 ;
      RECT 30.8 -79.355 31.2 -20.12 ;
      RECT 30 -182.675 30.4 -79.445 ;
      RECT 29.2 -63.5 29.6 -48.905 ;
      RECT 29.2 -45.08 29.6 -15.74 ;
      RECT 28.4 -182.675 28.8 -73.605 ;
      RECT 28.4 -64 28.8 -49.36 ;
      RECT 28.4 -45.51 28.8 -12.47 ;
      RECT 25.5 -80.215 25.9 -20.12 ;
      RECT 24.7 -79.355 25.1 -20.12 ;
      RECT 23.9 -182.675 24.3 -79.445 ;
      RECT 23.1 -63.5 23.5 -48.905 ;
      RECT 23.1 -45.08 23.5 -15.74 ;
      RECT 22.3 -182.675 22.7 -73.605 ;
      RECT 22.3 -64 22.7 -49.36 ;
      RECT 22.3 -45.51 22.7 -12.47 ;
      RECT 19.4 -80.215 19.8 -20.12 ;
      RECT 18.6 -79.355 19 -20.12 ;
      RECT 17.8 -182.675 18.2 -79.445 ;
      RECT 17 -63.5 17.4 -48.905 ;
      RECT 17 -45.08 17.4 -15.74 ;
      RECT 16.2 -182.675 16.6 -73.605 ;
      RECT 16.2 -64 16.6 -49.36 ;
      RECT 16.2 -45.51 16.6 -12.47 ;
      RECT 13.3 -80.215 13.7 -20.12 ;
      RECT 12.5 -79.355 12.9 -20.12 ;
      RECT 11.7 -182.675 12.1 -79.445 ;
      RECT 10.9 -63.5 11.3 -48.905 ;
      RECT 10.9 -45.08 11.3 -15.74 ;
      RECT 10.1 -182.675 10.5 -73.605 ;
      RECT 10.1 -64 10.5 -49.36 ;
      RECT 10.1 -45.51 10.5 -12.47 ;
      RECT 8 -87.06 8.4 -20.12 ;
      RECT 7.2 -80.215 7.6 -20.12 ;
      RECT 6.4 -182.675 6.8 -87.15 ;
      RECT 6.4 -79.355 6.8 -20.12 ;
      RECT 5.6 -182.675 6 -79.445 ;
      RECT 4.8 -63.5 5.2 -48.905 ;
      RECT 4.8 -45.08 5.2 -15.74 ;
      RECT 4 -182.675 4.4 -73.605 ;
      RECT 4 -64 4.4 -49.36 ;
      RECT 4 -45.51 4.4 -12.47 ;
  END
END sram22_512x64m4w8

END LIBRARY
